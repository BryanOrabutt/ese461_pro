module mult (clk, rst, A, B, out, start_mac);
  input clk;
  input rst; 
  input wire start_mac;
  input signed [15:0]A, B;
  output signed [15:0]out;
  reg signed [31:0] PRODUCT;
  reg [15:0]x1,x2;

  assign out = {PRODUCT[31], PRODUCT[22:8]};

always @(posedge clk ) begin
    if (rst) begin
      PRODUCT = 0;
        x1 = 0;
        x2 = 0;
    end else begin
	if (start_mac) begin
        x1 =((A[15]==0)?{1'b0,A[14:0]}:{1'b0,~(A[14:0]-1'b1)});
        x2 =((B[15]==0)?{1'b0,B[14:0]}:{1'b0,~(B[14:0]-1'b1)});
        PRODUCT=
              (A[15]^B[15]==0)?
              (
                (x2[0]? {15'b0,x1[15:0]}:      32'b0)+
                (x2[1]? {14'b0,x1[15:0], 1'b0}:32'b0)+
                (x2[2]? {13'b0,x1[15:0], 2'b0}:32'b0)+
                (x2[3]? {12'b0,x1[15:0], 3'b0}:32'b0)+
                (x2[4]? {11'b0,x1[15:0], 4'b0}:32'b0)+
                (x2[5]? {10'b0,x1[15:0], 5'b0}:32'b0)+
                (x2[6]? {9 'b0,x1[15:0], 6'b0}:32'b0)+
                (x2[7]? {8 'b0,x1[15:0], 7'b0}:32'b0)+
                (x2[8]? {7 'b0,x1[15:0], 8'b0}:32'b0)+
                (x2[9]? {6 'b0,x1[15:0], 9'b0}:32'b0)+
                (x2[10]?{5 'b0,x1[15:0],10'b0}:32'b0)+
                (x2[11]?{4 'b0,x1[15:0],11'b0}:32'b0)+
                (x2[12]?{3 'b0,x1[15:0],12'b0}:32'b0)+
                (x2[13]?{2 'b0,x1[15:0],13'b0}:32'b0)+
                (x2[14]?{1 'b0,x1[15:0],14'b0}:32'b0)+
                (x2[15]?{      x1[15:0],15'b0}:32'b0)
              ):(~(
                (x2[0]? {15'b0,x1[15:0]}:      32'b0)+
                (x2[1]? {14'b0,x1[15:0], 1'b0}:32'b0)+
                (x2[2]? {13'b0,x1[15:0], 2'b0}:32'b0)+
                (x2[3]? {12'b0,x1[15:0], 3'b0}:32'b0)+
                (x2[4]? {11'b0,x1[15:0], 4'b0}:32'b0)+
                (x2[5]? {10'b0,x1[15:0], 5'b0}:32'b0)+
                (x2[6]? {9 'b0,x1[15:0], 6'b0}:32'b0)+
                (x2[7]? {8 'b0,x1[15:0], 7'b0}:32'b0)+
                (x2[8]? {7 'b0,x1[15:0], 8'b0}:32'b0)+
                (x2[9]? {6 'b0,x1[15:0], 9'b0}:32'b0)+
                (x2[10]?{5 'b0,x1[15:0],10'b0}:32'b0)+
                (x2[11]?{4 'b0,x1[15:0],11'b0}:32'b0)+
                (x2[12]?{3 'b0,x1[15:0],12'b0}:32'b0)+
                (x2[13]?{2 'b0,x1[15:0],13'b0}:32'b0)+
                (x2[14]?{1 'b0,x1[15:0],14'b0}:32'b0)+
                (x2[15]?{      x1[15:0],15'b0}:32'b0))   
              );
        PRODUCT[31]=A[15]^B[15];
        PRODUCT=PRODUCT[31]?PRODUCT+1'b1:PRODUCT;
        //PRODUCT <= A*B;
		end
    end
  end
endmodule





