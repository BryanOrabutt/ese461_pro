

module ReadOnlyMemory_I(output reg [15:0] data_out, input [16:0] address);
always@(address)begin
	case(address) 
17'h0:	data_out=16'h1;
17'h1:	data_out=16'h0;
17'h2:	data_out=16'h0;
17'h3:	data_out=16'h0;
17'h4:	data_out=16'h0;
17'h5:	data_out=16'h0;
17'h6:	data_out=16'h0;
17'h7:	data_out=16'h0;
17'h8:	data_out=16'h0;
17'h9:	data_out=16'h0;
17'ha:	data_out=16'h0;
17'hb:	data_out=16'h0;
17'hc:	data_out=16'h0;
17'hd:	data_out=16'h0;
17'he:	data_out=16'h0;
17'hf:	data_out=16'h0;
17'h10:	data_out=16'h0;
17'h11:	data_out=16'h0;
17'h12:	data_out=16'h0;
17'h13:	data_out=16'h0;
17'h14:	data_out=16'h0;
17'h15:	data_out=16'h0;
17'h16:	data_out=16'h0;
17'h17:	data_out=16'h0;
17'h18:	data_out=16'h0;
17'h19:	data_out=16'h0;
17'h1a:	data_out=16'h0;
17'h1b:	data_out=16'h0;
17'h1c:	data_out=16'h0;
17'h1d:	data_out=16'h0;
17'h1e:	data_out=16'h0;
17'h1f:	data_out=16'h0;
17'h20:	data_out=16'h0;
17'h21:	data_out=16'h0;
17'h22:	data_out=16'h0;
17'h23:	data_out=16'h0;
17'h24:	data_out=16'h0;
17'h25:	data_out=16'h0;
17'h26:	data_out=16'h0;
17'h27:	data_out=16'h0;
17'h28:	data_out=16'h0;
17'h29:	data_out=16'h0;
17'h2a:	data_out=16'h0;
17'h2b:	data_out=16'h0;
17'h2c:	data_out=16'h0;
17'h2d:	data_out=16'h0;
17'h2e:	data_out=16'h0;
17'h2f:	data_out=16'h0;
17'h30:	data_out=16'h0;
17'h31:	data_out=16'h0;
17'h32:	data_out=16'h0;
17'h33:	data_out=16'h0;
17'h34:	data_out=16'h0;
17'h35:	data_out=16'h0;
17'h36:	data_out=16'h0;
17'h37:	data_out=16'h0;
17'h38:	data_out=16'h0;
17'h39:	data_out=16'h0;
17'h3a:	data_out=16'h0;
17'h3b:	data_out=16'h0;
17'h3c:	data_out=16'h0;
17'h3d:	data_out=16'h0;
17'h3e:	data_out=16'h0;
17'h3f:	data_out=16'h0;
17'h40:	data_out=16'h0;
17'h41:	data_out=16'h0;
17'h42:	data_out=16'h0;
17'h43:	data_out=16'h0;
17'h44:	data_out=16'h0;
17'h45:	data_out=16'h0;
17'h46:	data_out=16'h0;
17'h47:	data_out=16'h0;
17'h48:	data_out=16'h0;
17'h49:	data_out=16'h0;
17'h4a:	data_out=16'h0;
17'h4b:	data_out=16'h0;
17'h4c:	data_out=16'h0;
17'h4d:	data_out=16'h0;
17'h4e:	data_out=16'h0;
17'h4f:	data_out=16'h0;
17'h50:	data_out=16'h0;
17'h51:	data_out=16'h0;
17'h52:	data_out=16'h0;
17'h53:	data_out=16'h0;
17'h54:	data_out=16'h0;
17'h55:	data_out=16'h0;
17'h56:	data_out=16'h0;
17'h57:	data_out=16'h0;
17'h58:	data_out=16'h0;
17'h59:	data_out=16'h0;
17'h5a:	data_out=16'h0;
17'h5b:	data_out=16'h0;
17'h5c:	data_out=16'h0;
17'h5d:	data_out=16'h0;
17'h5e:	data_out=16'h0;
17'h5f:	data_out=16'h0;
17'h60:	data_out=16'h0;
17'h61:	data_out=16'h0;
17'h62:	data_out=16'h0;
17'h63:	data_out=16'h0;
17'h64:	data_out=16'h0;
17'h65:	data_out=16'h0;
17'h66:	data_out=16'h0;
17'h67:	data_out=16'h0;
17'h68:	data_out=16'h0;
17'h69:	data_out=16'h0;
17'h6a:	data_out=16'h0;
17'h6b:	data_out=16'h0;
17'h6c:	data_out=16'h0;
17'h6d:	data_out=16'h0;
17'h6e:	data_out=16'h0;
17'h6f:	data_out=16'h0;
17'h70:	data_out=16'h0;
17'h71:	data_out=16'h0;
17'h72:	data_out=16'h0;
17'h73:	data_out=16'h0;
17'h74:	data_out=16'h0;
17'h75:	data_out=16'h0;
17'h76:	data_out=16'h0;
17'h77:	data_out=16'h0;
17'h78:	data_out=16'h0;
17'h79:	data_out=16'h0;
17'h7a:	data_out=16'h0;
17'h7b:	data_out=16'h0;
17'h7c:	data_out=16'h0;
17'h7d:	data_out=16'h0;
17'h7e:	data_out=16'h0;
17'h7f:	data_out=16'h0;
17'h80:	data_out=16'h0;
17'h81:	data_out=16'h0;
17'h82:	data_out=16'h0;
17'h83:	data_out=16'h0;
17'h84:	data_out=16'h0;
17'h85:	data_out=16'h0;
17'h86:	data_out=16'h0;
17'h87:	data_out=16'h0;
17'h88:	data_out=16'h0;
17'h89:	data_out=16'h0;
17'h8a:	data_out=16'h0;
17'h8b:	data_out=16'h0;
17'h8c:	data_out=16'h0;
17'h8d:	data_out=16'h0;
17'h8e:	data_out=16'h0;
17'h8f:	data_out=16'h0;
17'h90:	data_out=16'h0;
17'h91:	data_out=16'h0;
17'h92:	data_out=16'h0;
17'h93:	data_out=16'h0;
17'h94:	data_out=16'h0;
17'h95:	data_out=16'h0;
17'h96:	data_out=16'h0;
17'h97:	data_out=16'h0;
17'h98:	data_out=16'h3;
17'h99:	data_out=16'h12;
17'h9a:	data_out=16'h12;
17'h9b:	data_out=16'h12;
17'h9c:	data_out=16'h7e;
17'h9d:	data_out=16'h89;
17'h9e:	data_out=16'hb0;
17'h9f:	data_out=16'h1a;
17'ha0:	data_out=16'ha7;
17'ha1:	data_out=16'h100;
17'ha2:	data_out=16'hf8;
17'ha3:	data_out=16'h7f;
17'ha4:	data_out=16'h0;
17'ha5:	data_out=16'h0;
17'ha6:	data_out=16'h0;
17'ha7:	data_out=16'h0;
17'ha8:	data_out=16'h0;
17'ha9:	data_out=16'h0;
17'haa:	data_out=16'h0;
17'hab:	data_out=16'h0;
17'hac:	data_out=16'h0;
17'had:	data_out=16'h0;
17'hae:	data_out=16'h0;
17'haf:	data_out=16'h0;
17'hb0:	data_out=16'h1e;
17'hb1:	data_out=16'h24;
17'hb2:	data_out=16'h5e;
17'hb3:	data_out=16'h9b;
17'hb4:	data_out=16'hab;
17'hb5:	data_out=16'hfe;
17'hb6:	data_out=16'hfe;
17'hb7:	data_out=16'hfe;
17'hb8:	data_out=16'hfe;
17'hb9:	data_out=16'hfe;
17'hba:	data_out=16'he2;
17'hbb:	data_out=16'had;
17'hbc:	data_out=16'hfe;
17'hbd:	data_out=16'hf3;
17'hbe:	data_out=16'hc4;
17'hbf:	data_out=16'h40;
17'hc0:	data_out=16'h0;
17'hc1:	data_out=16'h0;
17'hc2:	data_out=16'h0;
17'hc3:	data_out=16'h0;
17'hc4:	data_out=16'h0;
17'hc5:	data_out=16'h0;
17'hc6:	data_out=16'h0;
17'hc7:	data_out=16'h0;
17'hc8:	data_out=16'h0;
17'hc9:	data_out=16'h0;
17'hca:	data_out=16'h0;
17'hcb:	data_out=16'h31;
17'hcc:	data_out=16'hef;
17'hcd:	data_out=16'hfe;
17'hce:	data_out=16'hfe;
17'hcf:	data_out=16'hfe;
17'hd0:	data_out=16'hfe;
17'hd1:	data_out=16'hfe;
17'hd2:	data_out=16'hfe;
17'hd3:	data_out=16'hfe;
17'hd4:	data_out=16'hfe;
17'hd5:	data_out=16'hfc;
17'hd6:	data_out=16'h5d;
17'hd7:	data_out=16'h52;
17'hd8:	data_out=16'h52;
17'hd9:	data_out=16'h38;
17'hda:	data_out=16'h27;
17'hdb:	data_out=16'h0;
17'hdc:	data_out=16'h0;
17'hdd:	data_out=16'h0;
17'hde:	data_out=16'h0;
17'hdf:	data_out=16'h0;
17'he0:	data_out=16'h0;
17'he1:	data_out=16'h0;
17'he2:	data_out=16'h0;
17'he3:	data_out=16'h0;
17'he4:	data_out=16'h0;
17'he5:	data_out=16'h0;
17'he6:	data_out=16'h0;
17'he7:	data_out=16'h12;
17'he8:	data_out=16'hdc;
17'he9:	data_out=16'hfe;
17'hea:	data_out=16'hfe;
17'heb:	data_out=16'hfe;
17'hec:	data_out=16'hfe;
17'hed:	data_out=16'hfe;
17'hee:	data_out=16'hc7;
17'hef:	data_out=16'hb7;
17'hf0:	data_out=16'hf8;
17'hf1:	data_out=16'hf2;
17'hf2:	data_out=16'h0;
17'hf3:	data_out=16'h0;
17'hf4:	data_out=16'h0;
17'hf5:	data_out=16'h0;
17'hf6:	data_out=16'h0;
17'hf7:	data_out=16'h0;
17'hf8:	data_out=16'h0;
17'hf9:	data_out=16'h0;
17'hfa:	data_out=16'h0;
17'hfb:	data_out=16'h0;
17'hfc:	data_out=16'h0;
17'hfd:	data_out=16'h0;
17'hfe:	data_out=16'h0;
17'hff:	data_out=16'h0;
17'h100:	data_out=16'h0;
17'h101:	data_out=16'h0;
17'h102:	data_out=16'h0;
17'h103:	data_out=16'h0;
17'h104:	data_out=16'h50;
17'h105:	data_out=16'h9d;
17'h106:	data_out=16'h6b;
17'h107:	data_out=16'hfe;
17'h108:	data_out=16'hfe;
17'h109:	data_out=16'hce;
17'h10a:	data_out=16'hb;
17'h10b:	data_out=16'h0;
17'h10c:	data_out=16'h2b;
17'h10d:	data_out=16'h9b;
17'h10e:	data_out=16'h0;
17'h10f:	data_out=16'h0;
17'h110:	data_out=16'h0;
17'h111:	data_out=16'h0;
17'h112:	data_out=16'h0;
17'h113:	data_out=16'h0;
17'h114:	data_out=16'h0;
17'h115:	data_out=16'h0;
17'h116:	data_out=16'h0;
17'h117:	data_out=16'h0;
17'h118:	data_out=16'h0;
17'h119:	data_out=16'h0;
17'h11a:	data_out=16'h0;
17'h11b:	data_out=16'h0;
17'h11c:	data_out=16'h0;
17'h11d:	data_out=16'h0;
17'h11e:	data_out=16'h0;
17'h11f:	data_out=16'h0;
17'h120:	data_out=16'h0;
17'h121:	data_out=16'he;
17'h122:	data_out=16'h1;
17'h123:	data_out=16'h9b;
17'h124:	data_out=16'hfe;
17'h125:	data_out=16'h5a;
17'h126:	data_out=16'h0;
17'h127:	data_out=16'h0;
17'h128:	data_out=16'h0;
17'h129:	data_out=16'h0;
17'h12a:	data_out=16'h0;
17'h12b:	data_out=16'h0;
17'h12c:	data_out=16'h0;
17'h12d:	data_out=16'h0;
17'h12e:	data_out=16'h0;
17'h12f:	data_out=16'h0;
17'h130:	data_out=16'h0;
17'h131:	data_out=16'h0;
17'h132:	data_out=16'h0;
17'h133:	data_out=16'h0;
17'h134:	data_out=16'h0;
17'h135:	data_out=16'h0;
17'h136:	data_out=16'h0;
17'h137:	data_out=16'h0;
17'h138:	data_out=16'h0;
17'h139:	data_out=16'h0;
17'h13a:	data_out=16'h0;
17'h13b:	data_out=16'h0;
17'h13c:	data_out=16'h0;
17'h13d:	data_out=16'h0;
17'h13e:	data_out=16'h0;
17'h13f:	data_out=16'h8c;
17'h140:	data_out=16'hfe;
17'h141:	data_out=16'hbf;
17'h142:	data_out=16'h2;
17'h143:	data_out=16'h0;
17'h144:	data_out=16'h0;
17'h145:	data_out=16'h0;
17'h146:	data_out=16'h0;
17'h147:	data_out=16'h0;
17'h148:	data_out=16'h0;
17'h149:	data_out=16'h0;
17'h14a:	data_out=16'h0;
17'h14b:	data_out=16'h0;
17'h14c:	data_out=16'h0;
17'h14d:	data_out=16'h0;
17'h14e:	data_out=16'h0;
17'h14f:	data_out=16'h0;
17'h150:	data_out=16'h0;
17'h151:	data_out=16'h0;
17'h152:	data_out=16'h0;
17'h153:	data_out=16'h0;
17'h154:	data_out=16'h0;
17'h155:	data_out=16'h0;
17'h156:	data_out=16'h0;
17'h157:	data_out=16'h0;
17'h158:	data_out=16'h0;
17'h159:	data_out=16'h0;
17'h15a:	data_out=16'h0;
17'h15b:	data_out=16'hb;
17'h15c:	data_out=16'hbf;
17'h15d:	data_out=16'hfe;
17'h15e:	data_out=16'h46;
17'h15f:	data_out=16'h0;
17'h160:	data_out=16'h0;
17'h161:	data_out=16'h0;
17'h162:	data_out=16'h0;
17'h163:	data_out=16'h0;
17'h164:	data_out=16'h0;
17'h165:	data_out=16'h0;
17'h166:	data_out=16'h0;
17'h167:	data_out=16'h0;
17'h168:	data_out=16'h0;
17'h169:	data_out=16'h0;
17'h16a:	data_out=16'h0;
17'h16b:	data_out=16'h0;
17'h16c:	data_out=16'h0;
17'h16d:	data_out=16'h0;
17'h16e:	data_out=16'h0;
17'h16f:	data_out=16'h0;
17'h170:	data_out=16'h0;
17'h171:	data_out=16'h0;
17'h172:	data_out=16'h0;
17'h173:	data_out=16'h0;
17'h174:	data_out=16'h0;
17'h175:	data_out=16'h0;
17'h176:	data_out=16'h0;
17'h177:	data_out=16'h0;
17'h178:	data_out=16'h23;
17'h179:	data_out=16'hf2;
17'h17a:	data_out=16'he2;
17'h17b:	data_out=16'ha1;
17'h17c:	data_out=16'h6c;
17'h17d:	data_out=16'h1;
17'h17e:	data_out=16'h0;
17'h17f:	data_out=16'h0;
17'h180:	data_out=16'h0;
17'h181:	data_out=16'h0;
17'h182:	data_out=16'h0;
17'h183:	data_out=16'h0;
17'h184:	data_out=16'h0;
17'h185:	data_out=16'h0;
17'h186:	data_out=16'h0;
17'h187:	data_out=16'h0;
17'h188:	data_out=16'h0;
17'h189:	data_out=16'h0;
17'h18a:	data_out=16'h0;
17'h18b:	data_out=16'h0;
17'h18c:	data_out=16'h0;
17'h18d:	data_out=16'h0;
17'h18e:	data_out=16'h0;
17'h18f:	data_out=16'h0;
17'h190:	data_out=16'h0;
17'h191:	data_out=16'h0;
17'h192:	data_out=16'h0;
17'h193:	data_out=16'h0;
17'h194:	data_out=16'h0;
17'h195:	data_out=16'h51;
17'h196:	data_out=16'hf1;
17'h197:	data_out=16'hfe;
17'h198:	data_out=16'hfe;
17'h199:	data_out=16'h77;
17'h19a:	data_out=16'h19;
17'h19b:	data_out=16'h0;
17'h19c:	data_out=16'h0;
17'h19d:	data_out=16'h0;
17'h19e:	data_out=16'h0;
17'h19f:	data_out=16'h0;
17'h1a0:	data_out=16'h0;
17'h1a1:	data_out=16'h0;
17'h1a2:	data_out=16'h0;
17'h1a3:	data_out=16'h0;
17'h1a4:	data_out=16'h0;
17'h1a5:	data_out=16'h0;
17'h1a6:	data_out=16'h0;
17'h1a7:	data_out=16'h0;
17'h1a8:	data_out=16'h0;
17'h1a9:	data_out=16'h0;
17'h1aa:	data_out=16'h0;
17'h1ab:	data_out=16'h0;
17'h1ac:	data_out=16'h0;
17'h1ad:	data_out=16'h0;
17'h1ae:	data_out=16'h0;
17'h1af:	data_out=16'h0;
17'h1b0:	data_out=16'h0;
17'h1b1:	data_out=16'h0;
17'h1b2:	data_out=16'h2d;
17'h1b3:	data_out=16'hbb;
17'h1b4:	data_out=16'hfe;
17'h1b5:	data_out=16'hfe;
17'h1b6:	data_out=16'h97;
17'h1b7:	data_out=16'h1b;
17'h1b8:	data_out=16'h0;
17'h1b9:	data_out=16'h0;
17'h1ba:	data_out=16'h0;
17'h1bb:	data_out=16'h0;
17'h1bc:	data_out=16'h0;
17'h1bd:	data_out=16'h0;
17'h1be:	data_out=16'h0;
17'h1bf:	data_out=16'h0;
17'h1c0:	data_out=16'h0;
17'h1c1:	data_out=16'h0;
17'h1c2:	data_out=16'h0;
17'h1c3:	data_out=16'h0;
17'h1c4:	data_out=16'h0;
17'h1c5:	data_out=16'h0;
17'h1c6:	data_out=16'h0;
17'h1c7:	data_out=16'h0;
17'h1c8:	data_out=16'h0;
17'h1c9:	data_out=16'h0;
17'h1ca:	data_out=16'h0;
17'h1cb:	data_out=16'h0;
17'h1cc:	data_out=16'h0;
17'h1cd:	data_out=16'h0;
17'h1ce:	data_out=16'h0;
17'h1cf:	data_out=16'h10;
17'h1d0:	data_out=16'h5d;
17'h1d1:	data_out=16'hfd;
17'h1d2:	data_out=16'hfe;
17'h1d3:	data_out=16'hbc;
17'h1d4:	data_out=16'h0;
17'h1d5:	data_out=16'h0;
17'h1d6:	data_out=16'h0;
17'h1d7:	data_out=16'h0;
17'h1d8:	data_out=16'h0;
17'h1d9:	data_out=16'h0;
17'h1da:	data_out=16'h0;
17'h1db:	data_out=16'h0;
17'h1dc:	data_out=16'h0;
17'h1dd:	data_out=16'h0;
17'h1de:	data_out=16'h0;
17'h1df:	data_out=16'h0;
17'h1e0:	data_out=16'h0;
17'h1e1:	data_out=16'h0;
17'h1e2:	data_out=16'h0;
17'h1e3:	data_out=16'h0;
17'h1e4:	data_out=16'h0;
17'h1e5:	data_out=16'h0;
17'h1e6:	data_out=16'h0;
17'h1e7:	data_out=16'h0;
17'h1e8:	data_out=16'h0;
17'h1e9:	data_out=16'h0;
17'h1ea:	data_out=16'h0;
17'h1eb:	data_out=16'h0;
17'h1ec:	data_out=16'h0;
17'h1ed:	data_out=16'hfa;
17'h1ee:	data_out=16'hfe;
17'h1ef:	data_out=16'hfa;
17'h1f0:	data_out=16'h40;
17'h1f1:	data_out=16'h0;
17'h1f2:	data_out=16'h0;
17'h1f3:	data_out=16'h0;
17'h1f4:	data_out=16'h0;
17'h1f5:	data_out=16'h0;
17'h1f6:	data_out=16'h0;
17'h1f7:	data_out=16'h0;
17'h1f8:	data_out=16'h0;
17'h1f9:	data_out=16'h0;
17'h1fa:	data_out=16'h0;
17'h1fb:	data_out=16'h0;
17'h1fc:	data_out=16'h0;
17'h1fd:	data_out=16'h0;
17'h1fe:	data_out=16'h0;
17'h1ff:	data_out=16'h0;
17'h200:	data_out=16'h0;
17'h201:	data_out=16'h0;
17'h202:	data_out=16'h0;
17'h203:	data_out=16'h0;
17'h204:	data_out=16'h0;
17'h205:	data_out=16'h0;
17'h206:	data_out=16'h2e;
17'h207:	data_out=16'h83;
17'h208:	data_out=16'hb8;
17'h209:	data_out=16'hfe;
17'h20a:	data_out=16'hfe;
17'h20b:	data_out=16'hd0;
17'h20c:	data_out=16'h2;
17'h20d:	data_out=16'h0;
17'h20e:	data_out=16'h0;
17'h20f:	data_out=16'h0;
17'h210:	data_out=16'h0;
17'h211:	data_out=16'h0;
17'h212:	data_out=16'h0;
17'h213:	data_out=16'h0;
17'h214:	data_out=16'h0;
17'h215:	data_out=16'h0;
17'h216:	data_out=16'h0;
17'h217:	data_out=16'h0;
17'h218:	data_out=16'h0;
17'h219:	data_out=16'h0;
17'h21a:	data_out=16'h0;
17'h21b:	data_out=16'h0;
17'h21c:	data_out=16'h0;
17'h21d:	data_out=16'h0;
17'h21e:	data_out=16'h0;
17'h21f:	data_out=16'h0;
17'h220:	data_out=16'h27;
17'h221:	data_out=16'h95;
17'h222:	data_out=16'he6;
17'h223:	data_out=16'hfe;
17'h224:	data_out=16'hfe;
17'h225:	data_out=16'hfe;
17'h226:	data_out=16'hfb;
17'h227:	data_out=16'hb7;
17'h228:	data_out=16'h0;
17'h229:	data_out=16'h0;
17'h22a:	data_out=16'h0;
17'h22b:	data_out=16'h0;
17'h22c:	data_out=16'h0;
17'h22d:	data_out=16'h0;
17'h22e:	data_out=16'h0;
17'h22f:	data_out=16'h0;
17'h230:	data_out=16'h0;
17'h231:	data_out=16'h0;
17'h232:	data_out=16'h0;
17'h233:	data_out=16'h0;
17'h234:	data_out=16'h0;
17'h235:	data_out=16'h0;
17'h236:	data_out=16'h0;
17'h237:	data_out=16'h0;
17'h238:	data_out=16'h0;
17'h239:	data_out=16'h0;
17'h23a:	data_out=16'h18;
17'h23b:	data_out=16'h72;
17'h23c:	data_out=16'hde;
17'h23d:	data_out=16'hfe;
17'h23e:	data_out=16'hfe;
17'h23f:	data_out=16'hfe;
17'h240:	data_out=16'hfe;
17'h241:	data_out=16'hca;
17'h242:	data_out=16'h4e;
17'h243:	data_out=16'h0;
17'h244:	data_out=16'h0;
17'h245:	data_out=16'h0;
17'h246:	data_out=16'h0;
17'h247:	data_out=16'h0;
17'h248:	data_out=16'h0;
17'h249:	data_out=16'h0;
17'h24a:	data_out=16'h0;
17'h24b:	data_out=16'h0;
17'h24c:	data_out=16'h0;
17'h24d:	data_out=16'h0;
17'h24e:	data_out=16'h0;
17'h24f:	data_out=16'h0;
17'h250:	data_out=16'h0;
17'h251:	data_out=16'h0;
17'h252:	data_out=16'h0;
17'h253:	data_out=16'h0;
17'h254:	data_out=16'h17;
17'h255:	data_out=16'h42;
17'h256:	data_out=16'hd6;
17'h257:	data_out=16'hfe;
17'h258:	data_out=16'hfe;
17'h259:	data_out=16'hfe;
17'h25a:	data_out=16'hfe;
17'h25b:	data_out=16'hc7;
17'h25c:	data_out=16'h51;
17'h25d:	data_out=16'h2;
17'h25e:	data_out=16'h0;
17'h25f:	data_out=16'h0;
17'h260:	data_out=16'h0;
17'h261:	data_out=16'h0;
17'h262:	data_out=16'h0;
17'h263:	data_out=16'h0;
17'h264:	data_out=16'h0;
17'h265:	data_out=16'h0;
17'h266:	data_out=16'h0;
17'h267:	data_out=16'h0;
17'h268:	data_out=16'h0;
17'h269:	data_out=16'h0;
17'h26a:	data_out=16'h0;
17'h26b:	data_out=16'h0;
17'h26c:	data_out=16'h0;
17'h26d:	data_out=16'h0;
17'h26e:	data_out=16'h12;
17'h26f:	data_out=16'hac;
17'h270:	data_out=16'hdc;
17'h271:	data_out=16'hfe;
17'h272:	data_out=16'hfe;
17'h273:	data_out=16'hfe;
17'h274:	data_out=16'hfe;
17'h275:	data_out=16'hc4;
17'h276:	data_out=16'h50;
17'h277:	data_out=16'h9;
17'h278:	data_out=16'h0;
17'h279:	data_out=16'h0;
17'h27a:	data_out=16'h0;
17'h27b:	data_out=16'h0;
17'h27c:	data_out=16'h0;
17'h27d:	data_out=16'h0;
17'h27e:	data_out=16'h0;
17'h27f:	data_out=16'h0;
17'h280:	data_out=16'h0;
17'h281:	data_out=16'h0;
17'h282:	data_out=16'h0;
17'h283:	data_out=16'h0;
17'h284:	data_out=16'h0;
17'h285:	data_out=16'h0;
17'h286:	data_out=16'h0;
17'h287:	data_out=16'h0;
17'h288:	data_out=16'h37;
17'h289:	data_out=16'had;
17'h28a:	data_out=16'he3;
17'h28b:	data_out=16'hfe;
17'h28c:	data_out=16'hfe;
17'h28d:	data_out=16'hfe;
17'h28e:	data_out=16'hfe;
17'h28f:	data_out=16'hf5;
17'h290:	data_out=16'h86;
17'h291:	data_out=16'hb;
17'h292:	data_out=16'h0;
17'h293:	data_out=16'h0;
17'h294:	data_out=16'h0;
17'h295:	data_out=16'h0;
17'h296:	data_out=16'h0;
17'h297:	data_out=16'h0;
17'h298:	data_out=16'h0;
17'h299:	data_out=16'h0;
17'h29a:	data_out=16'h0;
17'h29b:	data_out=16'h0;
17'h29c:	data_out=16'h0;
17'h29d:	data_out=16'h0;
17'h29e:	data_out=16'h0;
17'h29f:	data_out=16'h0;
17'h2a0:	data_out=16'h0;
17'h2a1:	data_out=16'h0;
17'h2a2:	data_out=16'h0;
17'h2a3:	data_out=16'h0;
17'h2a4:	data_out=16'h89;
17'h2a5:	data_out=16'hfe;
17'h2a6:	data_out=16'hfe;
17'h2a7:	data_out=16'hfe;
17'h2a8:	data_out=16'hd5;
17'h2a9:	data_out=16'h88;
17'h2aa:	data_out=16'h85;
17'h2ab:	data_out=16'h10;
17'h2ac:	data_out=16'h0;
17'h2ad:	data_out=16'h0;
17'h2ae:	data_out=16'h0;
17'h2af:	data_out=16'h0;
17'h2b0:	data_out=16'h0;
17'h2b1:	data_out=16'h0;
17'h2b2:	data_out=16'h0;
17'h2b3:	data_out=16'h0;
17'h2b4:	data_out=16'h0;
17'h2b5:	data_out=16'h0;
17'h2b6:	data_out=16'h0;
17'h2b7:	data_out=16'h0;
17'h2b8:	data_out=16'h0;
17'h2b9:	data_out=16'h0;
17'h2ba:	data_out=16'h0;
17'h2bb:	data_out=16'h0;
17'h2bc:	data_out=16'h0;
17'h2bd:	data_out=16'h0;
17'h2be:	data_out=16'h0;
17'h2bf:	data_out=16'h0;
17'h2c0:	data_out=16'h0;
17'h2c1:	data_out=16'h0;
17'h2c2:	data_out=16'h0;
17'h2c3:	data_out=16'h0;
17'h2c4:	data_out=16'h0;
17'h2c5:	data_out=16'h0;
17'h2c6:	data_out=16'h0;
17'h2c7:	data_out=16'h0;
17'h2c8:	data_out=16'h0;
17'h2c9:	data_out=16'h0;
17'h2ca:	data_out=16'h0;
17'h2cb:	data_out=16'h0;
17'h2cc:	data_out=16'h0;
17'h2cd:	data_out=16'h0;
17'h2ce:	data_out=16'h0;
17'h2cf:	data_out=16'h0;
17'h2d0:	data_out=16'h0;
17'h2d1:	data_out=16'h0;
17'h2d2:	data_out=16'h0;
17'h2d3:	data_out=16'h0;
17'h2d4:	data_out=16'h0;
17'h2d5:	data_out=16'h0;
17'h2d6:	data_out=16'h0;
17'h2d7:	data_out=16'h0;
17'h2d8:	data_out=16'h0;
17'h2d9:	data_out=16'h0;
17'h2da:	data_out=16'h0;
17'h2db:	data_out=16'h0;
17'h2dc:	data_out=16'h0;
17'h2dd:	data_out=16'h0;
17'h2de:	data_out=16'h0;
17'h2df:	data_out=16'h0;
17'h2e0:	data_out=16'h0;
17'h2e1:	data_out=16'h0;
17'h2e2:	data_out=16'h0;
17'h2e3:	data_out=16'h0;
17'h2e4:	data_out=16'h0;
17'h2e5:	data_out=16'h0;
17'h2e6:	data_out=16'h0;
17'h2e7:	data_out=16'h0;
17'h2e8:	data_out=16'h0;
17'h2e9:	data_out=16'h0;
17'h2ea:	data_out=16'h0;
17'h2eb:	data_out=16'h0;
17'h2ec:	data_out=16'h0;
17'h2ed:	data_out=16'h0;
17'h2ee:	data_out=16'h0;
17'h2ef:	data_out=16'h0;
17'h2f0:	data_out=16'h0;
17'h2f1:	data_out=16'h0;
17'h2f2:	data_out=16'h0;
17'h2f3:	data_out=16'h0;
17'h2f4:	data_out=16'h0;
17'h2f5:	data_out=16'h0;
17'h2f6:	data_out=16'h0;
17'h2f7:	data_out=16'h0;
17'h2f8:	data_out=16'h0;
17'h2f9:	data_out=16'h0;
17'h2fa:	data_out=16'h0;
17'h2fb:	data_out=16'h0;
17'h2fc:	data_out=16'h0;
17'h2fd:	data_out=16'h0;
17'h2fe:	data_out=16'h0;
17'h2ff:	data_out=16'h0;
17'h300:	data_out=16'h0;
17'h301:	data_out=16'h0;
17'h302:	data_out=16'h0;
17'h303:	data_out=16'h0;
17'h304:	data_out=16'h0;
17'h305:	data_out=16'h0;
17'h306:	data_out=16'h0;
17'h307:	data_out=16'h0;
17'h308:	data_out=16'h0;
17'h309:	data_out=16'h0;
17'h30a:	data_out=16'h0;
17'h30b:	data_out=16'h0;
17'h30c:	data_out=16'h0;
17'h30d:	data_out=16'h0;
17'h30e:	data_out=16'h0;
17'h30f:	data_out=16'h0;
17'h310:	data_out=16'h0;
17'h311:	data_out=16'h0;
17'h312:	data_out=16'h0;
17'h313:	data_out=16'h0;
17'h314:	data_out=16'h0;
17'h315:	data_out=16'h0;
17'h316:	data_out=16'h0;
17'h317:	data_out=16'h0;
17'h318:	data_out=16'h0;
17'h319:	data_out=16'h0;
17'h31a:	data_out=16'h0;
17'h31b:	data_out=16'h0;
17'h31c:	data_out=16'h0;
17'h31d:	data_out=16'h0;
17'h31e:	data_out=16'h0;
17'h31f:	data_out=16'h0;
17'h320:	data_out=16'h0;
17'h321:	data_out=16'h0;
17'h322:	data_out=16'h0;
17'h323:	data_out=16'h0;
17'h324:	data_out=16'h0;
17'h325:	data_out=16'h0;
17'h326:	data_out=16'h0;
17'h327:	data_out=16'h0;
17'h328:	data_out=16'h0;
17'h329:	data_out=16'h0;
17'h32a:	data_out=16'h0;
17'h32b:	data_out=16'h0;
17'h32c:	data_out=16'h0;
17'h32d:	data_out=16'h0;
17'h32e:	data_out=16'h0;
17'h32f:	data_out=16'h0;
17'h330:	data_out=16'h0;
17'h331:	data_out=16'h0;
17'h332:	data_out=16'h0;
17'h333:	data_out=16'h0;
17'h334:	data_out=16'h0;
17'h335:	data_out=16'h0;
17'h336:	data_out=16'h0;
17'h337:	data_out=16'h0;
17'h338:	data_out=16'h0;
17'h339:	data_out=16'h0;
17'h33a:	data_out=16'h0;
17'h33b:	data_out=16'h0;
17'h33c:	data_out=16'h0;
17'h33d:	data_out=16'h0;
17'h33e:	data_out=16'h0;
17'h33f:	data_out=16'h0;
17'h340:	data_out=16'h0;
17'h341:	data_out=16'h0;
17'h342:	data_out=16'h0;
17'h343:	data_out=16'h0;
17'h344:	data_out=16'h0;
17'h345:	data_out=16'h0;
17'h346:	data_out=16'h0;
17'h347:	data_out=16'h0;
17'h348:	data_out=16'h0;
17'h349:	data_out=16'h0;
17'h34a:	data_out=16'h0;
17'h34b:	data_out=16'h0;
17'h34c:	data_out=16'h0;
17'h34d:	data_out=16'h0;
17'h34e:	data_out=16'h0;
17'h34f:	data_out=16'h0;
17'h350:	data_out=16'h0;
17'h351:	data_out=16'h0;
17'h352:	data_out=16'h0;
17'h353:	data_out=16'h0;
17'h354:	data_out=16'h0;
17'h355:	data_out=16'h0;
17'h356:	data_out=16'h0;
17'h357:	data_out=16'h0;
17'h358:	data_out=16'h0;
17'h359:	data_out=16'h0;
17'h35a:	data_out=16'h0;
17'h35b:	data_out=16'h0;
17'h35c:	data_out=16'h0;
17'h35d:	data_out=16'h0;
17'h35e:	data_out=16'h0;
17'h35f:	data_out=16'h0;
17'h360:	data_out=16'h0;
17'h361:	data_out=16'h0;
17'h362:	data_out=16'h0;
17'h363:	data_out=16'h0;
17'h364:	data_out=16'h0;
17'h365:	data_out=16'h0;
17'h366:	data_out=16'h0;
17'h367:	data_out=16'h0;
17'h368:	data_out=16'h0;
17'h369:	data_out=16'h0;
17'h36a:	data_out=16'h0;
17'h36b:	data_out=16'h0;
17'h36c:	data_out=16'h0;
17'h36d:	data_out=16'h0;
17'h36e:	data_out=16'h0;
17'h36f:	data_out=16'h0;
17'h370:	data_out=16'h0;
17'h371:	data_out=16'h0;
17'h372:	data_out=16'h0;
17'h373:	data_out=16'h0;
17'h374:	data_out=16'h0;
17'h375:	data_out=16'h0;
17'h376:	data_out=16'h0;
17'h377:	data_out=16'h0;
17'h378:	data_out=16'h0;
17'h379:	data_out=16'h0;
17'h37a:	data_out=16'h0;
17'h37b:	data_out=16'h0;
17'h37c:	data_out=16'h0;
17'h37d:	data_out=16'h0;
17'h37e:	data_out=16'h0;
17'h37f:	data_out=16'h0;
17'h380:	data_out=16'h0;
17'h381:	data_out=16'h0;
17'h382:	data_out=16'h0;
17'h383:	data_out=16'h0;
17'h384:	data_out=16'h0;
17'h385:	data_out=16'h0;
17'h386:	data_out=16'h0;
17'h387:	data_out=16'h0;
17'h388:	data_out=16'h0;
17'h389:	data_out=16'h0;
17'h38a:	data_out=16'h0;
17'h38b:	data_out=16'h0;
17'h38c:	data_out=16'h0;
17'h38d:	data_out=16'h0;
17'h38e:	data_out=16'h0;
17'h38f:	data_out=16'h33;
17'h390:	data_out=16'ha0;
17'h391:	data_out=16'hfe;
17'h392:	data_out=16'ha0;
17'h393:	data_out=16'h32;
17'h394:	data_out=16'h0;
17'h395:	data_out=16'h0;
17'h396:	data_out=16'h0;
17'h397:	data_out=16'h0;
17'h398:	data_out=16'h0;
17'h399:	data_out=16'h0;
17'h39a:	data_out=16'h0;
17'h39b:	data_out=16'h0;
17'h39c:	data_out=16'h0;
17'h39d:	data_out=16'h0;
17'h39e:	data_out=16'h0;
17'h39f:	data_out=16'h0;
17'h3a0:	data_out=16'h0;
17'h3a1:	data_out=16'h0;
17'h3a2:	data_out=16'h0;
17'h3a3:	data_out=16'h0;
17'h3a4:	data_out=16'h0;
17'h3a5:	data_out=16'h0;
17'h3a6:	data_out=16'h0;
17'h3a7:	data_out=16'h0;
17'h3a8:	data_out=16'h0;
17'h3a9:	data_out=16'h0;
17'h3aa:	data_out=16'h30;
17'h3ab:	data_out=16'hef;
17'h3ac:	data_out=16'hfd;
17'h3ad:	data_out=16'hfd;
17'h3ae:	data_out=16'hfd;
17'h3af:	data_out=16'hee;
17'h3b0:	data_out=16'h0;
17'h3b1:	data_out=16'h0;
17'h3b2:	data_out=16'h0;
17'h3b3:	data_out=16'h0;
17'h3b4:	data_out=16'h0;
17'h3b5:	data_out=16'h0;
17'h3b6:	data_out=16'h0;
17'h3b7:	data_out=16'h0;
17'h3b8:	data_out=16'h0;
17'h3b9:	data_out=16'h0;
17'h3ba:	data_out=16'h0;
17'h3bb:	data_out=16'h0;
17'h3bc:	data_out=16'h0;
17'h3bd:	data_out=16'h0;
17'h3be:	data_out=16'h0;
17'h3bf:	data_out=16'h0;
17'h3c0:	data_out=16'h0;
17'h3c1:	data_out=16'h0;
17'h3c2:	data_out=16'h0;
17'h3c3:	data_out=16'h0;
17'h3c4:	data_out=16'h0;
17'h3c5:	data_out=16'h36;
17'h3c6:	data_out=16'he4;
17'h3c7:	data_out=16'hfe;
17'h3c8:	data_out=16'hfd;
17'h3c9:	data_out=16'hf0;
17'h3ca:	data_out=16'hea;
17'h3cb:	data_out=16'hfd;
17'h3cc:	data_out=16'h39;
17'h3cd:	data_out=16'h6;
17'h3ce:	data_out=16'h0;
17'h3cf:	data_out=16'h0;
17'h3d0:	data_out=16'h0;
17'h3d1:	data_out=16'h0;
17'h3d2:	data_out=16'h0;
17'h3d3:	data_out=16'h0;
17'h3d4:	data_out=16'h0;
17'h3d5:	data_out=16'h0;
17'h3d6:	data_out=16'h0;
17'h3d7:	data_out=16'h0;
17'h3d8:	data_out=16'h0;
17'h3d9:	data_out=16'h0;
17'h3da:	data_out=16'h0;
17'h3db:	data_out=16'h0;
17'h3dc:	data_out=16'h0;
17'h3dd:	data_out=16'h0;
17'h3de:	data_out=16'h0;
17'h3df:	data_out=16'ha;
17'h3e0:	data_out=16'h3c;
17'h3e1:	data_out=16'he1;
17'h3e2:	data_out=16'hfd;
17'h3e3:	data_out=16'hfe;
17'h3e4:	data_out=16'hfd;
17'h3e5:	data_out=16'hcb;
17'h3e6:	data_out=16'h54;
17'h3e7:	data_out=16'hfd;
17'h3e8:	data_out=16'hfe;
17'h3e9:	data_out=16'h7a;
17'h3ea:	data_out=16'h0;
17'h3eb:	data_out=16'h0;
17'h3ec:	data_out=16'h0;
17'h3ed:	data_out=16'h0;
17'h3ee:	data_out=16'h0;
17'h3ef:	data_out=16'h0;
17'h3f0:	data_out=16'h0;
17'h3f1:	data_out=16'h0;
17'h3f2:	data_out=16'h0;
17'h3f3:	data_out=16'h0;
17'h3f4:	data_out=16'h0;
17'h3f5:	data_out=16'h0;
17'h3f6:	data_out=16'h0;
17'h3f7:	data_out=16'h0;
17'h3f8:	data_out=16'h0;
17'h3f9:	data_out=16'h0;
17'h3fa:	data_out=16'h0;
17'h3fb:	data_out=16'ha4;
17'h3fc:	data_out=16'hfd;
17'h3fd:	data_out=16'hfd;
17'h3fe:	data_out=16'hfd;
17'h3ff:	data_out=16'hfe;
17'h400:	data_out=16'hfd;
17'h401:	data_out=16'hfd;
17'h402:	data_out=16'h60;
17'h403:	data_out=16'hbe;
17'h404:	data_out=16'hfe;
17'h405:	data_out=16'ha8;
17'h406:	data_out=16'h0;
17'h407:	data_out=16'h0;
17'h408:	data_out=16'h0;
17'h409:	data_out=16'h0;
17'h40a:	data_out=16'h0;
17'h40b:	data_out=16'h0;
17'h40c:	data_out=16'h0;
17'h40d:	data_out=16'h0;
17'h40e:	data_out=16'h0;
17'h40f:	data_out=16'h0;
17'h410:	data_out=16'h0;
17'h411:	data_out=16'h0;
17'h412:	data_out=16'h0;
17'h413:	data_out=16'h0;
17'h414:	data_out=16'h0;
17'h415:	data_out=16'h0;
17'h416:	data_out=16'h33;
17'h417:	data_out=16'hef;
17'h418:	data_out=16'hfe;
17'h419:	data_out=16'hfe;
17'h41a:	data_out=16'hbf;
17'h41b:	data_out=16'h72;
17'h41c:	data_out=16'hfe;
17'h41d:	data_out=16'he5;
17'h41e:	data_out=16'h2f;
17'h41f:	data_out=16'h4f;
17'h420:	data_out=16'h100;
17'h421:	data_out=16'ha9;
17'h422:	data_out=16'h0;
17'h423:	data_out=16'h0;
17'h424:	data_out=16'h0;
17'h425:	data_out=16'h0;
17'h426:	data_out=16'h0;
17'h427:	data_out=16'h0;
17'h428:	data_out=16'h0;
17'h429:	data_out=16'h0;
17'h42a:	data_out=16'h0;
17'h42b:	data_out=16'h0;
17'h42c:	data_out=16'h0;
17'h42d:	data_out=16'h0;
17'h42e:	data_out=16'h0;
17'h42f:	data_out=16'h0;
17'h430:	data_out=16'h0;
17'h431:	data_out=16'h30;
17'h432:	data_out=16'hef;
17'h433:	data_out=16'hfd;
17'h434:	data_out=16'hfd;
17'h435:	data_out=16'hb4;
17'h436:	data_out=16'hc;
17'h437:	data_out=16'h4b;
17'h438:	data_out=16'h79;
17'h439:	data_out=16'h15;
17'h43a:	data_out=16'h0;
17'h43b:	data_out=16'h0;
17'h43c:	data_out=16'hfe;
17'h43d:	data_out=16'hf4;
17'h43e:	data_out=16'h32;
17'h43f:	data_out=16'h0;
17'h440:	data_out=16'h0;
17'h441:	data_out=16'h0;
17'h442:	data_out=16'h0;
17'h443:	data_out=16'h0;
17'h444:	data_out=16'h0;
17'h445:	data_out=16'h0;
17'h446:	data_out=16'h0;
17'h447:	data_out=16'h0;
17'h448:	data_out=16'h0;
17'h449:	data_out=16'h0;
17'h44a:	data_out=16'h0;
17'h44b:	data_out=16'h0;
17'h44c:	data_out=16'h26;
17'h44d:	data_out=16'ha6;
17'h44e:	data_out=16'hfe;
17'h44f:	data_out=16'hea;
17'h450:	data_out=16'hd1;
17'h451:	data_out=16'h54;
17'h452:	data_out=16'h0;
17'h453:	data_out=16'h0;
17'h454:	data_out=16'h0;
17'h455:	data_out=16'h0;
17'h456:	data_out=16'h0;
17'h457:	data_out=16'h0;
17'h458:	data_out=16'hfe;
17'h459:	data_out=16'hfd;
17'h45a:	data_out=16'ha6;
17'h45b:	data_out=16'h0;
17'h45c:	data_out=16'h0;
17'h45d:	data_out=16'h0;
17'h45e:	data_out=16'h0;
17'h45f:	data_out=16'h0;
17'h460:	data_out=16'h0;
17'h461:	data_out=16'h0;
17'h462:	data_out=16'h0;
17'h463:	data_out=16'h0;
17'h464:	data_out=16'h0;
17'h465:	data_out=16'h0;
17'h466:	data_out=16'h0;
17'h467:	data_out=16'h7;
17'h468:	data_out=16'hb3;
17'h469:	data_out=16'hfd;
17'h46a:	data_out=16'hf1;
17'h46b:	data_out=16'h47;
17'h46c:	data_out=16'h13;
17'h46d:	data_out=16'h1c;
17'h46e:	data_out=16'h0;
17'h46f:	data_out=16'h0;
17'h470:	data_out=16'h0;
17'h471:	data_out=16'h0;
17'h472:	data_out=16'h0;
17'h473:	data_out=16'h0;
17'h474:	data_out=16'hfe;
17'h475:	data_out=16'hfd;
17'h476:	data_out=16'hc4;
17'h477:	data_out=16'h0;
17'h478:	data_out=16'h0;
17'h479:	data_out=16'h0;
17'h47a:	data_out=16'h0;
17'h47b:	data_out=16'h0;
17'h47c:	data_out=16'h0;
17'h47d:	data_out=16'h0;
17'h47e:	data_out=16'h0;
17'h47f:	data_out=16'h0;
17'h480:	data_out=16'h0;
17'h481:	data_out=16'h0;
17'h482:	data_out=16'h0;
17'h483:	data_out=16'h39;
17'h484:	data_out=16'hfd;
17'h485:	data_out=16'hfd;
17'h486:	data_out=16'h3f;
17'h487:	data_out=16'h0;
17'h488:	data_out=16'h0;
17'h489:	data_out=16'h0;
17'h48a:	data_out=16'h0;
17'h48b:	data_out=16'h0;
17'h48c:	data_out=16'h0;
17'h48d:	data_out=16'h0;
17'h48e:	data_out=16'h0;
17'h48f:	data_out=16'h0;
17'h490:	data_out=16'hfe;
17'h491:	data_out=16'hfd;
17'h492:	data_out=16'hc4;
17'h493:	data_out=16'h0;
17'h494:	data_out=16'h0;
17'h495:	data_out=16'h0;
17'h496:	data_out=16'h0;
17'h497:	data_out=16'h0;
17'h498:	data_out=16'h0;
17'h499:	data_out=16'h0;
17'h49a:	data_out=16'h0;
17'h49b:	data_out=16'h0;
17'h49c:	data_out=16'h0;
17'h49d:	data_out=16'h0;
17'h49e:	data_out=16'h0;
17'h49f:	data_out=16'hc7;
17'h4a0:	data_out=16'hfe;
17'h4a1:	data_out=16'hbf;
17'h4a2:	data_out=16'h0;
17'h4a3:	data_out=16'h0;
17'h4a4:	data_out=16'h0;
17'h4a5:	data_out=16'h0;
17'h4a6:	data_out=16'h0;
17'h4a7:	data_out=16'h0;
17'h4a8:	data_out=16'h0;
17'h4a9:	data_out=16'h0;
17'h4aa:	data_out=16'h0;
17'h4ab:	data_out=16'h0;
17'h4ac:	data_out=16'h100;
17'h4ad:	data_out=16'hfe;
17'h4ae:	data_out=16'hc5;
17'h4af:	data_out=16'h0;
17'h4b0:	data_out=16'h0;
17'h4b1:	data_out=16'h0;
17'h4b2:	data_out=16'h0;
17'h4b3:	data_out=16'h0;
17'h4b4:	data_out=16'h0;
17'h4b5:	data_out=16'h0;
17'h4b6:	data_out=16'h0;
17'h4b7:	data_out=16'h0;
17'h4b8:	data_out=16'h0;
17'h4b9:	data_out=16'h0;
17'h4ba:	data_out=16'h4c;
17'h4bb:	data_out=16'hf7;
17'h4bc:	data_out=16'hfd;
17'h4bd:	data_out=16'h70;
17'h4be:	data_out=16'h0;
17'h4bf:	data_out=16'h0;
17'h4c0:	data_out=16'h0;
17'h4c1:	data_out=16'h0;
17'h4c2:	data_out=16'h0;
17'h4c3:	data_out=16'h0;
17'h4c4:	data_out=16'h0;
17'h4c5:	data_out=16'h0;
17'h4c6:	data_out=16'h0;
17'h4c7:	data_out=16'h0;
17'h4c8:	data_out=16'hfe;
17'h4c9:	data_out=16'hfd;
17'h4ca:	data_out=16'h95;
17'h4cb:	data_out=16'h0;
17'h4cc:	data_out=16'h0;
17'h4cd:	data_out=16'h0;
17'h4ce:	data_out=16'h0;
17'h4cf:	data_out=16'h0;
17'h4d0:	data_out=16'h0;
17'h4d1:	data_out=16'h0;
17'h4d2:	data_out=16'h0;
17'h4d3:	data_out=16'h0;
17'h4d4:	data_out=16'h0;
17'h4d5:	data_out=16'h0;
17'h4d6:	data_out=16'h55;
17'h4d7:	data_out=16'hfd;
17'h4d8:	data_out=16'he7;
17'h4d9:	data_out=16'h19;
17'h4da:	data_out=16'h0;
17'h4db:	data_out=16'h0;
17'h4dc:	data_out=16'h0;
17'h4dd:	data_out=16'h0;
17'h4de:	data_out=16'h0;
17'h4df:	data_out=16'h0;
17'h4e0:	data_out=16'h0;
17'h4e1:	data_out=16'h0;
17'h4e2:	data_out=16'h7;
17'h4e3:	data_out=16'h88;
17'h4e4:	data_out=16'hfe;
17'h4e5:	data_out=16'hbb;
17'h4e6:	data_out=16'hc;
17'h4e7:	data_out=16'h0;
17'h4e8:	data_out=16'h0;
17'h4e9:	data_out=16'h0;
17'h4ea:	data_out=16'h0;
17'h4eb:	data_out=16'h0;
17'h4ec:	data_out=16'h0;
17'h4ed:	data_out=16'h0;
17'h4ee:	data_out=16'h0;
17'h4ef:	data_out=16'h0;
17'h4f0:	data_out=16'h0;
17'h4f1:	data_out=16'h0;
17'h4f2:	data_out=16'h55;
17'h4f3:	data_out=16'hfd;
17'h4f4:	data_out=16'he0;
17'h4f5:	data_out=16'h0;
17'h4f6:	data_out=16'h0;
17'h4f7:	data_out=16'h0;
17'h4f8:	data_out=16'h0;
17'h4f9:	data_out=16'h0;
17'h4fa:	data_out=16'h0;
17'h4fb:	data_out=16'h0;
17'h4fc:	data_out=16'h0;
17'h4fd:	data_out=16'h7;
17'h4fe:	data_out=16'h84;
17'h4ff:	data_out=16'hfd;
17'h500:	data_out=16'he2;
17'h501:	data_out=16'h47;
17'h502:	data_out=16'h0;
17'h503:	data_out=16'h0;
17'h504:	data_out=16'h0;
17'h505:	data_out=16'h0;
17'h506:	data_out=16'h0;
17'h507:	data_out=16'h0;
17'h508:	data_out=16'h0;
17'h509:	data_out=16'h0;
17'h50a:	data_out=16'h0;
17'h50b:	data_out=16'h0;
17'h50c:	data_out=16'h0;
17'h50d:	data_out=16'h0;
17'h50e:	data_out=16'h55;
17'h50f:	data_out=16'hfd;
17'h510:	data_out=16'h92;
17'h511:	data_out=16'h0;
17'h512:	data_out=16'h0;
17'h513:	data_out=16'h0;
17'h514:	data_out=16'h0;
17'h515:	data_out=16'h0;
17'h516:	data_out=16'h0;
17'h517:	data_out=16'h0;
17'h518:	data_out=16'h30;
17'h519:	data_out=16'ha6;
17'h51a:	data_out=16'hfd;
17'h51b:	data_out=16'hae;
17'h51c:	data_out=16'h0;
17'h51d:	data_out=16'h0;
17'h51e:	data_out=16'h0;
17'h51f:	data_out=16'h0;
17'h520:	data_out=16'h0;
17'h521:	data_out=16'h0;
17'h522:	data_out=16'h0;
17'h523:	data_out=16'h0;
17'h524:	data_out=16'h0;
17'h525:	data_out=16'h0;
17'h526:	data_out=16'h0;
17'h527:	data_out=16'h0;
17'h528:	data_out=16'h0;
17'h529:	data_out=16'h0;
17'h52a:	data_out=16'h56;
17'h52b:	data_out=16'hfe;
17'h52c:	data_out=16'he2;
17'h52d:	data_out=16'h0;
17'h52e:	data_out=16'h0;
17'h52f:	data_out=16'h0;
17'h530:	data_out=16'h0;
17'h531:	data_out=16'h0;
17'h532:	data_out=16'h0;
17'h533:	data_out=16'h72;
17'h534:	data_out=16'hef;
17'h535:	data_out=16'hfe;
17'h536:	data_out=16'ha3;
17'h537:	data_out=16'h0;
17'h538:	data_out=16'h0;
17'h539:	data_out=16'h0;
17'h53a:	data_out=16'h0;
17'h53b:	data_out=16'h0;
17'h53c:	data_out=16'h0;
17'h53d:	data_out=16'h0;
17'h53e:	data_out=16'h0;
17'h53f:	data_out=16'h0;
17'h540:	data_out=16'h0;
17'h541:	data_out=16'h0;
17'h542:	data_out=16'h0;
17'h543:	data_out=16'h0;
17'h544:	data_out=16'h0;
17'h545:	data_out=16'h0;
17'h546:	data_out=16'h55;
17'h547:	data_out=16'hfd;
17'h548:	data_out=16'hfa;
17'h549:	data_out=16'h93;
17'h54a:	data_out=16'h30;
17'h54b:	data_out=16'h1d;
17'h54c:	data_out=16'h55;
17'h54d:	data_out=16'hb3;
17'h54e:	data_out=16'he2;
17'h54f:	data_out=16'hfe;
17'h550:	data_out=16'he0;
17'h551:	data_out=16'ha8;
17'h552:	data_out=16'h38;
17'h553:	data_out=16'h0;
17'h554:	data_out=16'h0;
17'h555:	data_out=16'h0;
17'h556:	data_out=16'h0;
17'h557:	data_out=16'h0;
17'h558:	data_out=16'h0;
17'h559:	data_out=16'h0;
17'h55a:	data_out=16'h0;
17'h55b:	data_out=16'h0;
17'h55c:	data_out=16'h0;
17'h55d:	data_out=16'h0;
17'h55e:	data_out=16'h0;
17'h55f:	data_out=16'h0;
17'h560:	data_out=16'h0;
17'h561:	data_out=16'h0;
17'h562:	data_out=16'h55;
17'h563:	data_out=16'hfd;
17'h564:	data_out=16'hfd;
17'h565:	data_out=16'hfd;
17'h566:	data_out=16'he6;
17'h567:	data_out=16'hd8;
17'h568:	data_out=16'hfd;
17'h569:	data_out=16'hfd;
17'h56a:	data_out=16'hfd;
17'h56b:	data_out=16'hc5;
17'h56c:	data_out=16'h83;
17'h56d:	data_out=16'h0;
17'h56e:	data_out=16'h0;
17'h56f:	data_out=16'h0;
17'h570:	data_out=16'h0;
17'h571:	data_out=16'h0;
17'h572:	data_out=16'h0;
17'h573:	data_out=16'h0;
17'h574:	data_out=16'h0;
17'h575:	data_out=16'h0;
17'h576:	data_out=16'h0;
17'h577:	data_out=16'h0;
17'h578:	data_out=16'h0;
17'h579:	data_out=16'h0;
17'h57a:	data_out=16'h0;
17'h57b:	data_out=16'h0;
17'h57c:	data_out=16'h0;
17'h57d:	data_out=16'h0;
17'h57e:	data_out=16'h1c;
17'h57f:	data_out=16'hc8;
17'h580:	data_out=16'hfd;
17'h581:	data_out=16'hfd;
17'h582:	data_out=16'hfe;
17'h583:	data_out=16'hfd;
17'h584:	data_out=16'hfd;
17'h585:	data_out=16'hea;
17'h586:	data_out=16'h92;
17'h587:	data_out=16'h0;
17'h588:	data_out=16'h0;
17'h589:	data_out=16'h0;
17'h58a:	data_out=16'h0;
17'h58b:	data_out=16'h0;
17'h58c:	data_out=16'h0;
17'h58d:	data_out=16'h0;
17'h58e:	data_out=16'h0;
17'h58f:	data_out=16'h0;
17'h590:	data_out=16'h0;
17'h591:	data_out=16'h0;
17'h592:	data_out=16'h0;
17'h593:	data_out=16'h0;
17'h594:	data_out=16'h0;
17'h595:	data_out=16'h0;
17'h596:	data_out=16'h0;
17'h597:	data_out=16'h0;
17'h598:	data_out=16'h0;
17'h599:	data_out=16'h0;
17'h59a:	data_out=16'h0;
17'h59b:	data_out=16'h19;
17'h59c:	data_out=16'h81;
17'h59d:	data_out=16'hfd;
17'h59e:	data_out=16'hfe;
17'h59f:	data_out=16'hfd;
17'h5a0:	data_out=16'h8e;
17'h5a1:	data_out=16'h25;
17'h5a2:	data_out=16'h0;
17'h5a3:	data_out=16'h0;
17'h5a4:	data_out=16'h0;
17'h5a5:	data_out=16'h0;
17'h5a6:	data_out=16'h0;
17'h5a7:	data_out=16'h0;
17'h5a8:	data_out=16'h0;
17'h5a9:	data_out=16'h0;
17'h5aa:	data_out=16'h0;
17'h5ab:	data_out=16'h0;
17'h5ac:	data_out=16'h0;
17'h5ad:	data_out=16'h0;
17'h5ae:	data_out=16'h0;
17'h5af:	data_out=16'h0;
17'h5b0:	data_out=16'h0;
17'h5b1:	data_out=16'h0;
17'h5b2:	data_out=16'h0;
17'h5b3:	data_out=16'h0;
17'h5b4:	data_out=16'h0;
17'h5b5:	data_out=16'h0;
17'h5b6:	data_out=16'h0;
17'h5b7:	data_out=16'h0;
17'h5b8:	data_out=16'h0;
17'h5b9:	data_out=16'h0;
17'h5ba:	data_out=16'h0;
17'h5bb:	data_out=16'h0;
17'h5bc:	data_out=16'h0;
17'h5bd:	data_out=16'h0;
17'h5be:	data_out=16'h0;
17'h5bf:	data_out=16'h0;
17'h5c0:	data_out=16'h0;
17'h5c1:	data_out=16'h0;
17'h5c2:	data_out=16'h0;
17'h5c3:	data_out=16'h0;
17'h5c4:	data_out=16'h0;
17'h5c5:	data_out=16'h0;
17'h5c6:	data_out=16'h0;
17'h5c7:	data_out=16'h0;
17'h5c8:	data_out=16'h0;
17'h5c9:	data_out=16'h0;
17'h5ca:	data_out=16'h0;
17'h5cb:	data_out=16'h0;
17'h5cc:	data_out=16'h0;
17'h5cd:	data_out=16'h0;
17'h5ce:	data_out=16'h0;
17'h5cf:	data_out=16'h0;
17'h5d0:	data_out=16'h0;
17'h5d1:	data_out=16'h0;
17'h5d2:	data_out=16'h0;
17'h5d3:	data_out=16'h0;
17'h5d4:	data_out=16'h0;
17'h5d5:	data_out=16'h0;
17'h5d6:	data_out=16'h0;
17'h5d7:	data_out=16'h0;
17'h5d8:	data_out=16'h0;
17'h5d9:	data_out=16'h0;
17'h5da:	data_out=16'h0;
17'h5db:	data_out=16'h0;
17'h5dc:	data_out=16'h0;
17'h5dd:	data_out=16'h0;
17'h5de:	data_out=16'h0;
17'h5df:	data_out=16'h0;
17'h5e0:	data_out=16'h0;
17'h5e1:	data_out=16'h0;
17'h5e2:	data_out=16'h0;
17'h5e3:	data_out=16'h0;
17'h5e4:	data_out=16'h0;
17'h5e5:	data_out=16'h0;
17'h5e6:	data_out=16'h0;
17'h5e7:	data_out=16'h0;
17'h5e8:	data_out=16'h0;
17'h5e9:	data_out=16'h0;
17'h5ea:	data_out=16'h0;
17'h5eb:	data_out=16'h0;
17'h5ec:	data_out=16'h0;
17'h5ed:	data_out=16'h0;
17'h5ee:	data_out=16'h0;
17'h5ef:	data_out=16'h0;
17'h5f0:	data_out=16'h0;
17'h5f1:	data_out=16'h0;
17'h5f2:	data_out=16'h0;
17'h5f3:	data_out=16'h0;
17'h5f4:	data_out=16'h0;
17'h5f5:	data_out=16'h0;
17'h5f6:	data_out=16'h0;
17'h5f7:	data_out=16'h0;
17'h5f8:	data_out=16'h0;
17'h5f9:	data_out=16'h0;
17'h5fa:	data_out=16'h0;
17'h5fb:	data_out=16'h0;
17'h5fc:	data_out=16'h0;
17'h5fd:	data_out=16'h0;
17'h5fe:	data_out=16'h0;
17'h5ff:	data_out=16'h0;
17'h600:	data_out=16'h0;
17'h601:	data_out=16'h0;
17'h602:	data_out=16'h0;
17'h603:	data_out=16'h0;
17'h604:	data_out=16'h0;
17'h605:	data_out=16'h0;
17'h606:	data_out=16'h0;
17'h607:	data_out=16'h0;
17'h608:	data_out=16'h0;
17'h609:	data_out=16'h0;
17'h60a:	data_out=16'h0;
17'h60b:	data_out=16'h0;
17'h60c:	data_out=16'h0;
17'h60d:	data_out=16'h0;
17'h60e:	data_out=16'h0;
17'h60f:	data_out=16'h0;
17'h610:	data_out=16'h0;
17'h611:	data_out=16'h0;
17'h612:	data_out=16'h0;
17'h613:	data_out=16'h0;
17'h614:	data_out=16'h0;
17'h615:	data_out=16'h0;
17'h616:	data_out=16'h0;
17'h617:	data_out=16'h0;
17'h618:	data_out=16'h0;
17'h619:	data_out=16'h0;
17'h61a:	data_out=16'h0;
17'h61b:	data_out=16'h0;
17'h61c:	data_out=16'h0;
17'h61d:	data_out=16'h0;
17'h61e:	data_out=16'h0;
17'h61f:	data_out=16'h0;
17'h620:	data_out=16'h0;
17'h621:	data_out=16'h0;
17'h622:	data_out=16'h0;
17'h623:	data_out=16'h0;
17'h624:	data_out=16'h0;
17'h625:	data_out=16'h0;
17'h626:	data_out=16'h0;
17'h627:	data_out=16'h0;
17'h628:	data_out=16'h0;
17'h629:	data_out=16'h0;
17'h62a:	data_out=16'h0;
17'h62b:	data_out=16'h0;
17'h62c:	data_out=16'h0;
17'h62d:	data_out=16'h0;
17'h62e:	data_out=16'h0;
17'h62f:	data_out=16'h0;
17'h630:	data_out=16'h0;
17'h631:	data_out=16'h0;
17'h632:	data_out=16'h0;
17'h633:	data_out=16'h0;
17'h634:	data_out=16'h0;
17'h635:	data_out=16'h0;
17'h636:	data_out=16'h0;
17'h637:	data_out=16'h0;
17'h638:	data_out=16'h0;
17'h639:	data_out=16'h0;
17'h63a:	data_out=16'h0;
17'h63b:	data_out=16'h0;
17'h63c:	data_out=16'h0;
17'h63d:	data_out=16'h0;
17'h63e:	data_out=16'h0;
17'h63f:	data_out=16'h0;
17'h640:	data_out=16'h0;
17'h641:	data_out=16'h0;
17'h642:	data_out=16'h0;
17'h643:	data_out=16'h0;
17'h644:	data_out=16'h0;
17'h645:	data_out=16'h0;
17'h646:	data_out=16'h0;
17'h647:	data_out=16'h0;
17'h648:	data_out=16'h0;
17'h649:	data_out=16'h0;
17'h64a:	data_out=16'h0;
17'h64b:	data_out=16'h0;
17'h64c:	data_out=16'h0;
17'h64d:	data_out=16'h0;
17'h64e:	data_out=16'h0;
17'h64f:	data_out=16'h0;
17'h650:	data_out=16'h0;
17'h651:	data_out=16'h0;
17'h652:	data_out=16'h0;
17'h653:	data_out=16'h0;
17'h654:	data_out=16'h0;
17'h655:	data_out=16'h0;
17'h656:	data_out=16'h0;
17'h657:	data_out=16'h0;
17'h658:	data_out=16'h0;
17'h659:	data_out=16'h0;
17'h65a:	data_out=16'h0;
17'h65b:	data_out=16'h0;
17'h65c:	data_out=16'h0;
17'h65d:	data_out=16'h0;
17'h65e:	data_out=16'h0;
17'h65f:	data_out=16'h0;
17'h660:	data_out=16'h0;
17'h661:	data_out=16'h0;
17'h662:	data_out=16'h0;
17'h663:	data_out=16'h0;
17'h664:	data_out=16'h0;
17'h665:	data_out=16'h0;
17'h666:	data_out=16'h0;
17'h667:	data_out=16'h0;
17'h668:	data_out=16'h0;
17'h669:	data_out=16'h0;
17'h66a:	data_out=16'h0;
17'h66b:	data_out=16'h0;
17'h66c:	data_out=16'h0;
17'h66d:	data_out=16'h0;
17'h66e:	data_out=16'h0;
17'h66f:	data_out=16'h0;
17'h670:	data_out=16'h0;
17'h671:	data_out=16'h0;
17'h672:	data_out=16'h0;
17'h673:	data_out=16'h0;
17'h674:	data_out=16'h0;
17'h675:	data_out=16'h0;
17'h676:	data_out=16'h0;
17'h677:	data_out=16'h0;
17'h678:	data_out=16'h0;
17'h679:	data_out=16'h0;
17'h67a:	data_out=16'h0;
17'h67b:	data_out=16'h0;
17'h67c:	data_out=16'h0;
17'h67d:	data_out=16'h0;
17'h67e:	data_out=16'h0;
17'h67f:	data_out=16'h0;
17'h680:	data_out=16'h0;
17'h681:	data_out=16'h0;
17'h682:	data_out=16'h0;
17'h683:	data_out=16'h0;
17'h684:	data_out=16'h0;
17'h685:	data_out=16'h0;
17'h686:	data_out=16'h0;
17'h687:	data_out=16'h0;
17'h688:	data_out=16'h0;
17'h689:	data_out=16'h0;
17'h68a:	data_out=16'h0;
17'h68b:	data_out=16'h0;
17'h68c:	data_out=16'h0;
17'h68d:	data_out=16'h0;
17'h68e:	data_out=16'h0;
17'h68f:	data_out=16'h0;
17'h690:	data_out=16'h0;
17'h691:	data_out=16'h0;
17'h692:	data_out=16'h0;
17'h693:	data_out=16'h0;
17'h694:	data_out=16'h0;
17'h695:	data_out=16'h0;
17'h696:	data_out=16'h0;
17'h697:	data_out=16'h0;
17'h698:	data_out=16'h0;
17'h699:	data_out=16'h0;
17'h69a:	data_out=16'h0;
17'h69b:	data_out=16'h0;
17'h69c:	data_out=16'h0;
17'h69d:	data_out=16'h0;
17'h69e:	data_out=16'h0;
17'h69f:	data_out=16'h0;
17'h6a0:	data_out=16'h0;
17'h6a1:	data_out=16'h0;
17'h6a2:	data_out=16'h0;
17'h6a3:	data_out=16'h0;
17'h6a4:	data_out=16'h0;
17'h6a5:	data_out=16'h0;
17'h6a6:	data_out=16'h0;
17'h6a7:	data_out=16'h0;
17'h6a8:	data_out=16'h0;
17'h6a9:	data_out=16'h0;
17'h6aa:	data_out=16'h0;
17'h6ab:	data_out=16'h0;
17'h6ac:	data_out=16'h0;
17'h6ad:	data_out=16'h0;
17'h6ae:	data_out=16'h0;
17'h6af:	data_out=16'h0;
17'h6b0:	data_out=16'h0;
17'h6b1:	data_out=16'h0;
17'h6b2:	data_out=16'h0;
17'h6b3:	data_out=16'h0;
17'h6b4:	data_out=16'h0;
17'h6b5:	data_out=16'h0;
17'h6b6:	data_out=16'h0;
17'h6b7:	data_out=16'h0;
17'h6b8:	data_out=16'h0;
17'h6b9:	data_out=16'h0;
17'h6ba:	data_out=16'h0;
17'h6bb:	data_out=16'h0;
17'h6bc:	data_out=16'h0;
17'h6bd:	data_out=16'h0;
17'h6be:	data_out=16'h0;
17'h6bf:	data_out=16'h0;
17'h6c0:	data_out=16'h43;
17'h6c1:	data_out=16'he9;
17'h6c2:	data_out=16'h27;
17'h6c3:	data_out=16'h0;
17'h6c4:	data_out=16'h0;
17'h6c5:	data_out=16'h0;
17'h6c6:	data_out=16'h0;
17'h6c7:	data_out=16'h0;
17'h6c8:	data_out=16'h0;
17'h6c9:	data_out=16'h0;
17'h6ca:	data_out=16'h0;
17'h6cb:	data_out=16'h0;
17'h6cc:	data_out=16'h3e;
17'h6cd:	data_out=16'h51;
17'h6ce:	data_out=16'h0;
17'h6cf:	data_out=16'h0;
17'h6d0:	data_out=16'h0;
17'h6d1:	data_out=16'h0;
17'h6d2:	data_out=16'h0;
17'h6d3:	data_out=16'h0;
17'h6d4:	data_out=16'h0;
17'h6d5:	data_out=16'h0;
17'h6d6:	data_out=16'h0;
17'h6d7:	data_out=16'h0;
17'h6d8:	data_out=16'h0;
17'h6d9:	data_out=16'h0;
17'h6da:	data_out=16'h0;
17'h6db:	data_out=16'h0;
17'h6dc:	data_out=16'h78;
17'h6dd:	data_out=16'hb5;
17'h6de:	data_out=16'h27;
17'h6df:	data_out=16'h0;
17'h6e0:	data_out=16'h0;
17'h6e1:	data_out=16'h0;
17'h6e2:	data_out=16'h0;
17'h6e3:	data_out=16'h0;
17'h6e4:	data_out=16'h0;
17'h6e5:	data_out=16'h0;
17'h6e6:	data_out=16'h0;
17'h6e7:	data_out=16'h0;
17'h6e8:	data_out=16'h7e;
17'h6e9:	data_out=16'ha4;
17'h6ea:	data_out=16'h0;
17'h6eb:	data_out=16'h0;
17'h6ec:	data_out=16'h0;
17'h6ed:	data_out=16'h0;
17'h6ee:	data_out=16'h0;
17'h6ef:	data_out=16'h0;
17'h6f0:	data_out=16'h0;
17'h6f1:	data_out=16'h0;
17'h6f2:	data_out=16'h0;
17'h6f3:	data_out=16'h0;
17'h6f4:	data_out=16'h0;
17'h6f5:	data_out=16'h0;
17'h6f6:	data_out=16'h0;
17'h6f7:	data_out=16'h2;
17'h6f8:	data_out=16'h9a;
17'h6f9:	data_out=16'hd3;
17'h6fa:	data_out=16'h28;
17'h6fb:	data_out=16'h0;
17'h6fc:	data_out=16'h0;
17'h6fd:	data_out=16'h0;
17'h6fe:	data_out=16'h0;
17'h6ff:	data_out=16'h0;
17'h700:	data_out=16'h0;
17'h701:	data_out=16'h0;
17'h702:	data_out=16'h0;
17'h703:	data_out=16'h0;
17'h704:	data_out=16'hdd;
17'h705:	data_out=16'ha4;
17'h706:	data_out=16'h0;
17'h707:	data_out=16'h0;
17'h708:	data_out=16'h0;
17'h709:	data_out=16'h0;
17'h70a:	data_out=16'h0;
17'h70b:	data_out=16'h0;
17'h70c:	data_out=16'h0;
17'h70d:	data_out=16'h0;
17'h70e:	data_out=16'h0;
17'h70f:	data_out=16'h0;
17'h710:	data_out=16'h0;
17'h711:	data_out=16'h0;
17'h712:	data_out=16'h0;
17'h713:	data_out=16'h1b;
17'h714:	data_out=16'hff;
17'h715:	data_out=16'ha3;
17'h716:	data_out=16'h0;
17'h717:	data_out=16'h0;
17'h718:	data_out=16'h0;
17'h719:	data_out=16'h0;
17'h71a:	data_out=16'h0;
17'h71b:	data_out=16'h0;
17'h71c:	data_out=16'h0;
17'h71d:	data_out=16'h0;
17'h71e:	data_out=16'h0;
17'h71f:	data_out=16'h0;
17'h720:	data_out=16'hdf;
17'h721:	data_out=16'ha4;
17'h722:	data_out=16'h0;
17'h723:	data_out=16'h0;
17'h724:	data_out=16'h0;
17'h725:	data_out=16'h0;
17'h726:	data_out=16'h0;
17'h727:	data_out=16'h0;
17'h728:	data_out=16'h0;
17'h729:	data_out=16'h0;
17'h72a:	data_out=16'h0;
17'h72b:	data_out=16'h0;
17'h72c:	data_out=16'h0;
17'h72d:	data_out=16'h0;
17'h72e:	data_out=16'h0;
17'h72f:	data_out=16'hb8;
17'h730:	data_out=16'hff;
17'h731:	data_out=16'h7d;
17'h732:	data_out=16'h0;
17'h733:	data_out=16'h0;
17'h734:	data_out=16'h0;
17'h735:	data_out=16'h0;
17'h736:	data_out=16'h0;
17'h737:	data_out=16'h0;
17'h738:	data_out=16'h0;
17'h739:	data_out=16'h0;
17'h73a:	data_out=16'h0;
17'h73b:	data_out=16'h2e;
17'h73c:	data_out=16'hf6;
17'h73d:	data_out=16'ha4;
17'h73e:	data_out=16'h0;
17'h73f:	data_out=16'h0;
17'h740:	data_out=16'h0;
17'h741:	data_out=16'h0;
17'h742:	data_out=16'h0;
17'h743:	data_out=16'h0;
17'h744:	data_out=16'h0;
17'h745:	data_out=16'h0;
17'h746:	data_out=16'h0;
17'h747:	data_out=16'h0;
17'h748:	data_out=16'h0;
17'h749:	data_out=16'h0;
17'h74a:	data_out=16'h0;
17'h74b:	data_out=16'hc7;
17'h74c:	data_out=16'hff;
17'h74d:	data_out=16'h38;
17'h74e:	data_out=16'h0;
17'h74f:	data_out=16'h0;
17'h750:	data_out=16'h0;
17'h751:	data_out=16'h0;
17'h752:	data_out=16'h0;
17'h753:	data_out=16'h0;
17'h754:	data_out=16'h0;
17'h755:	data_out=16'h0;
17'h756:	data_out=16'h0;
17'h757:	data_out=16'h78;
17'h758:	data_out=16'hff;
17'h759:	data_out=16'ha4;
17'h75a:	data_out=16'h0;
17'h75b:	data_out=16'h0;
17'h75c:	data_out=16'h0;
17'h75d:	data_out=16'h0;
17'h75e:	data_out=16'h0;
17'h75f:	data_out=16'h0;
17'h760:	data_out=16'h0;
17'h761:	data_out=16'h0;
17'h762:	data_out=16'h0;
17'h763:	data_out=16'h0;
17'h764:	data_out=16'h0;
17'h765:	data_out=16'h0;
17'h766:	data_out=16'h17;
17'h767:	data_out=16'he8;
17'h768:	data_out=16'hff;
17'h769:	data_out=16'h1d;
17'h76a:	data_out=16'h0;
17'h76b:	data_out=16'h0;
17'h76c:	data_out=16'h0;
17'h76d:	data_out=16'h0;
17'h76e:	data_out=16'h0;
17'h76f:	data_out=16'h0;
17'h770:	data_out=16'h0;
17'h771:	data_out=16'h0;
17'h772:	data_out=16'h0;
17'h773:	data_out=16'ha0;
17'h774:	data_out=16'hff;
17'h775:	data_out=16'h78;
17'h776:	data_out=16'h0;
17'h777:	data_out=16'h0;
17'h778:	data_out=16'h0;
17'h779:	data_out=16'h0;
17'h77a:	data_out=16'h0;
17'h77b:	data_out=16'h0;
17'h77c:	data_out=16'h0;
17'h77d:	data_out=16'h0;
17'h77e:	data_out=16'h0;
17'h77f:	data_out=16'h0;
17'h780:	data_out=16'h0;
17'h781:	data_out=16'h0;
17'h782:	data_out=16'ha4;
17'h783:	data_out=16'hff;
17'h784:	data_out=16'hd9;
17'h785:	data_out=16'h10;
17'h786:	data_out=16'h0;
17'h787:	data_out=16'h0;
17'h788:	data_out=16'h0;
17'h789:	data_out=16'h0;
17'h78a:	data_out=16'h0;
17'h78b:	data_out=16'h0;
17'h78c:	data_out=16'h0;
17'h78d:	data_out=16'h0;
17'h78e:	data_out=16'h0;
17'h78f:	data_out=16'ha0;
17'h790:	data_out=16'hff;
17'h791:	data_out=16'h43;
17'h792:	data_out=16'h0;
17'h793:	data_out=16'h0;
17'h794:	data_out=16'h0;
17'h795:	data_out=16'h0;
17'h796:	data_out=16'h0;
17'h797:	data_out=16'h0;
17'h798:	data_out=16'h0;
17'h799:	data_out=16'h0;
17'h79a:	data_out=16'h0;
17'h79b:	data_out=16'he;
17'h79c:	data_out=16'h56;
17'h79d:	data_out=16'hb3;
17'h79e:	data_out=16'hf9;
17'h79f:	data_out=16'hff;
17'h7a0:	data_out=16'h5b;
17'h7a1:	data_out=16'h0;
17'h7a2:	data_out=16'h0;
17'h7a3:	data_out=16'h0;
17'h7a4:	data_out=16'h0;
17'h7a5:	data_out=16'h0;
17'h7a6:	data_out=16'h0;
17'h7a7:	data_out=16'h0;
17'h7a8:	data_out=16'h0;
17'h7a9:	data_out=16'h0;
17'h7aa:	data_out=16'h0;
17'h7ab:	data_out=16'ha0;
17'h7ac:	data_out=16'hff;
17'h7ad:	data_out=16'h55;
17'h7ae:	data_out=16'h0;
17'h7af:	data_out=16'h0;
17'h7b0:	data_out=16'h0;
17'h7b1:	data_out=16'h2f;
17'h7b2:	data_out=16'h31;
17'h7b3:	data_out=16'h74;
17'h7b4:	data_out=16'h91;
17'h7b5:	data_out=16'h97;
17'h7b6:	data_out=16'hf2;
17'h7b7:	data_out=16'hf4;
17'h7b8:	data_out=16'heb;
17'h7b9:	data_out=16'hb4;
17'h7ba:	data_out=16'hf2;
17'h7bb:	data_out=16'hfd;
17'h7bc:	data_out=16'h28;
17'h7bd:	data_out=16'h0;
17'h7be:	data_out=16'h0;
17'h7bf:	data_out=16'h0;
17'h7c0:	data_out=16'h0;
17'h7c1:	data_out=16'h0;
17'h7c2:	data_out=16'h0;
17'h7c3:	data_out=16'h0;
17'h7c4:	data_out=16'h0;
17'h7c5:	data_out=16'h0;
17'h7c6:	data_out=16'h0;
17'h7c7:	data_out=16'h97;
17'h7c8:	data_out=16'hfe;
17'h7c9:	data_out=16'hee;
17'h7ca:	data_out=16'hd0;
17'h7cb:	data_out=16'hd0;
17'h7cc:	data_out=16'hd0;
17'h7cd:	data_out=16'hfe;
17'h7ce:	data_out=16'hff;
17'h7cf:	data_out=16'hfb;
17'h7d0:	data_out=16'hf1;
17'h7d1:	data_out=16'hc7;
17'h7d2:	data_out=16'h90;
17'h7d3:	data_out=16'h5b;
17'h7d4:	data_out=16'h1c;
17'h7d5:	data_out=16'h5;
17'h7d6:	data_out=16'hea;
17'h7d7:	data_out=16'hfb;
17'h7d8:	data_out=16'h0;
17'h7d9:	data_out=16'h0;
17'h7da:	data_out=16'h0;
17'h7db:	data_out=16'h0;
17'h7dc:	data_out=16'h0;
17'h7dd:	data_out=16'h0;
17'h7de:	data_out=16'h0;
17'h7df:	data_out=16'h0;
17'h7e0:	data_out=16'h0;
17'h7e1:	data_out=16'h0;
17'h7e2:	data_out=16'h0;
17'h7e3:	data_out=16'h0;
17'h7e4:	data_out=16'h77;
17'h7e5:	data_out=16'hb2;
17'h7e6:	data_out=16'hb2;
17'h7e7:	data_out=16'hb2;
17'h7e8:	data_out=16'hb2;
17'h7e9:	data_out=16'hb2;
17'h7ea:	data_out=16'h62;
17'h7eb:	data_out=16'h38;
17'h7ec:	data_out=16'h0;
17'h7ed:	data_out=16'h0;
17'h7ee:	data_out=16'h0;
17'h7ef:	data_out=16'h0;
17'h7f0:	data_out=16'h0;
17'h7f1:	data_out=16'h66;
17'h7f2:	data_out=16'hff;
17'h7f3:	data_out=16'hdd;
17'h7f4:	data_out=16'h0;
17'h7f5:	data_out=16'h0;
17'h7f6:	data_out=16'h0;
17'h7f7:	data_out=16'h0;
17'h7f8:	data_out=16'h0;
17'h7f9:	data_out=16'h0;
17'h7fa:	data_out=16'h0;
17'h7fb:	data_out=16'h0;
17'h7fc:	data_out=16'h0;
17'h7fd:	data_out=16'h0;
17'h7fe:	data_out=16'h0;
17'h7ff:	data_out=16'h0;
17'h800:	data_out=16'h0;
17'h801:	data_out=16'h0;
17'h802:	data_out=16'h0;
17'h803:	data_out=16'h0;
17'h804:	data_out=16'h0;
17'h805:	data_out=16'h0;
17'h806:	data_out=16'h0;
17'h807:	data_out=16'h0;
17'h808:	data_out=16'h0;
17'h809:	data_out=16'h0;
17'h80a:	data_out=16'h0;
17'h80b:	data_out=16'h0;
17'h80c:	data_out=16'h0;
17'h80d:	data_out=16'haa;
17'h80e:	data_out=16'hff;
17'h80f:	data_out=16'h8a;
17'h810:	data_out=16'h0;
17'h811:	data_out=16'h0;
17'h812:	data_out=16'h0;
17'h813:	data_out=16'h0;
17'h814:	data_out=16'h0;
17'h815:	data_out=16'h0;
17'h816:	data_out=16'h0;
17'h817:	data_out=16'h0;
17'h818:	data_out=16'h0;
17'h819:	data_out=16'h0;
17'h81a:	data_out=16'h0;
17'h81b:	data_out=16'h0;
17'h81c:	data_out=16'h0;
17'h81d:	data_out=16'h0;
17'h81e:	data_out=16'h0;
17'h81f:	data_out=16'h0;
17'h820:	data_out=16'h0;
17'h821:	data_out=16'h0;
17'h822:	data_out=16'h0;
17'h823:	data_out=16'h0;
17'h824:	data_out=16'h0;
17'h825:	data_out=16'h0;
17'h826:	data_out=16'h0;
17'h827:	data_out=16'h0;
17'h828:	data_out=16'h0;
17'h829:	data_out=16'haa;
17'h82a:	data_out=16'hff;
17'h82b:	data_out=16'h39;
17'h82c:	data_out=16'h0;
17'h82d:	data_out=16'h0;
17'h82e:	data_out=16'h0;
17'h82f:	data_out=16'h0;
17'h830:	data_out=16'h0;
17'h831:	data_out=16'h0;
17'h832:	data_out=16'h0;
17'h833:	data_out=16'h0;
17'h834:	data_out=16'h0;
17'h835:	data_out=16'h0;
17'h836:	data_out=16'h0;
17'h837:	data_out=16'h0;
17'h838:	data_out=16'h0;
17'h839:	data_out=16'h0;
17'h83a:	data_out=16'h0;
17'h83b:	data_out=16'h0;
17'h83c:	data_out=16'h0;
17'h83d:	data_out=16'h0;
17'h83e:	data_out=16'h0;
17'h83f:	data_out=16'h0;
17'h840:	data_out=16'h0;
17'h841:	data_out=16'h0;
17'h842:	data_out=16'h0;
17'h843:	data_out=16'h0;
17'h844:	data_out=16'h0;
17'h845:	data_out=16'haa;
17'h846:	data_out=16'hff;
17'h847:	data_out=16'h39;
17'h848:	data_out=16'h0;
17'h849:	data_out=16'h0;
17'h84a:	data_out=16'h0;
17'h84b:	data_out=16'h0;
17'h84c:	data_out=16'h0;
17'h84d:	data_out=16'h0;
17'h84e:	data_out=16'h0;
17'h84f:	data_out=16'h0;
17'h850:	data_out=16'h0;
17'h851:	data_out=16'h0;
17'h852:	data_out=16'h0;
17'h853:	data_out=16'h0;
17'h854:	data_out=16'h0;
17'h855:	data_out=16'h0;
17'h856:	data_out=16'h0;
17'h857:	data_out=16'h0;
17'h858:	data_out=16'h0;
17'h859:	data_out=16'h0;
17'h85a:	data_out=16'h0;
17'h85b:	data_out=16'h0;
17'h85c:	data_out=16'h0;
17'h85d:	data_out=16'h0;
17'h85e:	data_out=16'h0;
17'h85f:	data_out=16'h0;
17'h860:	data_out=16'h0;
17'h861:	data_out=16'haa;
17'h862:	data_out=16'h100;
17'h863:	data_out=16'h5e;
17'h864:	data_out=16'h0;
17'h865:	data_out=16'h0;
17'h866:	data_out=16'h0;
17'h867:	data_out=16'h0;
17'h868:	data_out=16'h0;
17'h869:	data_out=16'h0;
17'h86a:	data_out=16'h0;
17'h86b:	data_out=16'h0;
17'h86c:	data_out=16'h0;
17'h86d:	data_out=16'h0;
17'h86e:	data_out=16'h0;
17'h86f:	data_out=16'h0;
17'h870:	data_out=16'h0;
17'h871:	data_out=16'h0;
17'h872:	data_out=16'h0;
17'h873:	data_out=16'h0;
17'h874:	data_out=16'h0;
17'h875:	data_out=16'h0;
17'h876:	data_out=16'h0;
17'h877:	data_out=16'h0;
17'h878:	data_out=16'h0;
17'h879:	data_out=16'h0;
17'h87a:	data_out=16'h0;
17'h87b:	data_out=16'h0;
17'h87c:	data_out=16'h0;
17'h87d:	data_out=16'haa;
17'h87e:	data_out=16'hff;
17'h87f:	data_out=16'h60;
17'h880:	data_out=16'h0;
17'h881:	data_out=16'h0;
17'h882:	data_out=16'h0;
17'h883:	data_out=16'h0;
17'h884:	data_out=16'h0;
17'h885:	data_out=16'h0;
17'h886:	data_out=16'h0;
17'h887:	data_out=16'h0;
17'h888:	data_out=16'h0;
17'h889:	data_out=16'h0;
17'h88a:	data_out=16'h0;
17'h88b:	data_out=16'h0;
17'h88c:	data_out=16'h0;
17'h88d:	data_out=16'h0;
17'h88e:	data_out=16'h0;
17'h88f:	data_out=16'h0;
17'h890:	data_out=16'h0;
17'h891:	data_out=16'h0;
17'h892:	data_out=16'h0;
17'h893:	data_out=16'h0;
17'h894:	data_out=16'h0;
17'h895:	data_out=16'h0;
17'h896:	data_out=16'h0;
17'h897:	data_out=16'h0;
17'h898:	data_out=16'h0;
17'h899:	data_out=16'haa;
17'h89a:	data_out=16'hff;
17'h89b:	data_out=16'h9a;
17'h89c:	data_out=16'h0;
17'h89d:	data_out=16'h0;
17'h89e:	data_out=16'h0;
17'h89f:	data_out=16'h0;
17'h8a0:	data_out=16'h0;
17'h8a1:	data_out=16'h0;
17'h8a2:	data_out=16'h0;
17'h8a3:	data_out=16'h0;
17'h8a4:	data_out=16'h0;
17'h8a5:	data_out=16'h0;
17'h8a6:	data_out=16'h0;
17'h8a7:	data_out=16'h0;
17'h8a8:	data_out=16'h0;
17'h8a9:	data_out=16'h0;
17'h8aa:	data_out=16'h0;
17'h8ab:	data_out=16'h0;
17'h8ac:	data_out=16'h0;
17'h8ad:	data_out=16'h0;
17'h8ae:	data_out=16'h0;
17'h8af:	data_out=16'h0;
17'h8b0:	data_out=16'h0;
17'h8b1:	data_out=16'h0;
17'h8b2:	data_out=16'h0;
17'h8b3:	data_out=16'h0;
17'h8b4:	data_out=16'h0;
17'h8b5:	data_out=16'haa;
17'h8b6:	data_out=16'h100;
17'h8b7:	data_out=16'h9a;
17'h8b8:	data_out=16'h0;
17'h8b9:	data_out=16'h0;
17'h8ba:	data_out=16'h0;
17'h8bb:	data_out=16'h0;
17'h8bc:	data_out=16'h0;
17'h8bd:	data_out=16'h0;
17'h8be:	data_out=16'h0;
17'h8bf:	data_out=16'h0;
17'h8c0:	data_out=16'h0;
17'h8c1:	data_out=16'h0;
17'h8c2:	data_out=16'h0;
17'h8c3:	data_out=16'h0;
17'h8c4:	data_out=16'h0;
17'h8c5:	data_out=16'h0;
17'h8c6:	data_out=16'h0;
17'h8c7:	data_out=16'h0;
17'h8c8:	data_out=16'h0;
17'h8c9:	data_out=16'h0;
17'h8ca:	data_out=16'h0;
17'h8cb:	data_out=16'h0;
17'h8cc:	data_out=16'h0;
17'h8cd:	data_out=16'h0;
17'h8ce:	data_out=16'h0;
17'h8cf:	data_out=16'h0;
17'h8d0:	data_out=16'h0;
17'h8d1:	data_out=16'h60;
17'h8d2:	data_out=16'hff;
17'h8d3:	data_out=16'h9a;
17'h8d4:	data_out=16'h0;
17'h8d5:	data_out=16'h0;
17'h8d6:	data_out=16'h0;
17'h8d7:	data_out=16'h0;
17'h8d8:	data_out=16'h0;
17'h8d9:	data_out=16'h0;
17'h8da:	data_out=16'h0;
17'h8db:	data_out=16'h0;
17'h8dc:	data_out=16'h0;
17'h8dd:	data_out=16'h0;
17'h8de:	data_out=16'h0;
17'h8df:	data_out=16'h0;
17'h8e0:	data_out=16'h0;
17'h8e1:	data_out=16'h0;
17'h8e2:	data_out=16'h0;
17'h8e3:	data_out=16'h0;
17'h8e4:	data_out=16'h0;
17'h8e5:	data_out=16'h0;
17'h8e6:	data_out=16'h0;
17'h8e7:	data_out=16'h0;
17'h8e8:	data_out=16'h0;
17'h8e9:	data_out=16'h0;
17'h8ea:	data_out=16'h0;
17'h8eb:	data_out=16'h0;
17'h8ec:	data_out=16'h0;
17'h8ed:	data_out=16'h0;
17'h8ee:	data_out=16'h0;
17'h8ef:	data_out=16'h0;
17'h8f0:	data_out=16'h0;
17'h8f1:	data_out=16'h0;
17'h8f2:	data_out=16'h0;
17'h8f3:	data_out=16'h0;
17'h8f4:	data_out=16'h0;
17'h8f5:	data_out=16'h0;
17'h8f6:	data_out=16'h0;
17'h8f7:	data_out=16'h0;
17'h8f8:	data_out=16'h0;
17'h8f9:	data_out=16'h0;
17'h8fa:	data_out=16'h0;
17'h8fb:	data_out=16'h0;
17'h8fc:	data_out=16'h0;
17'h8fd:	data_out=16'h0;
17'h8fe:	data_out=16'h0;
17'h8ff:	data_out=16'h0;
17'h900:	data_out=16'h0;
17'h901:	data_out=16'h0;
17'h902:	data_out=16'h0;
17'h903:	data_out=16'h0;
17'h904:	data_out=16'h0;
17'h905:	data_out=16'h0;
17'h906:	data_out=16'h0;
17'h907:	data_out=16'h0;
17'h908:	data_out=16'h0;
17'h909:	data_out=16'h0;
17'h90a:	data_out=16'h0;
17'h90b:	data_out=16'h0;
17'h90c:	data_out=16'h0;
17'h90d:	data_out=16'h0;
17'h90e:	data_out=16'h0;
17'h90f:	data_out=16'h0;
17'h910:	data_out=16'h0;
17'h911:	data_out=16'h0;
17'h912:	data_out=16'h0;
17'h913:	data_out=16'h0;
17'h914:	data_out=16'h0;
17'h915:	data_out=16'h0;
17'h916:	data_out=16'h0;
17'h917:	data_out=16'h0;
17'h918:	data_out=16'h0;
17'h919:	data_out=16'h0;
17'h91a:	data_out=16'h0;
17'h91b:	data_out=16'h0;
17'h91c:	data_out=16'h0;
17'h91d:	data_out=16'h0;
17'h91e:	data_out=16'h0;
17'h91f:	data_out=16'h0;
17'h920:	data_out=16'h0;
17'h921:	data_out=16'h0;
17'h922:	data_out=16'h0;
17'h923:	data_out=16'h0;
17'h924:	data_out=16'h0;
17'h925:	data_out=16'h0;
17'h926:	data_out=16'h0;
17'h927:	data_out=16'h0;
17'h928:	data_out=16'h0;
17'h929:	data_out=16'h0;
17'h92a:	data_out=16'h0;
17'h92b:	data_out=16'h0;
17'h92c:	data_out=16'h0;
17'h92d:	data_out=16'h0;
17'h92e:	data_out=16'h0;
17'h92f:	data_out=16'h0;
17'h930:	data_out=16'h0;
17'h931:	data_out=16'h0;
17'h932:	data_out=16'h0;
17'h933:	data_out=16'h0;
17'h934:	data_out=16'h0;
17'h935:	data_out=16'h0;
17'h936:	data_out=16'h0;
17'h937:	data_out=16'h0;
17'h938:	data_out=16'h0;
17'h939:	data_out=16'h0;
17'h93a:	data_out=16'h0;
17'h93b:	data_out=16'h0;
17'h93c:	data_out=16'h0;
17'h93d:	data_out=16'h0;
17'h93e:	data_out=16'h0;
17'h93f:	data_out=16'h0;
17'h940:	data_out=16'h0;
17'h941:	data_out=16'h0;
17'h942:	data_out=16'h0;
17'h943:	data_out=16'h0;
17'h944:	data_out=16'h0;
17'h945:	data_out=16'h0;
17'h946:	data_out=16'h0;
17'h947:	data_out=16'h0;
17'h948:	data_out=16'h0;
17'h949:	data_out=16'h0;
17'h94a:	data_out=16'h0;
17'h94b:	data_out=16'h0;
17'h94c:	data_out=16'h0;
17'h94d:	data_out=16'h0;
17'h94e:	data_out=16'h0;
17'h94f:	data_out=16'h0;
17'h950:	data_out=16'h0;
17'h951:	data_out=16'h0;
17'h952:	data_out=16'h0;
17'h953:	data_out=16'h0;
17'h954:	data_out=16'h0;
17'h955:	data_out=16'h0;
17'h956:	data_out=16'h0;
17'h957:	data_out=16'h0;
17'h958:	data_out=16'h0;
17'h959:	data_out=16'h0;
17'h95a:	data_out=16'h0;
17'h95b:	data_out=16'h0;
17'h95c:	data_out=16'h0;
17'h95d:	data_out=16'h0;
17'h95e:	data_out=16'h0;
17'h95f:	data_out=16'h0;
17'h960:	data_out=16'h0;
17'h961:	data_out=16'h0;
17'h962:	data_out=16'h0;
17'h963:	data_out=16'h0;
17'h964:	data_out=16'h0;
17'h965:	data_out=16'h0;
17'h966:	data_out=16'h0;
17'h967:	data_out=16'h0;
17'h968:	data_out=16'h0;
17'h969:	data_out=16'h0;
17'h96a:	data_out=16'h0;
17'h96b:	data_out=16'h0;
17'h96c:	data_out=16'h0;
17'h96d:	data_out=16'h0;
17'h96e:	data_out=16'h0;
17'h96f:	data_out=16'h0;
17'h970:	data_out=16'h0;
17'h971:	data_out=16'h0;
17'h972:	data_out=16'h0;
17'h973:	data_out=16'h0;
17'h974:	data_out=16'h0;
17'h975:	data_out=16'h0;
17'h976:	data_out=16'h0;
17'h977:	data_out=16'h0;
17'h978:	data_out=16'h0;
17'h979:	data_out=16'h0;
17'h97a:	data_out=16'h0;
17'h97b:	data_out=16'h0;
17'h97c:	data_out=16'h0;
17'h97d:	data_out=16'h0;
17'h97e:	data_out=16'h0;
17'h97f:	data_out=16'h0;
17'h980:	data_out=16'h0;
17'h981:	data_out=16'h0;
17'h982:	data_out=16'h0;
17'h983:	data_out=16'h0;
17'h984:	data_out=16'h0;
17'h985:	data_out=16'h0;
17'h986:	data_out=16'h0;
17'h987:	data_out=16'h0;
17'h988:	data_out=16'h0;
17'h989:	data_out=16'h0;
17'h98a:	data_out=16'h0;
17'h98b:	data_out=16'h0;
17'h98c:	data_out=16'h0;
17'h98d:	data_out=16'h0;
17'h98e:	data_out=16'h0;
17'h98f:	data_out=16'h0;
17'h990:	data_out=16'h0;
17'h991:	data_out=16'h0;
17'h992:	data_out=16'h0;
17'h993:	data_out=16'h0;
17'h994:	data_out=16'h0;
17'h995:	data_out=16'h0;
17'h996:	data_out=16'h0;
17'h997:	data_out=16'h0;
17'h998:	data_out=16'h0;
17'h999:	data_out=16'h0;
17'h99a:	data_out=16'h0;
17'h99b:	data_out=16'h0;
17'h99c:	data_out=16'h0;
17'h99d:	data_out=16'h0;
17'h99e:	data_out=16'h0;
17'h99f:	data_out=16'h0;
17'h9a0:	data_out=16'h0;
17'h9a1:	data_out=16'h0;
17'h9a2:	data_out=16'h0;
17'h9a3:	data_out=16'h0;
17'h9a4:	data_out=16'h0;
17'h9a5:	data_out=16'h0;
17'h9a6:	data_out=16'h0;
17'h9a7:	data_out=16'h0;
17'h9a8:	data_out=16'h0;
17'h9a9:	data_out=16'h0;
17'h9aa:	data_out=16'h0;
17'h9ab:	data_out=16'h0;
17'h9ac:	data_out=16'h0;
17'h9ad:	data_out=16'h0;
17'h9ae:	data_out=16'h0;
17'h9af:	data_out=16'h0;
17'h9b0:	data_out=16'h0;
17'h9b1:	data_out=16'h0;
17'h9b2:	data_out=16'h0;
17'h9b3:	data_out=16'h0;
17'h9b4:	data_out=16'h0;
17'h9b5:	data_out=16'h0;
17'h9b6:	data_out=16'h0;
17'h9b7:	data_out=16'h0;
17'h9b8:	data_out=16'h0;
17'h9b9:	data_out=16'h0;
17'h9ba:	data_out=16'h0;
17'h9bb:	data_out=16'h0;
17'h9bc:	data_out=16'h0;
17'h9bd:	data_out=16'h0;
17'h9be:	data_out=16'h0;
17'h9bf:	data_out=16'h0;
17'h9c0:	data_out=16'h0;
17'h9c1:	data_out=16'h0;
17'h9c2:	data_out=16'h0;
17'h9c3:	data_out=16'h0;
17'h9c4:	data_out=16'h0;
17'h9c5:	data_out=16'h0;
17'h9c6:	data_out=16'h0;
17'h9c7:	data_out=16'h0;
17'h9c8:	data_out=16'h0;
17'h9c9:	data_out=16'h0;
17'h9ca:	data_out=16'h0;
17'h9cb:	data_out=16'h0;
17'h9cc:	data_out=16'h0;
17'h9cd:	data_out=16'h0;
17'h9ce:	data_out=16'h7c;
17'h9cf:	data_out=16'hfe;
17'h9d0:	data_out=16'h100;
17'h9d1:	data_out=16'h3f;
17'h9d2:	data_out=16'h0;
17'h9d3:	data_out=16'h0;
17'h9d4:	data_out=16'h0;
17'h9d5:	data_out=16'h0;
17'h9d6:	data_out=16'h0;
17'h9d7:	data_out=16'h0;
17'h9d8:	data_out=16'h0;
17'h9d9:	data_out=16'h0;
17'h9da:	data_out=16'h0;
17'h9db:	data_out=16'h0;
17'h9dc:	data_out=16'h0;
17'h9dd:	data_out=16'h0;
17'h9de:	data_out=16'h0;
17'h9df:	data_out=16'h0;
17'h9e0:	data_out=16'h0;
17'h9e1:	data_out=16'h0;
17'h9e2:	data_out=16'h0;
17'h9e3:	data_out=16'h0;
17'h9e4:	data_out=16'h0;
17'h9e5:	data_out=16'h0;
17'h9e6:	data_out=16'h0;
17'h9e7:	data_out=16'h0;
17'h9e8:	data_out=16'h0;
17'h9e9:	data_out=16'h60;
17'h9ea:	data_out=16'hf5;
17'h9eb:	data_out=16'hfc;
17'h9ec:	data_out=16'hfe;
17'h9ed:	data_out=16'h3e;
17'h9ee:	data_out=16'h0;
17'h9ef:	data_out=16'h0;
17'h9f0:	data_out=16'h0;
17'h9f1:	data_out=16'h0;
17'h9f2:	data_out=16'h0;
17'h9f3:	data_out=16'h0;
17'h9f4:	data_out=16'h0;
17'h9f5:	data_out=16'h0;
17'h9f6:	data_out=16'h0;
17'h9f7:	data_out=16'h0;
17'h9f8:	data_out=16'h0;
17'h9f9:	data_out=16'h0;
17'h9fa:	data_out=16'h0;
17'h9fb:	data_out=16'h0;
17'h9fc:	data_out=16'h0;
17'h9fd:	data_out=16'h0;
17'h9fe:	data_out=16'h0;
17'h9ff:	data_out=16'h0;
17'ha00:	data_out=16'h0;
17'ha01:	data_out=16'h0;
17'ha02:	data_out=16'h0;
17'ha03:	data_out=16'h0;
17'ha04:	data_out=16'h0;
17'ha05:	data_out=16'h7f;
17'ha06:	data_out=16'hfc;
17'ha07:	data_out=16'hfc;
17'ha08:	data_out=16'hfe;
17'ha09:	data_out=16'h3e;
17'ha0a:	data_out=16'h0;
17'ha0b:	data_out=16'h0;
17'ha0c:	data_out=16'h0;
17'ha0d:	data_out=16'h0;
17'ha0e:	data_out=16'h0;
17'ha0f:	data_out=16'h0;
17'ha10:	data_out=16'h0;
17'ha11:	data_out=16'h0;
17'ha12:	data_out=16'h0;
17'ha13:	data_out=16'h0;
17'ha14:	data_out=16'h0;
17'ha15:	data_out=16'h0;
17'ha16:	data_out=16'h0;
17'ha17:	data_out=16'h0;
17'ha18:	data_out=16'h0;
17'ha19:	data_out=16'h0;
17'ha1a:	data_out=16'h0;
17'ha1b:	data_out=16'h0;
17'ha1c:	data_out=16'h0;
17'ha1d:	data_out=16'h0;
17'ha1e:	data_out=16'h0;
17'ha1f:	data_out=16'h0;
17'ha20:	data_out=16'h44;
17'ha21:	data_out=16'hed;
17'ha22:	data_out=16'hfc;
17'ha23:	data_out=16'hd4;
17'ha24:	data_out=16'h1f;
17'ha25:	data_out=16'h8;
17'ha26:	data_out=16'h0;
17'ha27:	data_out=16'h0;
17'ha28:	data_out=16'h0;
17'ha29:	data_out=16'h0;
17'ha2a:	data_out=16'h0;
17'ha2b:	data_out=16'h0;
17'ha2c:	data_out=16'h0;
17'ha2d:	data_out=16'h0;
17'ha2e:	data_out=16'h0;
17'ha2f:	data_out=16'h0;
17'ha30:	data_out=16'h0;
17'ha31:	data_out=16'h0;
17'ha32:	data_out=16'h0;
17'ha33:	data_out=16'h0;
17'ha34:	data_out=16'h0;
17'ha35:	data_out=16'h0;
17'ha36:	data_out=16'h0;
17'ha37:	data_out=16'h0;
17'ha38:	data_out=16'h0;
17'ha39:	data_out=16'h0;
17'ha3a:	data_out=16'h0;
17'ha3b:	data_out=16'h3c;
17'ha3c:	data_out=16'he5;
17'ha3d:	data_out=16'hfc;
17'ha3e:	data_out=16'hfc;
17'ha3f:	data_out=16'h5e;
17'ha40:	data_out=16'h0;
17'ha41:	data_out=16'h0;
17'ha42:	data_out=16'h0;
17'ha43:	data_out=16'h0;
17'ha44:	data_out=16'h0;
17'ha45:	data_out=16'h0;
17'ha46:	data_out=16'h0;
17'ha47:	data_out=16'h0;
17'ha48:	data_out=16'h0;
17'ha49:	data_out=16'h0;
17'ha4a:	data_out=16'h0;
17'ha4b:	data_out=16'h0;
17'ha4c:	data_out=16'h0;
17'ha4d:	data_out=16'h0;
17'ha4e:	data_out=16'h0;
17'ha4f:	data_out=16'h0;
17'ha50:	data_out=16'h0;
17'ha51:	data_out=16'h0;
17'ha52:	data_out=16'h0;
17'ha53:	data_out=16'h0;
17'ha54:	data_out=16'h0;
17'ha55:	data_out=16'h0;
17'ha56:	data_out=16'h0;
17'ha57:	data_out=16'h9c;
17'ha58:	data_out=16'hfe;
17'ha59:	data_out=16'hfe;
17'ha5a:	data_out=16'hbe;
17'ha5b:	data_out=16'h0;
17'ha5c:	data_out=16'h0;
17'ha5d:	data_out=16'h0;
17'ha5e:	data_out=16'h0;
17'ha5f:	data_out=16'h0;
17'ha60:	data_out=16'h0;
17'ha61:	data_out=16'h0;
17'ha62:	data_out=16'h0;
17'ha63:	data_out=16'h0;
17'ha64:	data_out=16'h0;
17'ha65:	data_out=16'h0;
17'ha66:	data_out=16'h0;
17'ha67:	data_out=16'h0;
17'ha68:	data_out=16'h0;
17'ha69:	data_out=16'h0;
17'ha6a:	data_out=16'h0;
17'ha6b:	data_out=16'h0;
17'ha6c:	data_out=16'h0;
17'ha6d:	data_out=16'h0;
17'ha6e:	data_out=16'h0;
17'ha6f:	data_out=16'h0;
17'ha70:	data_out=16'h0;
17'ha71:	data_out=16'h0;
17'ha72:	data_out=16'h14;
17'ha73:	data_out=16'hfe;
17'ha74:	data_out=16'hfc;
17'ha75:	data_out=16'hec;
17'ha76:	data_out=16'h42;
17'ha77:	data_out=16'h0;
17'ha78:	data_out=16'h0;
17'ha79:	data_out=16'h0;
17'ha7a:	data_out=16'h0;
17'ha7b:	data_out=16'h0;
17'ha7c:	data_out=16'h0;
17'ha7d:	data_out=16'h0;
17'ha7e:	data_out=16'h0;
17'ha7f:	data_out=16'h0;
17'ha80:	data_out=16'h0;
17'ha81:	data_out=16'h0;
17'ha82:	data_out=16'h0;
17'ha83:	data_out=16'h0;
17'ha84:	data_out=16'h0;
17'ha85:	data_out=16'h0;
17'ha86:	data_out=16'h0;
17'ha87:	data_out=16'h0;
17'ha88:	data_out=16'h0;
17'ha89:	data_out=16'h0;
17'ha8a:	data_out=16'h0;
17'ha8b:	data_out=16'h0;
17'ha8c:	data_out=16'h0;
17'ha8d:	data_out=16'h20;
17'ha8e:	data_out=16'hce;
17'ha8f:	data_out=16'hfe;
17'ha90:	data_out=16'hfc;
17'ha91:	data_out=16'h7e;
17'ha92:	data_out=16'h0;
17'ha93:	data_out=16'h0;
17'ha94:	data_out=16'h0;
17'ha95:	data_out=16'h0;
17'ha96:	data_out=16'h0;
17'ha97:	data_out=16'h0;
17'ha98:	data_out=16'h0;
17'ha99:	data_out=16'h0;
17'ha9a:	data_out=16'h0;
17'ha9b:	data_out=16'h0;
17'ha9c:	data_out=16'h0;
17'ha9d:	data_out=16'h0;
17'ha9e:	data_out=16'h0;
17'ha9f:	data_out=16'h0;
17'haa0:	data_out=16'h0;
17'haa1:	data_out=16'h0;
17'haa2:	data_out=16'h0;
17'haa3:	data_out=16'h0;
17'haa4:	data_out=16'h0;
17'haa5:	data_out=16'h0;
17'haa6:	data_out=16'h0;
17'haa7:	data_out=16'h0;
17'haa8:	data_out=16'h0;
17'haa9:	data_out=16'h68;
17'haaa:	data_out=16'hfc;
17'haab:	data_out=16'hfe;
17'haac:	data_out=16'hb9;
17'haad:	data_out=16'hf;
17'haae:	data_out=16'h0;
17'haaf:	data_out=16'h0;
17'hab0:	data_out=16'h0;
17'hab1:	data_out=16'h0;
17'hab2:	data_out=16'h0;
17'hab3:	data_out=16'h0;
17'hab4:	data_out=16'h0;
17'hab5:	data_out=16'h0;
17'hab6:	data_out=16'h0;
17'hab7:	data_out=16'h0;
17'hab8:	data_out=16'h0;
17'hab9:	data_out=16'h0;
17'haba:	data_out=16'h0;
17'habb:	data_out=16'h0;
17'habc:	data_out=16'h0;
17'habd:	data_out=16'h0;
17'habe:	data_out=16'h0;
17'habf:	data_out=16'h0;
17'hac0:	data_out=16'h0;
17'hac1:	data_out=16'h0;
17'hac2:	data_out=16'h0;
17'hac3:	data_out=16'h0;
17'hac4:	data_out=16'h50;
17'hac5:	data_out=16'hf1;
17'hac6:	data_out=16'hfc;
17'hac7:	data_out=16'hc2;
17'hac8:	data_out=16'h17;
17'hac9:	data_out=16'h0;
17'haca:	data_out=16'h0;
17'hacb:	data_out=16'h0;
17'hacc:	data_out=16'h0;
17'hacd:	data_out=16'h0;
17'hace:	data_out=16'h0;
17'hacf:	data_out=16'h0;
17'had0:	data_out=16'h0;
17'had1:	data_out=16'h0;
17'had2:	data_out=16'h0;
17'had3:	data_out=16'h0;
17'had4:	data_out=16'h0;
17'had5:	data_out=16'h0;
17'had6:	data_out=16'h0;
17'had7:	data_out=16'h0;
17'had8:	data_out=16'h0;
17'had9:	data_out=16'h0;
17'hada:	data_out=16'h0;
17'hadb:	data_out=16'h0;
17'hadc:	data_out=16'h0;
17'hadd:	data_out=16'h0;
17'hade:	data_out=16'h0;
17'hadf:	data_out=16'h20;
17'hae0:	data_out=16'hfe;
17'hae1:	data_out=16'hfe;
17'hae2:	data_out=16'hfe;
17'hae3:	data_out=16'ha0;
17'hae4:	data_out=16'h0;
17'hae5:	data_out=16'h0;
17'hae6:	data_out=16'h0;
17'hae7:	data_out=16'h0;
17'hae8:	data_out=16'h0;
17'hae9:	data_out=16'h0;
17'haea:	data_out=16'h0;
17'haeb:	data_out=16'h0;
17'haec:	data_out=16'h0;
17'haed:	data_out=16'h0;
17'haee:	data_out=16'h0;
17'haef:	data_out=16'h0;
17'haf0:	data_out=16'h0;
17'haf1:	data_out=16'h0;
17'haf2:	data_out=16'h0;
17'haf3:	data_out=16'h0;
17'haf4:	data_out=16'h0;
17'haf5:	data_out=16'h0;
17'haf6:	data_out=16'h0;
17'haf7:	data_out=16'h0;
17'haf8:	data_out=16'h0;
17'haf9:	data_out=16'h0;
17'hafa:	data_out=16'h0;
17'hafb:	data_out=16'h98;
17'hafc:	data_out=16'hfc;
17'hafd:	data_out=16'hfc;
17'hafe:	data_out=16'hfc;
17'haff:	data_out=16'h27;
17'hb00:	data_out=16'h0;
17'hb01:	data_out=16'h0;
17'hb02:	data_out=16'h0;
17'hb03:	data_out=16'h0;
17'hb04:	data_out=16'h0;
17'hb05:	data_out=16'h0;
17'hb06:	data_out=16'h0;
17'hb07:	data_out=16'h0;
17'hb08:	data_out=16'h0;
17'hb09:	data_out=16'h0;
17'hb0a:	data_out=16'h0;
17'hb0b:	data_out=16'h0;
17'hb0c:	data_out=16'h0;
17'hb0d:	data_out=16'h0;
17'hb0e:	data_out=16'h0;
17'hb0f:	data_out=16'h0;
17'hb10:	data_out=16'h0;
17'hb11:	data_out=16'h0;
17'hb12:	data_out=16'h0;
17'hb13:	data_out=16'h0;
17'hb14:	data_out=16'h0;
17'hb15:	data_out=16'h0;
17'hb16:	data_out=16'h30;
17'hb17:	data_out=16'hde;
17'hb18:	data_out=16'hfc;
17'hb19:	data_out=16'hfc;
17'hb1a:	data_out=16'had;
17'hb1b:	data_out=16'h0;
17'hb1c:	data_out=16'h0;
17'hb1d:	data_out=16'h0;
17'hb1e:	data_out=16'h0;
17'hb1f:	data_out=16'h0;
17'hb20:	data_out=16'h0;
17'hb21:	data_out=16'h0;
17'hb22:	data_out=16'h0;
17'hb23:	data_out=16'h0;
17'hb24:	data_out=16'h0;
17'hb25:	data_out=16'h0;
17'hb26:	data_out=16'h0;
17'hb27:	data_out=16'h0;
17'hb28:	data_out=16'h0;
17'hb29:	data_out=16'h0;
17'hb2a:	data_out=16'h0;
17'hb2b:	data_out=16'h0;
17'hb2c:	data_out=16'h0;
17'hb2d:	data_out=16'h0;
17'hb2e:	data_out=16'h0;
17'hb2f:	data_out=16'h0;
17'hb30:	data_out=16'h0;
17'hb31:	data_out=16'h0;
17'hb32:	data_out=16'heb;
17'hb33:	data_out=16'hfc;
17'hb34:	data_out=16'hfc;
17'hb35:	data_out=16'hc5;
17'hb36:	data_out=16'hc;
17'hb37:	data_out=16'h0;
17'hb38:	data_out=16'h0;
17'hb39:	data_out=16'h0;
17'hb3a:	data_out=16'h0;
17'hb3b:	data_out=16'h0;
17'hb3c:	data_out=16'h0;
17'hb3d:	data_out=16'h0;
17'hb3e:	data_out=16'h0;
17'hb3f:	data_out=16'h0;
17'hb40:	data_out=16'h0;
17'hb41:	data_out=16'h0;
17'hb42:	data_out=16'h0;
17'hb43:	data_out=16'h0;
17'hb44:	data_out=16'h0;
17'hb45:	data_out=16'h0;
17'hb46:	data_out=16'h0;
17'hb47:	data_out=16'h0;
17'hb48:	data_out=16'h0;
17'hb49:	data_out=16'h0;
17'hb4a:	data_out=16'h0;
17'hb4b:	data_out=16'h0;
17'hb4c:	data_out=16'h0;
17'hb4d:	data_out=16'h0;
17'hb4e:	data_out=16'hfe;
17'hb4f:	data_out=16'hfc;
17'hb50:	data_out=16'hfc;
17'hb51:	data_out=16'h59;
17'hb52:	data_out=16'h0;
17'hb53:	data_out=16'h0;
17'hb54:	data_out=16'h0;
17'hb55:	data_out=16'h0;
17'hb56:	data_out=16'h0;
17'hb57:	data_out=16'h0;
17'hb58:	data_out=16'h0;
17'hb59:	data_out=16'h0;
17'hb5a:	data_out=16'h0;
17'hb5b:	data_out=16'h0;
17'hb5c:	data_out=16'h0;
17'hb5d:	data_out=16'h0;
17'hb5e:	data_out=16'h0;
17'hb5f:	data_out=16'h0;
17'hb60:	data_out=16'h0;
17'hb61:	data_out=16'h0;
17'hb62:	data_out=16'h0;
17'hb63:	data_out=16'h0;
17'hb64:	data_out=16'h0;
17'hb65:	data_out=16'h0;
17'hb66:	data_out=16'h0;
17'hb67:	data_out=16'h0;
17'hb68:	data_out=16'h0;
17'hb69:	data_out=16'ha0;
17'hb6a:	data_out=16'h100;
17'hb6b:	data_out=16'hfe;
17'hb6c:	data_out=16'hfe;
17'hb6d:	data_out=16'h1f;
17'hb6e:	data_out=16'h0;
17'hb6f:	data_out=16'h0;
17'hb70:	data_out=16'h0;
17'hb71:	data_out=16'h0;
17'hb72:	data_out=16'h0;
17'hb73:	data_out=16'h0;
17'hb74:	data_out=16'h0;
17'hb75:	data_out=16'h0;
17'hb76:	data_out=16'h0;
17'hb77:	data_out=16'h0;
17'hb78:	data_out=16'h0;
17'hb79:	data_out=16'h0;
17'hb7a:	data_out=16'h0;
17'hb7b:	data_out=16'h0;
17'hb7c:	data_out=16'h0;
17'hb7d:	data_out=16'h0;
17'hb7e:	data_out=16'h0;
17'hb7f:	data_out=16'h0;
17'hb80:	data_out=16'h0;
17'hb81:	data_out=16'h0;
17'hb82:	data_out=16'h0;
17'hb83:	data_out=16'h0;
17'hb84:	data_out=16'h30;
17'hb85:	data_out=16'he5;
17'hb86:	data_out=16'hfe;
17'hb87:	data_out=16'hf8;
17'hb88:	data_out=16'h8d;
17'hb89:	data_out=16'h8;
17'hb8a:	data_out=16'h0;
17'hb8b:	data_out=16'h0;
17'hb8c:	data_out=16'h0;
17'hb8d:	data_out=16'h0;
17'hb8e:	data_out=16'h0;
17'hb8f:	data_out=16'h0;
17'hb90:	data_out=16'h0;
17'hb91:	data_out=16'h0;
17'hb92:	data_out=16'h0;
17'hb93:	data_out=16'h0;
17'hb94:	data_out=16'h0;
17'hb95:	data_out=16'h0;
17'hb96:	data_out=16'h0;
17'hb97:	data_out=16'h0;
17'hb98:	data_out=16'h0;
17'hb99:	data_out=16'h0;
17'hb9a:	data_out=16'h0;
17'hb9b:	data_out=16'h0;
17'hb9c:	data_out=16'h0;
17'hb9d:	data_out=16'h0;
17'hb9e:	data_out=16'h0;
17'hb9f:	data_out=16'h0;
17'hba0:	data_out=16'h40;
17'hba1:	data_out=16'hfc;
17'hba2:	data_out=16'hfe;
17'hba3:	data_out=16'hdd;
17'hba4:	data_out=16'h0;
17'hba5:	data_out=16'h0;
17'hba6:	data_out=16'h0;
17'hba7:	data_out=16'h0;
17'hba8:	data_out=16'h0;
17'hba9:	data_out=16'h0;
17'hbaa:	data_out=16'h0;
17'hbab:	data_out=16'h0;
17'hbac:	data_out=16'h0;
17'hbad:	data_out=16'h0;
17'hbae:	data_out=16'h0;
17'hbaf:	data_out=16'h0;
17'hbb0:	data_out=16'h0;
17'hbb1:	data_out=16'h0;
17'hbb2:	data_out=16'h0;
17'hbb3:	data_out=16'h0;
17'hbb4:	data_out=16'h0;
17'hbb5:	data_out=16'h0;
17'hbb6:	data_out=16'h0;
17'hbb7:	data_out=16'h0;
17'hbb8:	data_out=16'h0;
17'hbb9:	data_out=16'h0;
17'hbba:	data_out=16'h0;
17'hbbb:	data_out=16'h0;
17'hbbc:	data_out=16'h40;
17'hbbd:	data_out=16'hfc;
17'hbbe:	data_out=16'hfe;
17'hbbf:	data_out=16'hdd;
17'hbc0:	data_out=16'h0;
17'hbc1:	data_out=16'h0;
17'hbc2:	data_out=16'h0;
17'hbc3:	data_out=16'h0;
17'hbc4:	data_out=16'h0;
17'hbc5:	data_out=16'h0;
17'hbc6:	data_out=16'h0;
17'hbc7:	data_out=16'h0;
17'hbc8:	data_out=16'h0;
17'hbc9:	data_out=16'h0;
17'hbca:	data_out=16'h0;
17'hbcb:	data_out=16'h0;
17'hbcc:	data_out=16'h0;
17'hbcd:	data_out=16'h0;
17'hbce:	data_out=16'h0;
17'hbcf:	data_out=16'h0;
17'hbd0:	data_out=16'h0;
17'hbd1:	data_out=16'h0;
17'hbd2:	data_out=16'h0;
17'hbd3:	data_out=16'h0;
17'hbd4:	data_out=16'h0;
17'hbd5:	data_out=16'h0;
17'hbd6:	data_out=16'h0;
17'hbd7:	data_out=16'h0;
17'hbd8:	data_out=16'h18;
17'hbd9:	data_out=16'hc2;
17'hbda:	data_out=16'hfe;
17'hbdb:	data_out=16'hdd;
17'hbdc:	data_out=16'h0;
17'hbdd:	data_out=16'h0;
17'hbde:	data_out=16'h0;
17'hbdf:	data_out=16'h0;
17'hbe0:	data_out=16'h0;
17'hbe1:	data_out=16'h0;
17'hbe2:	data_out=16'h0;
17'hbe3:	data_out=16'h0;
17'hbe4:	data_out=16'h0;
17'hbe5:	data_out=16'h0;
17'hbe6:	data_out=16'h0;
17'hbe7:	data_out=16'h0;
17'hbe8:	data_out=16'h0;
17'hbe9:	data_out=16'h0;
17'hbea:	data_out=16'h0;
17'hbeb:	data_out=16'h0;
17'hbec:	data_out=16'h0;
17'hbed:	data_out=16'h0;
17'hbee:	data_out=16'h0;
17'hbef:	data_out=16'h0;
17'hbf0:	data_out=16'h0;
17'hbf1:	data_out=16'h0;
17'hbf2:	data_out=16'h0;
17'hbf3:	data_out=16'h0;
17'hbf4:	data_out=16'h0;
17'hbf5:	data_out=16'h0;
17'hbf6:	data_out=16'h0;
17'hbf7:	data_out=16'h0;
17'hbf8:	data_out=16'h0;
17'hbf9:	data_out=16'h0;
17'hbfa:	data_out=16'h0;
17'hbfb:	data_out=16'h0;
17'hbfc:	data_out=16'h0;
17'hbfd:	data_out=16'h0;
17'hbfe:	data_out=16'h0;
17'hbff:	data_out=16'h0;
17'hc00:	data_out=16'h0;
17'hc01:	data_out=16'h0;
17'hc02:	data_out=16'h0;
17'hc03:	data_out=16'h0;
17'hc04:	data_out=16'h0;
17'hc05:	data_out=16'h0;
17'hc06:	data_out=16'h0;
17'hc07:	data_out=16'h0;
17'hc08:	data_out=16'h0;
17'hc09:	data_out=16'h0;
17'hc0a:	data_out=16'h0;
17'hc0b:	data_out=16'h0;
17'hc0c:	data_out=16'h0;
17'hc0d:	data_out=16'h0;
17'hc0e:	data_out=16'h0;
17'hc0f:	data_out=16'h0;
17'hc10:	data_out=16'h0;
17'hc11:	data_out=16'h0;
17'hc12:	data_out=16'h0;
17'hc13:	data_out=16'h0;
17'hc14:	data_out=16'h0;
17'hc15:	data_out=16'h0;
17'hc16:	data_out=16'h0;
17'hc17:	data_out=16'h0;
17'hc18:	data_out=16'h0;
17'hc19:	data_out=16'h0;
17'hc1a:	data_out=16'h0;
17'hc1b:	data_out=16'h0;
17'hc1c:	data_out=16'h0;
17'hc1d:	data_out=16'h0;
17'hc1e:	data_out=16'h0;
17'hc1f:	data_out=16'h0;
17'hc20:	data_out=16'h0;
17'hc21:	data_out=16'h0;
17'hc22:	data_out=16'h0;
17'hc23:	data_out=16'h0;
17'hc24:	data_out=16'h0;
17'hc25:	data_out=16'h0;
17'hc26:	data_out=16'h0;
17'hc27:	data_out=16'h0;
17'hc28:	data_out=16'h0;
17'hc29:	data_out=16'h0;
17'hc2a:	data_out=16'h0;
17'hc2b:	data_out=16'h0;
17'hc2c:	data_out=16'h0;
17'hc2d:	data_out=16'h0;
17'hc2e:	data_out=16'h0;
17'hc2f:	data_out=16'h0;
17'hc30:	data_out=16'h0;
17'hc31:	data_out=16'h0;
17'hc32:	data_out=16'h0;
17'hc33:	data_out=16'h0;
17'hc34:	data_out=16'h0;
17'hc35:	data_out=16'h0;
17'hc36:	data_out=16'h0;
17'hc37:	data_out=16'h0;
17'hc38:	data_out=16'h0;
17'hc39:	data_out=16'h0;
17'hc3a:	data_out=16'h0;
17'hc3b:	data_out=16'h0;
17'hc3c:	data_out=16'h0;
17'hc3d:	data_out=16'h0;
17'hc3e:	data_out=16'h0;
17'hc3f:	data_out=16'h0;
17'hc40:	data_out=16'h0;
17'hc41:	data_out=16'h0;
17'hc42:	data_out=16'h0;
17'hc43:	data_out=16'h0;
17'hc44:	data_out=16'h0;
17'hc45:	data_out=16'h0;
17'hc46:	data_out=16'h0;
17'hc47:	data_out=16'h0;
17'hc48:	data_out=16'h0;
17'hc49:	data_out=16'h0;
17'hc4a:	data_out=16'h0;
17'hc4b:	data_out=16'h0;
17'hc4c:	data_out=16'h0;
17'hc4d:	data_out=16'h0;
17'hc4e:	data_out=16'h0;
17'hc4f:	data_out=16'h0;
17'hc50:	data_out=16'h0;
17'hc51:	data_out=16'h0;
17'hc52:	data_out=16'h0;
17'hc53:	data_out=16'h0;
17'hc54:	data_out=16'h0;
17'hc55:	data_out=16'h0;
17'hc56:	data_out=16'h0;
17'hc57:	data_out=16'h0;
17'hc58:	data_out=16'h0;
17'hc59:	data_out=16'h0;
17'hc5a:	data_out=16'h0;
17'hc5b:	data_out=16'h0;
17'hc5c:	data_out=16'h0;
17'hc5d:	data_out=16'h0;
17'hc5e:	data_out=16'h0;
17'hc5f:	data_out=16'h0;
17'hc60:	data_out=16'h0;
17'hc61:	data_out=16'h0;
17'hc62:	data_out=16'h0;
17'hc63:	data_out=16'h0;
17'hc64:	data_out=16'h0;
17'hc65:	data_out=16'h0;
17'hc66:	data_out=16'h0;
17'hc67:	data_out=16'h0;
17'hc68:	data_out=16'h0;
17'hc69:	data_out=16'h0;
17'hc6a:	data_out=16'h0;
17'hc6b:	data_out=16'h0;
17'hc6c:	data_out=16'h0;
17'hc6d:	data_out=16'h0;
17'hc6e:	data_out=16'h0;
17'hc6f:	data_out=16'h0;
17'hc70:	data_out=16'h0;
17'hc71:	data_out=16'h0;
17'hc72:	data_out=16'h0;
17'hc73:	data_out=16'h0;
17'hc74:	data_out=16'h0;
17'hc75:	data_out=16'h0;
17'hc76:	data_out=16'h0;
17'hc77:	data_out=16'h0;
17'hc78:	data_out=16'h0;
17'hc79:	data_out=16'h0;
17'hc7a:	data_out=16'h0;
17'hc7b:	data_out=16'h0;
17'hc7c:	data_out=16'h0;
17'hc7d:	data_out=16'h0;
17'hc7e:	data_out=16'h0;
17'hc7f:	data_out=16'h0;
17'hc80:	data_out=16'h0;
17'hc81:	data_out=16'h0;
17'hc82:	data_out=16'h0;
17'hc83:	data_out=16'h0;
17'hc84:	data_out=16'h0;
17'hc85:	data_out=16'h0;
17'hc86:	data_out=16'h0;
17'hc87:	data_out=16'h0;
17'hc88:	data_out=16'h0;
17'hc89:	data_out=16'h0;
17'hc8a:	data_out=16'h0;
17'hc8b:	data_out=16'h0;
17'hc8c:	data_out=16'h0;
17'hc8d:	data_out=16'h0;
17'hc8e:	data_out=16'h0;
17'hc8f:	data_out=16'h0;
17'hc90:	data_out=16'h0;
17'hc91:	data_out=16'h0;
17'hc92:	data_out=16'h0;
17'hc93:	data_out=16'h0;
17'hc94:	data_out=16'h0;
17'hc95:	data_out=16'h0;
17'hc96:	data_out=16'h0;
17'hc97:	data_out=16'h0;
17'hc98:	data_out=16'h0;
17'hc99:	data_out=16'h0;
17'hc9a:	data_out=16'h0;
17'hc9b:	data_out=16'h0;
17'hc9c:	data_out=16'h0;
17'hc9d:	data_out=16'h0;
17'hc9e:	data_out=16'h0;
17'hc9f:	data_out=16'h0;
17'hca0:	data_out=16'h0;
17'hca1:	data_out=16'h0;
17'hca2:	data_out=16'h0;
17'hca3:	data_out=16'h0;
17'hca4:	data_out=16'h0;
17'hca5:	data_out=16'h0;
17'hca6:	data_out=16'h0;
17'hca7:	data_out=16'h0;
17'hca8:	data_out=16'h0;
17'hca9:	data_out=16'h0;
17'hcaa:	data_out=16'h0;
17'hcab:	data_out=16'h0;
17'hcac:	data_out=16'h0;
17'hcad:	data_out=16'h0;
17'hcae:	data_out=16'h0;
17'hcaf:	data_out=16'h0;
17'hcb0:	data_out=16'h0;
17'hcb1:	data_out=16'h0;
17'hcb2:	data_out=16'h0;
17'hcb3:	data_out=16'h0;
17'hcb4:	data_out=16'h0;
17'hcb5:	data_out=16'h0;
17'hcb6:	data_out=16'h0;
17'hcb7:	data_out=16'h0;
17'hcb8:	data_out=16'h0;
17'hcb9:	data_out=16'h0;
17'hcba:	data_out=16'h0;
17'hcbb:	data_out=16'h0;
17'hcbc:	data_out=16'h0;
17'hcbd:	data_out=16'h0;
17'hcbe:	data_out=16'h0;
17'hcbf:	data_out=16'h0;
17'hcc0:	data_out=16'h0;
17'hcc1:	data_out=16'h0;
17'hcc2:	data_out=16'h0;
17'hcc3:	data_out=16'h0;
17'hcc4:	data_out=16'h0;
17'hcc5:	data_out=16'h0;
17'hcc6:	data_out=16'h0;
17'hcc7:	data_out=16'h0;
17'hcc8:	data_out=16'h0;
17'hcc9:	data_out=16'h0;
17'hcca:	data_out=16'h0;
17'hccb:	data_out=16'h0;
17'hccc:	data_out=16'h0;
17'hccd:	data_out=16'h0;
17'hcce:	data_out=16'h0;
17'hccf:	data_out=16'h0;
17'hcd0:	data_out=16'h0;
17'hcd1:	data_out=16'h0;
17'hcd2:	data_out=16'h0;
17'hcd3:	data_out=16'h0;
17'hcd4:	data_out=16'h0;
17'hcd5:	data_out=16'h0;
17'hcd6:	data_out=16'h0;
17'hcd7:	data_out=16'h0;
17'hcd8:	data_out=16'h0;
17'hcd9:	data_out=16'h0;
17'hcda:	data_out=16'h0;
17'hcdb:	data_out=16'h0;
17'hcdc:	data_out=16'h0;
17'hcdd:	data_out=16'h0;
17'hcde:	data_out=16'h0;
17'hcdf:	data_out=16'h0;
17'hce0:	data_out=16'h0;
17'hce1:	data_out=16'h0;
17'hce2:	data_out=16'h0;
17'hce3:	data_out=16'h0;
17'hce4:	data_out=16'h0;
17'hce5:	data_out=16'h0;
17'hce6:	data_out=16'h0;
17'hce7:	data_out=16'h0;
17'hce8:	data_out=16'h0;
17'hce9:	data_out=16'h0;
17'hcea:	data_out=16'h0;
17'hceb:	data_out=16'h0;
17'hcec:	data_out=16'h0;
17'hced:	data_out=16'h0;
17'hcee:	data_out=16'h0;
17'hcef:	data_out=16'h0;
17'hcf0:	data_out=16'h0;
17'hcf1:	data_out=16'h0;
17'hcf2:	data_out=16'h0;
17'hcf3:	data_out=16'h0;
17'hcf4:	data_out=16'h0;
17'hcf5:	data_out=16'h0;
17'hcf6:	data_out=16'h0;
17'hcf7:	data_out=16'h0;
17'hcf8:	data_out=16'h0;
17'hcf9:	data_out=16'h0;
17'hcfa:	data_out=16'h0;
17'hcfb:	data_out=16'h0;
17'hcfc:	data_out=16'h0;
17'hcfd:	data_out=16'h0;
17'hcfe:	data_out=16'h0;
17'hcff:	data_out=16'h0;
17'hd00:	data_out=16'h0;
17'hd01:	data_out=16'h0;
17'hd02:	data_out=16'h0;
17'hd03:	data_out=16'h0;
17'hd04:	data_out=16'h0;
17'hd05:	data_out=16'h0;
17'hd06:	data_out=16'h0;
17'hd07:	data_out=16'h0;
17'hd08:	data_out=16'h0;
17'hd09:	data_out=16'h0;
17'hd0a:	data_out=16'h0;
17'hd0b:	data_out=16'h0;
17'hd0c:	data_out=16'h0;
17'hd0d:	data_out=16'h0;
17'hd0e:	data_out=16'h0;
17'hd0f:	data_out=16'h0;
17'hd10:	data_out=16'h37;
17'hd11:	data_out=16'h95;
17'hd12:	data_out=16'hd3;
17'hd13:	data_out=16'hfe;
17'hd14:	data_out=16'hfe;
17'hd15:	data_out=16'h71;
17'hd16:	data_out=16'h57;
17'hd17:	data_out=16'h95;
17'hd18:	data_out=16'h37;
17'hd19:	data_out=16'h0;
17'hd1a:	data_out=16'h0;
17'hd1b:	data_out=16'h0;
17'hd1c:	data_out=16'h0;
17'hd1d:	data_out=16'h0;
17'hd1e:	data_out=16'h0;
17'hd1f:	data_out=16'h0;
17'hd20:	data_out=16'h0;
17'hd21:	data_out=16'h0;
17'hd22:	data_out=16'h0;
17'hd23:	data_out=16'h0;
17'hd24:	data_out=16'h0;
17'hd25:	data_out=16'h0;
17'hd26:	data_out=16'h0;
17'hd27:	data_out=16'h0;
17'hd28:	data_out=16'h0;
17'hd29:	data_out=16'h0;
17'hd2a:	data_out=16'h0;
17'hd2b:	data_out=16'h57;
17'hd2c:	data_out=16'he9;
17'hd2d:	data_out=16'hfd;
17'hd2e:	data_out=16'hfe;
17'hd2f:	data_out=16'hbe;
17'hd30:	data_out=16'hd3;
17'hd31:	data_out=16'hfd;
17'hd32:	data_out=16'hfd;
17'hd33:	data_out=16'hfe;
17'hd34:	data_out=16'ha9;
17'hd35:	data_out=16'h0;
17'hd36:	data_out=16'h0;
17'hd37:	data_out=16'h0;
17'hd38:	data_out=16'h0;
17'hd39:	data_out=16'h0;
17'hd3a:	data_out=16'h0;
17'hd3b:	data_out=16'h0;
17'hd3c:	data_out=16'h0;
17'hd3d:	data_out=16'h0;
17'hd3e:	data_out=16'h0;
17'hd3f:	data_out=16'h0;
17'hd40:	data_out=16'h0;
17'hd41:	data_out=16'h0;
17'hd42:	data_out=16'h0;
17'hd43:	data_out=16'h0;
17'hd44:	data_out=16'h0;
17'hd45:	data_out=16'h4;
17'hd46:	data_out=16'h39;
17'hd47:	data_out=16'hf3;
17'hd48:	data_out=16'hfd;
17'hd49:	data_out=16'hbf;
17'hd4a:	data_out=16'h41;
17'hd4b:	data_out=16'h5;
17'hd4c:	data_out=16'hc;
17'hd4d:	data_out=16'hb7;
17'hd4e:	data_out=16'hfd;
17'hd4f:	data_out=16'hfe;
17'hd50:	data_out=16'h74;
17'hd51:	data_out=16'h0;
17'hd52:	data_out=16'h0;
17'hd53:	data_out=16'h0;
17'hd54:	data_out=16'h0;
17'hd55:	data_out=16'h0;
17'hd56:	data_out=16'h0;
17'hd57:	data_out=16'h0;
17'hd58:	data_out=16'h0;
17'hd59:	data_out=16'h0;
17'hd5a:	data_out=16'h0;
17'hd5b:	data_out=16'h0;
17'hd5c:	data_out=16'h0;
17'hd5d:	data_out=16'h0;
17'hd5e:	data_out=16'h0;
17'hd5f:	data_out=16'h0;
17'hd60:	data_out=16'h0;
17'hd61:	data_out=16'h60;
17'hd62:	data_out=16'hfd;
17'hd63:	data_out=16'hfd;
17'hd64:	data_out=16'hb8;
17'hd65:	data_out=16'he;
17'hd66:	data_out=16'h0;
17'hd67:	data_out=16'h0;
17'hd68:	data_out=16'h5c;
17'hd69:	data_out=16'hfd;
17'hd6a:	data_out=16'hfd;
17'hd6b:	data_out=16'he2;
17'hd6c:	data_out=16'h15;
17'hd6d:	data_out=16'h0;
17'hd6e:	data_out=16'h0;
17'hd6f:	data_out=16'h0;
17'hd70:	data_out=16'h0;
17'hd71:	data_out=16'h0;
17'hd72:	data_out=16'h0;
17'hd73:	data_out=16'h0;
17'hd74:	data_out=16'h0;
17'hd75:	data_out=16'h0;
17'hd76:	data_out=16'h0;
17'hd77:	data_out=16'h0;
17'hd78:	data_out=16'h0;
17'hd79:	data_out=16'h0;
17'hd7a:	data_out=16'h0;
17'hd7b:	data_out=16'h0;
17'hd7c:	data_out=16'h85;
17'hd7d:	data_out=16'hfe;
17'hd7e:	data_out=16'hfd;
17'hd7f:	data_out=16'h93;
17'hd80:	data_out=16'he;
17'hd81:	data_out=16'h0;
17'hd82:	data_out=16'h0;
17'hd83:	data_out=16'h0;
17'hd84:	data_out=16'hd8;
17'hd85:	data_out=16'hfd;
17'hd86:	data_out=16'hfd;
17'hd87:	data_out=16'h4f;
17'hd88:	data_out=16'h0;
17'hd89:	data_out=16'h0;
17'hd8a:	data_out=16'h0;
17'hd8b:	data_out=16'h0;
17'hd8c:	data_out=16'h0;
17'hd8d:	data_out=16'h0;
17'hd8e:	data_out=16'h0;
17'hd8f:	data_out=16'h0;
17'hd90:	data_out=16'h0;
17'hd91:	data_out=16'h0;
17'hd92:	data_out=16'h0;
17'hd93:	data_out=16'h0;
17'hd94:	data_out=16'h0;
17'hd95:	data_out=16'h0;
17'hd96:	data_out=16'h0;
17'hd97:	data_out=16'h7e;
17'hd98:	data_out=16'hfe;
17'hd99:	data_out=16'hf8;
17'hd9a:	data_out=16'hb1;
17'hd9b:	data_out=16'h9;
17'hd9c:	data_out=16'h0;
17'hd9d:	data_out=16'h0;
17'hd9e:	data_out=16'h8;
17'hd9f:	data_out=16'h4e;
17'hda0:	data_out=16'hf6;
17'hda1:	data_out=16'hfe;
17'hda2:	data_out=16'h82;
17'hda3:	data_out=16'h0;
17'hda4:	data_out=16'h0;
17'hda5:	data_out=16'h0;
17'hda6:	data_out=16'h0;
17'hda7:	data_out=16'h0;
17'hda8:	data_out=16'h0;
17'hda9:	data_out=16'h0;
17'hdaa:	data_out=16'h0;
17'hdab:	data_out=16'h0;
17'hdac:	data_out=16'h0;
17'hdad:	data_out=16'h0;
17'hdae:	data_out=16'h0;
17'hdaf:	data_out=16'h0;
17'hdb0:	data_out=16'h0;
17'hdb1:	data_out=16'h0;
17'hdb2:	data_out=16'h10;
17'hdb3:	data_out=16'he9;
17'hdb4:	data_out=16'hfd;
17'hdb5:	data_out=16'hb1;
17'hdb6:	data_out=16'h0;
17'hdb7:	data_out=16'h0;
17'hdb8:	data_out=16'h0;
17'hdb9:	data_out=16'h24;
17'hdba:	data_out=16'hca;
17'hdbb:	data_out=16'hfd;
17'hdbc:	data_out=16'hfd;
17'hdbd:	data_out=16'haa;
17'hdbe:	data_out=16'hb;
17'hdbf:	data_out=16'h0;
17'hdc0:	data_out=16'h0;
17'hdc1:	data_out=16'h0;
17'hdc2:	data_out=16'h0;
17'hdc3:	data_out=16'h0;
17'hdc4:	data_out=16'h0;
17'hdc5:	data_out=16'h0;
17'hdc6:	data_out=16'h0;
17'hdc7:	data_out=16'h0;
17'hdc8:	data_out=16'h0;
17'hdc9:	data_out=16'h0;
17'hdca:	data_out=16'h0;
17'hdcb:	data_out=16'h0;
17'hdcc:	data_out=16'h0;
17'hdcd:	data_out=16'h0;
17'hdce:	data_out=16'h16;
17'hdcf:	data_out=16'hfd;
17'hdd0:	data_out=16'hfd;
17'hdd1:	data_out=16'h1e;
17'hdd2:	data_out=16'h16;
17'hdd3:	data_out=16'h77;
17'hdd4:	data_out=16'hc6;
17'hdd5:	data_out=16'hf2;
17'hdd6:	data_out=16'hfe;
17'hdd7:	data_out=16'hfd;
17'hdd8:	data_out=16'hfc;
17'hdd9:	data_out=16'h4d;
17'hdda:	data_out=16'h0;
17'hddb:	data_out=16'h0;
17'hddc:	data_out=16'h0;
17'hddd:	data_out=16'h0;
17'hdde:	data_out=16'h0;
17'hddf:	data_out=16'h0;
17'hde0:	data_out=16'h0;
17'hde1:	data_out=16'h0;
17'hde2:	data_out=16'h0;
17'hde3:	data_out=16'h0;
17'hde4:	data_out=16'h0;
17'hde5:	data_out=16'h0;
17'hde6:	data_out=16'h0;
17'hde7:	data_out=16'h0;
17'hde8:	data_out=16'h0;
17'hde9:	data_out=16'h0;
17'hdea:	data_out=16'h10;
17'hdeb:	data_out=16'he8;
17'hdec:	data_out=16'hfd;
17'hded:	data_out=16'hfe;
17'hdee:	data_out=16'hfd;
17'hdef:	data_out=16'hfd;
17'hdf0:	data_out=16'hfd;
17'hdf1:	data_out=16'he3;
17'hdf2:	data_out=16'he4;
17'hdf3:	data_out=16'hfd;
17'hdf4:	data_out=16'he8;
17'hdf5:	data_out=16'h0;
17'hdf6:	data_out=16'h0;
17'hdf7:	data_out=16'h0;
17'hdf8:	data_out=16'h0;
17'hdf9:	data_out=16'h0;
17'hdfa:	data_out=16'h0;
17'hdfb:	data_out=16'h0;
17'hdfc:	data_out=16'h0;
17'hdfd:	data_out=16'h0;
17'hdfe:	data_out=16'h0;
17'hdff:	data_out=16'h0;
17'he00:	data_out=16'h0;
17'he01:	data_out=16'h0;
17'he02:	data_out=16'h0;
17'he03:	data_out=16'h0;
17'he04:	data_out=16'h0;
17'he05:	data_out=16'h0;
17'he06:	data_out=16'h0;
17'he07:	data_out=16'h37;
17'he08:	data_out=16'hec;
17'he09:	data_out=16'hfe;
17'he0a:	data_out=16'hda;
17'he0b:	data_out=16'h8b;
17'he0c:	data_out=16'h2a;
17'he0d:	data_out=16'h18;
17'he0e:	data_out=16'hc1;
17'he0f:	data_out=16'hfd;
17'he10:	data_out=16'h90;
17'he11:	data_out=16'h0;
17'he12:	data_out=16'h0;
17'he13:	data_out=16'h0;
17'he14:	data_out=16'h0;
17'he15:	data_out=16'h0;
17'he16:	data_out=16'h0;
17'he17:	data_out=16'h0;
17'he18:	data_out=16'h0;
17'he19:	data_out=16'h0;
17'he1a:	data_out=16'h0;
17'he1b:	data_out=16'h0;
17'he1c:	data_out=16'h0;
17'he1d:	data_out=16'h0;
17'he1e:	data_out=16'h0;
17'he1f:	data_out=16'h0;
17'he20:	data_out=16'h0;
17'he21:	data_out=16'h0;
17'he22:	data_out=16'h0;
17'he23:	data_out=16'h0;
17'he24:	data_out=16'h0;
17'he25:	data_out=16'h0;
17'he26:	data_out=16'h0;
17'he27:	data_out=16'h0;
17'he28:	data_out=16'h0;
17'he29:	data_out=16'h3e;
17'he2a:	data_out=16'h100;
17'he2b:	data_out=16'hfe;
17'he2c:	data_out=16'h6d;
17'he2d:	data_out=16'h0;
17'he2e:	data_out=16'h0;
17'he2f:	data_out=16'h0;
17'he30:	data_out=16'h0;
17'he31:	data_out=16'h0;
17'he32:	data_out=16'h0;
17'he33:	data_out=16'h0;
17'he34:	data_out=16'h0;
17'he35:	data_out=16'h0;
17'he36:	data_out=16'h0;
17'he37:	data_out=16'h0;
17'he38:	data_out=16'h0;
17'he39:	data_out=16'h0;
17'he3a:	data_out=16'h0;
17'he3b:	data_out=16'h0;
17'he3c:	data_out=16'h0;
17'he3d:	data_out=16'h0;
17'he3e:	data_out=16'h0;
17'he3f:	data_out=16'h0;
17'he40:	data_out=16'h0;
17'he41:	data_out=16'h0;
17'he42:	data_out=16'h0;
17'he43:	data_out=16'h0;
17'he44:	data_out=16'h0;
17'he45:	data_out=16'h47;
17'he46:	data_out=16'hfe;
17'he47:	data_out=16'hfd;
17'he48:	data_out=16'h15;
17'he49:	data_out=16'h0;
17'he4a:	data_out=16'h0;
17'he4b:	data_out=16'h0;
17'he4c:	data_out=16'h0;
17'he4d:	data_out=16'h0;
17'he4e:	data_out=16'h0;
17'he4f:	data_out=16'h0;
17'he50:	data_out=16'h0;
17'he51:	data_out=16'h0;
17'he52:	data_out=16'h0;
17'he53:	data_out=16'h0;
17'he54:	data_out=16'h0;
17'he55:	data_out=16'h0;
17'he56:	data_out=16'h0;
17'he57:	data_out=16'h0;
17'he58:	data_out=16'h0;
17'he59:	data_out=16'h0;
17'he5a:	data_out=16'h0;
17'he5b:	data_out=16'h0;
17'he5c:	data_out=16'h0;
17'he5d:	data_out=16'h0;
17'he5e:	data_out=16'h0;
17'he5f:	data_out=16'h0;
17'he60:	data_out=16'h0;
17'he61:	data_out=16'h0;
17'he62:	data_out=16'hfe;
17'he63:	data_out=16'hfd;
17'he64:	data_out=16'h15;
17'he65:	data_out=16'h0;
17'he66:	data_out=16'h0;
17'he67:	data_out=16'h0;
17'he68:	data_out=16'h0;
17'he69:	data_out=16'h0;
17'he6a:	data_out=16'h0;
17'he6b:	data_out=16'h0;
17'he6c:	data_out=16'h0;
17'he6d:	data_out=16'h0;
17'he6e:	data_out=16'h0;
17'he6f:	data_out=16'h0;
17'he70:	data_out=16'h0;
17'he71:	data_out=16'h0;
17'he72:	data_out=16'h0;
17'he73:	data_out=16'h0;
17'he74:	data_out=16'h0;
17'he75:	data_out=16'h0;
17'he76:	data_out=16'h0;
17'he77:	data_out=16'h0;
17'he78:	data_out=16'h0;
17'he79:	data_out=16'h0;
17'he7a:	data_out=16'h0;
17'he7b:	data_out=16'h0;
17'he7c:	data_out=16'h0;
17'he7d:	data_out=16'h47;
17'he7e:	data_out=16'hfe;
17'he7f:	data_out=16'hfd;
17'he80:	data_out=16'h15;
17'he81:	data_out=16'h0;
17'he82:	data_out=16'h0;
17'he83:	data_out=16'h0;
17'he84:	data_out=16'h0;
17'he85:	data_out=16'h0;
17'he86:	data_out=16'h0;
17'he87:	data_out=16'h0;
17'he88:	data_out=16'h0;
17'he89:	data_out=16'h0;
17'he8a:	data_out=16'h0;
17'he8b:	data_out=16'h0;
17'he8c:	data_out=16'h0;
17'he8d:	data_out=16'h0;
17'he8e:	data_out=16'h0;
17'he8f:	data_out=16'h0;
17'he90:	data_out=16'h0;
17'he91:	data_out=16'h0;
17'he92:	data_out=16'h0;
17'he93:	data_out=16'h0;
17'he94:	data_out=16'h0;
17'he95:	data_out=16'h0;
17'he96:	data_out=16'h0;
17'he97:	data_out=16'h0;
17'he98:	data_out=16'h0;
17'he99:	data_out=16'h6a;
17'he9a:	data_out=16'hfe;
17'he9b:	data_out=16'hfd;
17'he9c:	data_out=16'h15;
17'he9d:	data_out=16'h0;
17'he9e:	data_out=16'h0;
17'he9f:	data_out=16'h0;
17'hea0:	data_out=16'h0;
17'hea1:	data_out=16'h0;
17'hea2:	data_out=16'h0;
17'hea3:	data_out=16'h0;
17'hea4:	data_out=16'h0;
17'hea5:	data_out=16'h0;
17'hea6:	data_out=16'h0;
17'hea7:	data_out=16'h0;
17'hea8:	data_out=16'h0;
17'hea9:	data_out=16'h0;
17'heaa:	data_out=16'h0;
17'heab:	data_out=16'h0;
17'heac:	data_out=16'h0;
17'head:	data_out=16'h0;
17'heae:	data_out=16'h0;
17'heaf:	data_out=16'h0;
17'heb0:	data_out=16'h0;
17'heb1:	data_out=16'h0;
17'heb2:	data_out=16'h0;
17'heb3:	data_out=16'h0;
17'heb4:	data_out=16'h0;
17'heb5:	data_out=16'h2d;
17'heb6:	data_out=16'h100;
17'heb7:	data_out=16'hfe;
17'heb8:	data_out=16'h15;
17'heb9:	data_out=16'h0;
17'heba:	data_out=16'h0;
17'hebb:	data_out=16'h0;
17'hebc:	data_out=16'h0;
17'hebd:	data_out=16'h0;
17'hebe:	data_out=16'h0;
17'hebf:	data_out=16'h0;
17'hec0:	data_out=16'h0;
17'hec1:	data_out=16'h0;
17'hec2:	data_out=16'h0;
17'hec3:	data_out=16'h0;
17'hec4:	data_out=16'h0;
17'hec5:	data_out=16'h0;
17'hec6:	data_out=16'h0;
17'hec7:	data_out=16'h0;
17'hec8:	data_out=16'h0;
17'hec9:	data_out=16'h0;
17'heca:	data_out=16'h0;
17'hecb:	data_out=16'h0;
17'hecc:	data_out=16'h0;
17'hecd:	data_out=16'h0;
17'hece:	data_out=16'h0;
17'hecf:	data_out=16'h0;
17'hed0:	data_out=16'h0;
17'hed1:	data_out=16'h0;
17'hed2:	data_out=16'hdb;
17'hed3:	data_out=16'hfd;
17'hed4:	data_out=16'h38;
17'hed5:	data_out=16'h0;
17'hed6:	data_out=16'h0;
17'hed7:	data_out=16'h0;
17'hed8:	data_out=16'h0;
17'hed9:	data_out=16'h0;
17'heda:	data_out=16'h0;
17'hedb:	data_out=16'h0;
17'hedc:	data_out=16'h0;
17'hedd:	data_out=16'h0;
17'hede:	data_out=16'h0;
17'hedf:	data_out=16'h0;
17'hee0:	data_out=16'h0;
17'hee1:	data_out=16'h0;
17'hee2:	data_out=16'h0;
17'hee3:	data_out=16'h0;
17'hee4:	data_out=16'h0;
17'hee5:	data_out=16'h0;
17'hee6:	data_out=16'h0;
17'hee7:	data_out=16'h0;
17'hee8:	data_out=16'h0;
17'hee9:	data_out=16'h0;
17'heea:	data_out=16'h0;
17'heeb:	data_out=16'h0;
17'heec:	data_out=16'h0;
17'heed:	data_out=16'h0;
17'heee:	data_out=16'h60;
17'heef:	data_out=16'hfd;
17'hef0:	data_out=16'hbe;
17'hef1:	data_out=16'h2a;
17'hef2:	data_out=16'h0;
17'hef3:	data_out=16'h0;
17'hef4:	data_out=16'h0;
17'hef5:	data_out=16'h0;
17'hef6:	data_out=16'h0;
17'hef7:	data_out=16'h0;
17'hef8:	data_out=16'h0;
17'hef9:	data_out=16'h0;
17'hefa:	data_out=16'h0;
17'hefb:	data_out=16'h0;
17'hefc:	data_out=16'h0;
17'hefd:	data_out=16'h0;
17'hefe:	data_out=16'h0;
17'heff:	data_out=16'h0;
17'hf00:	data_out=16'h0;
17'hf01:	data_out=16'h0;
17'hf02:	data_out=16'h0;
17'hf03:	data_out=16'h0;
17'hf04:	data_out=16'h0;
17'hf05:	data_out=16'h0;
17'hf06:	data_out=16'h0;
17'hf07:	data_out=16'h0;
17'hf08:	data_out=16'h0;
17'hf09:	data_out=16'h0;
17'hf0a:	data_out=16'he;
17'hf0b:	data_out=16'hb9;
17'hf0c:	data_out=16'hfd;
17'hf0d:	data_out=16'hab;
17'hf0e:	data_out=16'hb;
17'hf0f:	data_out=16'h0;
17'hf10:	data_out=16'h0;
17'hf11:	data_out=16'h0;
17'hf12:	data_out=16'h0;
17'hf13:	data_out=16'h0;
17'hf14:	data_out=16'h0;
17'hf15:	data_out=16'h0;
17'hf16:	data_out=16'h0;
17'hf17:	data_out=16'h0;
17'hf18:	data_out=16'h0;
17'hf19:	data_out=16'h0;
17'hf1a:	data_out=16'h0;
17'hf1b:	data_out=16'h0;
17'hf1c:	data_out=16'h0;
17'hf1d:	data_out=16'h0;
17'hf1e:	data_out=16'h0;
17'hf1f:	data_out=16'h0;
17'hf20:	data_out=16'h0;
17'hf21:	data_out=16'h0;
17'hf22:	data_out=16'h0;
17'hf23:	data_out=16'h0;
17'hf24:	data_out=16'h0;
17'hf25:	data_out=16'h0;
17'hf26:	data_out=16'h0;
17'hf27:	data_out=16'he;
17'hf28:	data_out=16'h94;
17'hf29:	data_out=16'hfd;
17'hf2a:	data_out=16'h2a;
17'hf2b:	data_out=16'h0;
17'hf2c:	data_out=16'h0;
17'hf2d:	data_out=16'h0;
17'hf2e:	data_out=16'h0;
17'hf2f:	data_out=16'h0;
17'hf30:	data_out=16'h0;
17'hf31:	data_out=16'h0;
17'hf32:	data_out=16'h0;
17'hf33:	data_out=16'h0;
17'hf34:	data_out=16'h0;
17'hf35:	data_out=16'h0;
17'hf36:	data_out=16'h0;
17'hf37:	data_out=16'h0;
17'hf38:	data_out=16'h0;
17'hf39:	data_out=16'h0;
17'hf3a:	data_out=16'h0;
17'hf3b:	data_out=16'h0;
17'hf3c:	data_out=16'h0;
17'hf3d:	data_out=16'h0;
17'hf3e:	data_out=16'h0;
17'hf3f:	data_out=16'h0;
17'hf40:	data_out=16'h0;
17'hf41:	data_out=16'h0;
17'hf42:	data_out=16'h0;
17'hf43:	data_out=16'h0;
17'hf44:	data_out=16'h0;
17'hf45:	data_out=16'h0;
17'hf46:	data_out=16'h0;
17'hf47:	data_out=16'h0;
17'hf48:	data_out=16'h0;
17'hf49:	data_out=16'h0;
17'hf4a:	data_out=16'h0;
17'hf4b:	data_out=16'h0;
17'hf4c:	data_out=16'h0;
17'hf4d:	data_out=16'h0;
17'hf4e:	data_out=16'h0;
17'hf4f:	data_out=16'h0;
17'hf50:	data_out=16'h0;
17'hf51:	data_out=16'h0;
17'hf52:	data_out=16'h0;
17'hf53:	data_out=16'h0;
17'hf54:	data_out=16'h0;
17'hf55:	data_out=16'h0;
17'hf56:	data_out=16'h0;
17'hf57:	data_out=16'h0;
17'hf58:	data_out=16'h0;
17'hf59:	data_out=16'h0;
17'hf5a:	data_out=16'h0;
17'hf5b:	data_out=16'h0;
17'hf5c:	data_out=16'h0;
17'hf5d:	data_out=16'h0;
17'hf5e:	data_out=16'h0;
17'hf5f:	data_out=16'h0;
17'hf60:	data_out=16'h0;
17'hf61:	data_out=16'h0;
17'hf62:	data_out=16'h0;
17'hf63:	data_out=16'h0;
17'hf64:	data_out=16'h0;
17'hf65:	data_out=16'h0;
17'hf66:	data_out=16'h0;
17'hf67:	data_out=16'h0;
17'hf68:	data_out=16'h0;
17'hf69:	data_out=16'h0;
17'hf6a:	data_out=16'h0;
17'hf6b:	data_out=16'h0;
17'hf6c:	data_out=16'h0;
17'hf6d:	data_out=16'h0;
17'hf6e:	data_out=16'h0;
17'hf6f:	data_out=16'h0;
17'hf70:	data_out=16'h0;
17'hf71:	data_out=16'h0;
17'hf72:	data_out=16'h0;
17'hf73:	data_out=16'h0;
17'hf74:	data_out=16'h0;
17'hf75:	data_out=16'h0;
17'hf76:	data_out=16'h0;
17'hf77:	data_out=16'h0;
17'hf78:	data_out=16'h0;
17'hf79:	data_out=16'h0;
17'hf7a:	data_out=16'h0;
17'hf7b:	data_out=16'h0;
17'hf7c:	data_out=16'h0;
17'hf7d:	data_out=16'h0;
17'hf7e:	data_out=16'h0;
17'hf7f:	data_out=16'h0;
17'hf80:	data_out=16'h0;
17'hf81:	data_out=16'h0;
17'hf82:	data_out=16'h0;
17'hf83:	data_out=16'h0;
17'hf84:	data_out=16'h0;
17'hf85:	data_out=16'h0;
17'hf86:	data_out=16'h0;
17'hf87:	data_out=16'h0;
17'hf88:	data_out=16'h0;
17'hf89:	data_out=16'h0;
17'hf8a:	data_out=16'h0;
17'hf8b:	data_out=16'h0;
17'hf8c:	data_out=16'h0;
17'hf8d:	data_out=16'h0;
17'hf8e:	data_out=16'h0;
17'hf8f:	data_out=16'h0;
17'hf90:	data_out=16'h0;
17'hf91:	data_out=16'h0;
17'hf92:	data_out=16'h0;
17'hf93:	data_out=16'h0;
17'hf94:	data_out=16'h0;
17'hf95:	data_out=16'h0;
17'hf96:	data_out=16'h0;
17'hf97:	data_out=16'h0;
17'hf98:	data_out=16'h0;
17'hf99:	data_out=16'h0;
17'hf9a:	data_out=16'h0;
17'hf9b:	data_out=16'h0;
17'hf9c:	data_out=16'h0;
17'hf9d:	data_out=16'h0;
17'hf9e:	data_out=16'h0;
17'hf9f:	data_out=16'h0;
17'hfa0:	data_out=16'h0;
17'hfa1:	data_out=16'h0;
17'hfa2:	data_out=16'h0;
17'hfa3:	data_out=16'h0;
17'hfa4:	data_out=16'h0;
17'hfa5:	data_out=16'h0;
17'hfa6:	data_out=16'h0;
17'hfa7:	data_out=16'h0;
17'hfa8:	data_out=16'h0;
17'hfa9:	data_out=16'h0;
17'hfaa:	data_out=16'h0;
17'hfab:	data_out=16'h0;
17'hfac:	data_out=16'h0;
17'hfad:	data_out=16'h0;
17'hfae:	data_out=16'h0;
17'hfaf:	data_out=16'h0;
17'hfb0:	data_out=16'h0;
17'hfb1:	data_out=16'h0;
17'hfb2:	data_out=16'h0;
17'hfb3:	data_out=16'h0;
17'hfb4:	data_out=16'h0;
17'hfb5:	data_out=16'h0;
17'hfb6:	data_out=16'h0;
17'hfb7:	data_out=16'h0;
17'hfb8:	data_out=16'h0;
17'hfb9:	data_out=16'h0;
17'hfba:	data_out=16'h0;
17'hfbb:	data_out=16'h0;
17'hfbc:	data_out=16'h0;
17'hfbd:	data_out=16'h0;
17'hfbe:	data_out=16'h0;
17'hfbf:	data_out=16'h0;
17'hfc0:	data_out=16'h0;
17'hfc1:	data_out=16'h0;
17'hfc2:	data_out=16'h0;
17'hfc3:	data_out=16'h0;
17'hfc4:	data_out=16'h0;
17'hfc5:	data_out=16'h0;
17'hfc6:	data_out=16'h0;
17'hfc7:	data_out=16'h0;
17'hfc8:	data_out=16'h0;
17'hfc9:	data_out=16'h0;
17'hfca:	data_out=16'h0;
17'hfcb:	data_out=16'h0;
17'hfcc:	data_out=16'h0;
17'hfcd:	data_out=16'h0;
17'hfce:	data_out=16'h0;
17'hfcf:	data_out=16'h0;
17'hfd0:	data_out=16'h0;
17'hfd1:	data_out=16'h0;
17'hfd2:	data_out=16'h0;
17'hfd3:	data_out=16'h0;
17'hfd4:	data_out=16'h0;
17'hfd5:	data_out=16'h0;
17'hfd6:	data_out=16'h0;
17'hfd7:	data_out=16'h0;
17'hfd8:	data_out=16'h0;
17'hfd9:	data_out=16'h0;
17'hfda:	data_out=16'h0;
17'hfdb:	data_out=16'h0;
17'hfdc:	data_out=16'h0;
17'hfdd:	data_out=16'h0;
17'hfde:	data_out=16'h0;
17'hfdf:	data_out=16'h0;
17'hfe0:	data_out=16'h0;
17'hfe1:	data_out=16'h0;
17'hfe2:	data_out=16'h0;
17'hfe3:	data_out=16'h0;
17'hfe4:	data_out=16'h0;
17'hfe5:	data_out=16'h0;
17'hfe6:	data_out=16'h0;
17'hfe7:	data_out=16'h0;
17'hfe8:	data_out=16'h0;
17'hfe9:	data_out=16'h0;
17'hfea:	data_out=16'h0;
17'hfeb:	data_out=16'hd;
17'hfec:	data_out=16'h19;
17'hfed:	data_out=16'h64;
17'hfee:	data_out=16'h7a;
17'hfef:	data_out=16'h7;
17'hff0:	data_out=16'h0;
17'hff1:	data_out=16'h0;
17'hff2:	data_out=16'h0;
17'hff3:	data_out=16'h0;
17'hff4:	data_out=16'h0;
17'hff5:	data_out=16'h0;
17'hff6:	data_out=16'h0;
17'hff7:	data_out=16'h0;
17'hff8:	data_out=16'h0;
17'hff9:	data_out=16'h0;
17'hffa:	data_out=16'h0;
17'hffb:	data_out=16'h0;
17'hffc:	data_out=16'h0;
17'hffd:	data_out=16'h0;
17'hffe:	data_out=16'h0;
17'hfff:	data_out=16'h0;
17'h1000:	data_out=16'h0;
17'h1001:	data_out=16'h0;
17'h1002:	data_out=16'h0;
17'h1003:	data_out=16'h0;
17'h1004:	data_out=16'h0;
17'h1005:	data_out=16'h21;
17'h1006:	data_out=16'h98;
17'h1007:	data_out=16'hd1;
17'h1008:	data_out=16'hfd;
17'h1009:	data_out=16'hfd;
17'h100a:	data_out=16'hfd;
17'h100b:	data_out=16'h93;
17'h100c:	data_out=16'h0;
17'h100d:	data_out=16'h0;
17'h100e:	data_out=16'h0;
17'h100f:	data_out=16'h0;
17'h1010:	data_out=16'h0;
17'h1011:	data_out=16'h0;
17'h1012:	data_out=16'h0;
17'h1013:	data_out=16'h0;
17'h1014:	data_out=16'h0;
17'h1015:	data_out=16'h0;
17'h1016:	data_out=16'h0;
17'h1017:	data_out=16'h0;
17'h1018:	data_out=16'h0;
17'h1019:	data_out=16'h0;
17'h101a:	data_out=16'h0;
17'h101b:	data_out=16'h0;
17'h101c:	data_out=16'h0;
17'h101d:	data_out=16'h0;
17'h101e:	data_out=16'h0;
17'h101f:	data_out=16'h28;
17'h1020:	data_out=16'h99;
17'h1021:	data_out=16'hf5;
17'h1022:	data_out=16'hfd;
17'h1023:	data_out=16'hfe;
17'h1024:	data_out=16'he1;
17'h1025:	data_out=16'hd4;
17'h1026:	data_out=16'hfd;
17'h1027:	data_out=16'he9;
17'h1028:	data_out=16'h28;
17'h1029:	data_out=16'h0;
17'h102a:	data_out=16'h0;
17'h102b:	data_out=16'h0;
17'h102c:	data_out=16'h0;
17'h102d:	data_out=16'h0;
17'h102e:	data_out=16'h0;
17'h102f:	data_out=16'h0;
17'h1030:	data_out=16'h0;
17'h1031:	data_out=16'h0;
17'h1032:	data_out=16'h0;
17'h1033:	data_out=16'h0;
17'h1034:	data_out=16'h0;
17'h1035:	data_out=16'h0;
17'h1036:	data_out=16'h0;
17'h1037:	data_out=16'h0;
17'h1038:	data_out=16'h0;
17'h1039:	data_out=16'hf;
17'h103a:	data_out=16'h99;
17'h103b:	data_out=16'hf0;
17'h103c:	data_out=16'hfd;
17'h103d:	data_out=16'hfd;
17'h103e:	data_out=16'hfd;
17'h103f:	data_out=16'hd9;
17'h1040:	data_out=16'h1f;
17'h1041:	data_out=16'h25;
17'h1042:	data_out=16'hfd;
17'h1043:	data_out=16'hfd;
17'h1044:	data_out=16'h3c;
17'h1045:	data_out=16'h0;
17'h1046:	data_out=16'h0;
17'h1047:	data_out=16'h0;
17'h1048:	data_out=16'h0;
17'h1049:	data_out=16'h0;
17'h104a:	data_out=16'h0;
17'h104b:	data_out=16'h0;
17'h104c:	data_out=16'h0;
17'h104d:	data_out=16'h0;
17'h104e:	data_out=16'h0;
17'h104f:	data_out=16'h0;
17'h1050:	data_out=16'h0;
17'h1051:	data_out=16'h0;
17'h1052:	data_out=16'h0;
17'h1053:	data_out=16'h0;
17'h1054:	data_out=16'h0;
17'h1055:	data_out=16'h60;
17'h1056:	data_out=16'hfd;
17'h1057:	data_out=16'hfd;
17'h1058:	data_out=16'hfd;
17'h1059:	data_out=16'hfd;
17'h105a:	data_out=16'hda;
17'h105b:	data_out=16'h1d;
17'h105c:	data_out=16'h0;
17'h105d:	data_out=16'h25;
17'h105e:	data_out=16'hfd;
17'h105f:	data_out=16'hfd;
17'h1060:	data_out=16'h3c;
17'h1061:	data_out=16'h0;
17'h1062:	data_out=16'h0;
17'h1063:	data_out=16'h0;
17'h1064:	data_out=16'h0;
17'h1065:	data_out=16'h0;
17'h1066:	data_out=16'h0;
17'h1067:	data_out=16'h0;
17'h1068:	data_out=16'h0;
17'h1069:	data_out=16'h0;
17'h106a:	data_out=16'h0;
17'h106b:	data_out=16'h0;
17'h106c:	data_out=16'h0;
17'h106d:	data_out=16'h0;
17'h106e:	data_out=16'h0;
17'h106f:	data_out=16'h0;
17'h1070:	data_out=16'h0;
17'h1071:	data_out=16'hb6;
17'h1072:	data_out=16'hfd;
17'h1073:	data_out=16'hfd;
17'h1074:	data_out=16'hdd;
17'h1075:	data_out=16'ha8;
17'h1076:	data_out=16'h1e;
17'h1077:	data_out=16'h0;
17'h1078:	data_out=16'h0;
17'h1079:	data_out=16'h4d;
17'h107a:	data_out=16'hfd;
17'h107b:	data_out=16'hfd;
17'h107c:	data_out=16'h3c;
17'h107d:	data_out=16'h0;
17'h107e:	data_out=16'h0;
17'h107f:	data_out=16'h0;
17'h1080:	data_out=16'h0;
17'h1081:	data_out=16'h0;
17'h1082:	data_out=16'h0;
17'h1083:	data_out=16'h0;
17'h1084:	data_out=16'h0;
17'h1085:	data_out=16'h0;
17'h1086:	data_out=16'h0;
17'h1087:	data_out=16'h0;
17'h1088:	data_out=16'h0;
17'h1089:	data_out=16'h0;
17'h108a:	data_out=16'h0;
17'h108b:	data_out=16'h0;
17'h108c:	data_out=16'h0;
17'h108d:	data_out=16'h1a;
17'h108e:	data_out=16'h81;
17'h108f:	data_out=16'h3a;
17'h1090:	data_out=16'h16;
17'h1091:	data_out=16'h0;
17'h1092:	data_out=16'h0;
17'h1093:	data_out=16'h0;
17'h1094:	data_out=16'h0;
17'h1095:	data_out=16'h64;
17'h1096:	data_out=16'hfd;
17'h1097:	data_out=16'hfd;
17'h1098:	data_out=16'h3c;
17'h1099:	data_out=16'h0;
17'h109a:	data_out=16'h0;
17'h109b:	data_out=16'h0;
17'h109c:	data_out=16'h0;
17'h109d:	data_out=16'h0;
17'h109e:	data_out=16'h0;
17'h109f:	data_out=16'h0;
17'h10a0:	data_out=16'h0;
17'h10a1:	data_out=16'h0;
17'h10a2:	data_out=16'h0;
17'h10a3:	data_out=16'h0;
17'h10a4:	data_out=16'h0;
17'h10a5:	data_out=16'h0;
17'h10a6:	data_out=16'h0;
17'h10a7:	data_out=16'h0;
17'h10a8:	data_out=16'h0;
17'h10a9:	data_out=16'h0;
17'h10aa:	data_out=16'h0;
17'h10ab:	data_out=16'h0;
17'h10ac:	data_out=16'h0;
17'h10ad:	data_out=16'h0;
17'h10ae:	data_out=16'h0;
17'h10af:	data_out=16'h0;
17'h10b0:	data_out=16'h0;
17'h10b1:	data_out=16'h9e;
17'h10b2:	data_out=16'hfd;
17'h10b3:	data_out=16'hfd;
17'h10b4:	data_out=16'h3c;
17'h10b5:	data_out=16'h0;
17'h10b6:	data_out=16'h0;
17'h10b7:	data_out=16'h0;
17'h10b8:	data_out=16'h0;
17'h10b9:	data_out=16'h0;
17'h10ba:	data_out=16'h0;
17'h10bb:	data_out=16'h0;
17'h10bc:	data_out=16'h0;
17'h10bd:	data_out=16'h0;
17'h10be:	data_out=16'h0;
17'h10bf:	data_out=16'h0;
17'h10c0:	data_out=16'h0;
17'h10c1:	data_out=16'h0;
17'h10c2:	data_out=16'h0;
17'h10c3:	data_out=16'h0;
17'h10c4:	data_out=16'h0;
17'h10c5:	data_out=16'h0;
17'h10c6:	data_out=16'h0;
17'h10c7:	data_out=16'h0;
17'h10c8:	data_out=16'h0;
17'h10c9:	data_out=16'h6e;
17'h10ca:	data_out=16'h79;
17'h10cb:	data_out=16'h7a;
17'h10cc:	data_out=16'h79;
17'h10cd:	data_out=16'hcb;
17'h10ce:	data_out=16'hfd;
17'h10cf:	data_out=16'hc3;
17'h10d0:	data_out=16'h3;
17'h10d1:	data_out=16'h0;
17'h10d2:	data_out=16'h0;
17'h10d3:	data_out=16'h0;
17'h10d4:	data_out=16'h0;
17'h10d5:	data_out=16'h0;
17'h10d6:	data_out=16'h0;
17'h10d7:	data_out=16'h0;
17'h10d8:	data_out=16'h0;
17'h10d9:	data_out=16'h0;
17'h10da:	data_out=16'h0;
17'h10db:	data_out=16'h0;
17'h10dc:	data_out=16'h0;
17'h10dd:	data_out=16'h0;
17'h10de:	data_out=16'h0;
17'h10df:	data_out=16'h0;
17'h10e0:	data_out=16'h0;
17'h10e1:	data_out=16'h0;
17'h10e2:	data_out=16'ha;
17'h10e3:	data_out=16'h35;
17'h10e4:	data_out=16'hb4;
17'h10e5:	data_out=16'hfe;
17'h10e6:	data_out=16'hfe;
17'h10e7:	data_out=16'h100;
17'h10e8:	data_out=16'hfe;
17'h10e9:	data_out=16'hfe;
17'h10ea:	data_out=16'he5;
17'h10eb:	data_out=16'h23;
17'h10ec:	data_out=16'h0;
17'h10ed:	data_out=16'h0;
17'h10ee:	data_out=16'h0;
17'h10ef:	data_out=16'h0;
17'h10f0:	data_out=16'h0;
17'h10f1:	data_out=16'h0;
17'h10f2:	data_out=16'h0;
17'h10f3:	data_out=16'h0;
17'h10f4:	data_out=16'h0;
17'h10f5:	data_out=16'h0;
17'h10f6:	data_out=16'h0;
17'h10f7:	data_out=16'h0;
17'h10f8:	data_out=16'h0;
17'h10f9:	data_out=16'h0;
17'h10fa:	data_out=16'h0;
17'h10fb:	data_out=16'h0;
17'h10fc:	data_out=16'h5;
17'h10fd:	data_out=16'h36;
17'h10fe:	data_out=16'he4;
17'h10ff:	data_out=16'hfd;
17'h1100:	data_out=16'hf4;
17'h1101:	data_out=16'he5;
17'h1102:	data_out=16'hab;
17'h1103:	data_out=16'hf3;
17'h1104:	data_out=16'hfd;
17'h1105:	data_out=16'hfd;
17'h1106:	data_out=16'he8;
17'h1107:	data_out=16'h75;
17'h1108:	data_out=16'h6;
17'h1109:	data_out=16'h0;
17'h110a:	data_out=16'h0;
17'h110b:	data_out=16'h0;
17'h110c:	data_out=16'h0;
17'h110d:	data_out=16'h0;
17'h110e:	data_out=16'h0;
17'h110f:	data_out=16'h0;
17'h1110:	data_out=16'h0;
17'h1111:	data_out=16'h0;
17'h1112:	data_out=16'h0;
17'h1113:	data_out=16'h0;
17'h1114:	data_out=16'h0;
17'h1115:	data_out=16'h0;
17'h1116:	data_out=16'h0;
17'h1117:	data_out=16'h6;
17'h1118:	data_out=16'h4e;
17'h1119:	data_out=16'hfd;
17'h111a:	data_out=16'hfd;
17'h111b:	data_out=16'h7d;
17'h111c:	data_out=16'h3b;
17'h111d:	data_out=16'h0;
17'h111e:	data_out=16'h12;
17'h111f:	data_out=16'hd1;
17'h1120:	data_out=16'hfd;
17'h1121:	data_out=16'hfd;
17'h1122:	data_out=16'hfd;
17'h1123:	data_out=16'hfd;
17'h1124:	data_out=16'h57;
17'h1125:	data_out=16'h7;
17'h1126:	data_out=16'h0;
17'h1127:	data_out=16'h0;
17'h1128:	data_out=16'h0;
17'h1129:	data_out=16'h0;
17'h112a:	data_out=16'h0;
17'h112b:	data_out=16'h0;
17'h112c:	data_out=16'h0;
17'h112d:	data_out=16'h0;
17'h112e:	data_out=16'h0;
17'h112f:	data_out=16'h0;
17'h1130:	data_out=16'h0;
17'h1131:	data_out=16'h0;
17'h1132:	data_out=16'h5;
17'h1133:	data_out=16'h88;
17'h1134:	data_out=16'hfd;
17'h1135:	data_out=16'hfd;
17'h1136:	data_out=16'hb5;
17'h1137:	data_out=16'h10;
17'h1138:	data_out=16'h0;
17'h1139:	data_out=16'h15;
17'h113a:	data_out=16'hcc;
17'h113b:	data_out=16'hfe;
17'h113c:	data_out=16'hf8;
17'h113d:	data_out=16'h82;
17'h113e:	data_out=16'hae;
17'h113f:	data_out=16'hfd;
17'h1140:	data_out=16'hfd;
17'h1141:	data_out=16'hb9;
17'h1142:	data_out=16'h42;
17'h1143:	data_out=16'h31;
17'h1144:	data_out=16'h31;
17'h1145:	data_out=16'h0;
17'h1146:	data_out=16'h0;
17'h1147:	data_out=16'h0;
17'h1148:	data_out=16'h0;
17'h1149:	data_out=16'h0;
17'h114a:	data_out=16'h0;
17'h114b:	data_out=16'h0;
17'h114c:	data_out=16'h0;
17'h114d:	data_out=16'h3;
17'h114e:	data_out=16'h89;
17'h114f:	data_out=16'hfd;
17'h1150:	data_out=16'hf2;
17'h1151:	data_out=16'h6a;
17'h1152:	data_out=16'h11;
17'h1153:	data_out=16'h0;
17'h1154:	data_out=16'h35;
17'h1155:	data_out=16'hc9;
17'h1156:	data_out=16'hfd;
17'h1157:	data_out=16'hd9;
17'h1158:	data_out=16'h41;
17'h1159:	data_out=16'h0;
17'h115a:	data_out=16'he;
17'h115b:	data_out=16'h48;
17'h115c:	data_out=16'ha4;
17'h115d:	data_out=16'hf2;
17'h115e:	data_out=16'hfd;
17'h115f:	data_out=16'hfd;
17'h1160:	data_out=16'he0;
17'h1161:	data_out=16'h0;
17'h1162:	data_out=16'h0;
17'h1163:	data_out=16'h0;
17'h1164:	data_out=16'h0;
17'h1165:	data_out=16'h0;
17'h1166:	data_out=16'h0;
17'h1167:	data_out=16'h0;
17'h1168:	data_out=16'h0;
17'h1169:	data_out=16'h69;
17'h116a:	data_out=16'hfd;
17'h116b:	data_out=16'hf3;
17'h116c:	data_out=16'h58;
17'h116d:	data_out=16'h12;
17'h116e:	data_out=16'h49;
17'h116f:	data_out=16'hab;
17'h1170:	data_out=16'hf5;
17'h1171:	data_out=16'hfd;
17'h1172:	data_out=16'h7e;
17'h1173:	data_out=16'h1d;
17'h1174:	data_out=16'h0;
17'h1175:	data_out=16'h0;
17'h1176:	data_out=16'h0;
17'h1177:	data_out=16'h0;
17'h1178:	data_out=16'h0;
17'h1179:	data_out=16'h59;
17'h117a:	data_out=16'hb5;
17'h117b:	data_out=16'hb5;
17'h117c:	data_out=16'h25;
17'h117d:	data_out=16'h0;
17'h117e:	data_out=16'h0;
17'h117f:	data_out=16'h0;
17'h1180:	data_out=16'h0;
17'h1181:	data_out=16'h0;
17'h1182:	data_out=16'h0;
17'h1183:	data_out=16'h0;
17'h1184:	data_out=16'h0;
17'h1185:	data_out=16'he8;
17'h1186:	data_out=16'hfd;
17'h1187:	data_out=16'hf6;
17'h1188:	data_out=16'hce;
17'h1189:	data_out=16'hd9;
17'h118a:	data_out=16'hfd;
17'h118b:	data_out=16'hfd;
17'h118c:	data_out=16'hfd;
17'h118d:	data_out=16'h7c;
17'h118e:	data_out=16'h3;
17'h118f:	data_out=16'h0;
17'h1190:	data_out=16'h0;
17'h1191:	data_out=16'h0;
17'h1192:	data_out=16'h0;
17'h1193:	data_out=16'h0;
17'h1194:	data_out=16'h0;
17'h1195:	data_out=16'h0;
17'h1196:	data_out=16'h0;
17'h1197:	data_out=16'h0;
17'h1198:	data_out=16'h0;
17'h1199:	data_out=16'h0;
17'h119a:	data_out=16'h0;
17'h119b:	data_out=16'h0;
17'h119c:	data_out=16'h0;
17'h119d:	data_out=16'h0;
17'h119e:	data_out=16'h0;
17'h119f:	data_out=16'h0;
17'h11a0:	data_out=16'h0;
17'h11a1:	data_out=16'hd0;
17'h11a2:	data_out=16'hfd;
17'h11a3:	data_out=16'hfd;
17'h11a4:	data_out=16'hfd;
17'h11a5:	data_out=16'hfd;
17'h11a6:	data_out=16'hb3;
17'h11a7:	data_out=16'h74;
17'h11a8:	data_out=16'h24;
17'h11a9:	data_out=16'h4;
17'h11aa:	data_out=16'h0;
17'h11ab:	data_out=16'h0;
17'h11ac:	data_out=16'h0;
17'h11ad:	data_out=16'h0;
17'h11ae:	data_out=16'h0;
17'h11af:	data_out=16'h0;
17'h11b0:	data_out=16'h0;
17'h11b1:	data_out=16'h0;
17'h11b2:	data_out=16'h0;
17'h11b3:	data_out=16'h0;
17'h11b4:	data_out=16'h0;
17'h11b5:	data_out=16'h0;
17'h11b6:	data_out=16'h0;
17'h11b7:	data_out=16'h0;
17'h11b8:	data_out=16'h0;
17'h11b9:	data_out=16'h0;
17'h11ba:	data_out=16'h0;
17'h11bb:	data_out=16'h0;
17'h11bc:	data_out=16'h0;
17'h11bd:	data_out=16'hd;
17'h11be:	data_out=16'h5d;
17'h11bf:	data_out=16'h90;
17'h11c0:	data_out=16'h79;
17'h11c1:	data_out=16'h17;
17'h11c2:	data_out=16'h6;
17'h11c3:	data_out=16'h0;
17'h11c4:	data_out=16'h0;
17'h11c5:	data_out=16'h0;
17'h11c6:	data_out=16'h0;
17'h11c7:	data_out=16'h0;
17'h11c8:	data_out=16'h0;
17'h11c9:	data_out=16'h0;
17'h11ca:	data_out=16'h0;
17'h11cb:	data_out=16'h0;
17'h11cc:	data_out=16'h0;
17'h11cd:	data_out=16'h0;
17'h11ce:	data_out=16'h0;
17'h11cf:	data_out=16'h0;
17'h11d0:	data_out=16'h0;
17'h11d1:	data_out=16'h0;
17'h11d2:	data_out=16'h0;
17'h11d3:	data_out=16'h0;
17'h11d4:	data_out=16'h0;
17'h11d5:	data_out=16'h0;
17'h11d6:	data_out=16'h0;
17'h11d7:	data_out=16'h0;
17'h11d8:	data_out=16'h0;
17'h11d9:	data_out=16'h0;
17'h11da:	data_out=16'h0;
17'h11db:	data_out=16'h0;
17'h11dc:	data_out=16'h0;
17'h11dd:	data_out=16'h0;
17'h11de:	data_out=16'h0;
17'h11df:	data_out=16'h0;
17'h11e0:	data_out=16'h0;
17'h11e1:	data_out=16'h0;
17'h11e2:	data_out=16'h0;
17'h11e3:	data_out=16'h0;
17'h11e4:	data_out=16'h0;
17'h11e5:	data_out=16'h0;
17'h11e6:	data_out=16'h0;
17'h11e7:	data_out=16'h0;
17'h11e8:	data_out=16'h0;
17'h11e9:	data_out=16'h0;
17'h11ea:	data_out=16'h0;
17'h11eb:	data_out=16'h0;
17'h11ec:	data_out=16'h0;
17'h11ed:	data_out=16'h0;
17'h11ee:	data_out=16'h0;
17'h11ef:	data_out=16'h0;
17'h11f0:	data_out=16'h0;
17'h11f1:	data_out=16'h0;
17'h11f2:	data_out=16'h0;
17'h11f3:	data_out=16'h0;
17'h11f4:	data_out=16'h0;
17'h11f5:	data_out=16'h0;
17'h11f6:	data_out=16'h0;
17'h11f7:	data_out=16'h0;
17'h11f8:	data_out=16'h0;
17'h11f9:	data_out=16'h0;
17'h11fa:	data_out=16'h0;
17'h11fb:	data_out=16'h0;
17'h11fc:	data_out=16'h0;
17'h11fd:	data_out=16'h0;
17'h11fe:	data_out=16'h0;
17'h11ff:	data_out=16'h0;
17'h1200:	data_out=16'h0;
17'h1201:	data_out=16'h0;
17'h1202:	data_out=16'h0;
17'h1203:	data_out=16'h0;
17'h1204:	data_out=16'h0;
17'h1205:	data_out=16'h0;
17'h1206:	data_out=16'h0;
17'h1207:	data_out=16'h0;
17'h1208:	data_out=16'h0;
17'h1209:	data_out=16'h0;
17'h120a:	data_out=16'h0;
17'h120b:	data_out=16'h0;
17'h120c:	data_out=16'h0;
17'h120d:	data_out=16'h0;
17'h120e:	data_out=16'h0;
17'h120f:	data_out=16'h0;
17'h1210:	data_out=16'h0;
17'h1211:	data_out=16'h0;
17'h1212:	data_out=16'h0;
17'h1213:	data_out=16'h0;
17'h1214:	data_out=16'h0;
17'h1215:	data_out=16'h0;
17'h1216:	data_out=16'h0;
17'h1217:	data_out=16'h0;
17'h1218:	data_out=16'h0;
17'h1219:	data_out=16'h0;
17'h121a:	data_out=16'h0;
17'h121b:	data_out=16'h0;
17'h121c:	data_out=16'h0;
17'h121d:	data_out=16'h0;
17'h121e:	data_out=16'h0;
17'h121f:	data_out=16'h0;
17'h1220:	data_out=16'h0;
17'h1221:	data_out=16'h0;
17'h1222:	data_out=16'h0;
17'h1223:	data_out=16'h0;
17'h1224:	data_out=16'h0;
17'h1225:	data_out=16'h0;
17'h1226:	data_out=16'h0;
17'h1227:	data_out=16'h0;
17'h1228:	data_out=16'h0;
17'h1229:	data_out=16'h0;
17'h122a:	data_out=16'h0;
17'h122b:	data_out=16'h0;
17'h122c:	data_out=16'h0;
17'h122d:	data_out=16'h0;
17'h122e:	data_out=16'h0;
17'h122f:	data_out=16'h0;
17'h1230:	data_out=16'h0;
17'h1231:	data_out=16'h0;
17'h1232:	data_out=16'h0;
17'h1233:	data_out=16'h0;
17'h1234:	data_out=16'h0;
17'h1235:	data_out=16'h0;
17'h1236:	data_out=16'h0;
17'h1237:	data_out=16'h0;
17'h1238:	data_out=16'h0;
17'h1239:	data_out=16'h0;
17'h123a:	data_out=16'h0;
17'h123b:	data_out=16'h0;
17'h123c:	data_out=16'h0;
17'h123d:	data_out=16'h0;
17'h123e:	data_out=16'h0;
17'h123f:	data_out=16'h0;
17'h1240:	data_out=16'h0;
17'h1241:	data_out=16'h0;
17'h1242:	data_out=16'h0;
17'h1243:	data_out=16'h0;
17'h1244:	data_out=16'h0;
17'h1245:	data_out=16'h0;
17'h1246:	data_out=16'h0;
17'h1247:	data_out=16'h0;
17'h1248:	data_out=16'h0;
17'h1249:	data_out=16'h0;
17'h124a:	data_out=16'h0;
17'h124b:	data_out=16'h0;
17'h124c:	data_out=16'h0;
17'h124d:	data_out=16'h0;
17'h124e:	data_out=16'h0;
17'h124f:	data_out=16'h0;
17'h1250:	data_out=16'h0;
17'h1251:	data_out=16'h0;
17'h1252:	data_out=16'h0;
17'h1253:	data_out=16'h0;
17'h1254:	data_out=16'h0;
17'h1255:	data_out=16'h0;
17'h1256:	data_out=16'h0;
17'h1257:	data_out=16'h0;
17'h1258:	data_out=16'h0;
17'h1259:	data_out=16'h0;
17'h125a:	data_out=16'h0;
17'h125b:	data_out=16'h0;
17'h125c:	data_out=16'h0;
17'h125d:	data_out=16'h0;
17'h125e:	data_out=16'h0;
17'h125f:	data_out=16'h0;
17'h1260:	data_out=16'h0;
17'h1261:	data_out=16'h0;
17'h1262:	data_out=16'h0;
17'h1263:	data_out=16'h0;
17'h1264:	data_out=16'h0;
17'h1265:	data_out=16'h0;
17'h1266:	data_out=16'h0;
17'h1267:	data_out=16'h0;
17'h1268:	data_out=16'h0;
17'h1269:	data_out=16'h0;
17'h126a:	data_out=16'h0;
17'h126b:	data_out=16'h0;
17'h126c:	data_out=16'h0;
17'h126d:	data_out=16'h0;
17'h126e:	data_out=16'h0;
17'h126f:	data_out=16'h0;
17'h1270:	data_out=16'h0;
17'h1271:	data_out=16'h0;
17'h1272:	data_out=16'h0;
17'h1273:	data_out=16'h0;
17'h1274:	data_out=16'h0;
17'h1275:	data_out=16'h0;
17'h1276:	data_out=16'h0;
17'h1277:	data_out=16'h0;
17'h1278:	data_out=16'h0;
17'h1279:	data_out=16'h0;
17'h127a:	data_out=16'h0;
17'h127b:	data_out=16'h0;
17'h127c:	data_out=16'h0;
17'h127d:	data_out=16'h0;
17'h127e:	data_out=16'h0;
17'h127f:	data_out=16'h0;
17'h1280:	data_out=16'h0;
17'h1281:	data_out=16'h0;
17'h1282:	data_out=16'h0;
17'h1283:	data_out=16'h0;
17'h1284:	data_out=16'h0;
17'h1285:	data_out=16'h0;
17'h1286:	data_out=16'h0;
17'h1287:	data_out=16'h0;
17'h1288:	data_out=16'h0;
17'h1289:	data_out=16'h0;
17'h128a:	data_out=16'h0;
17'h128b:	data_out=16'h0;
17'h128c:	data_out=16'h0;
17'h128d:	data_out=16'h0;
17'h128e:	data_out=16'h0;
17'h128f:	data_out=16'h0;
17'h1290:	data_out=16'h0;
17'h1291:	data_out=16'h0;
17'h1292:	data_out=16'h0;
17'h1293:	data_out=16'h0;
17'h1294:	data_out=16'h0;
17'h1295:	data_out=16'h0;
17'h1296:	data_out=16'h0;
17'h1297:	data_out=16'h0;
17'h1298:	data_out=16'h0;
17'h1299:	data_out=16'h0;
17'h129a:	data_out=16'h0;
17'h129b:	data_out=16'h0;
17'h129c:	data_out=16'h0;
17'h129d:	data_out=16'h0;
17'h129e:	data_out=16'h0;
17'h129f:	data_out=16'h0;
17'h12a0:	data_out=16'h0;
17'h12a1:	data_out=16'h0;
17'h12a2:	data_out=16'h0;
17'h12a3:	data_out=16'h0;
17'h12a4:	data_out=16'h0;
17'h12a5:	data_out=16'h0;
17'h12a6:	data_out=16'h0;
17'h12a7:	data_out=16'h0;
17'h12a8:	data_out=16'h0;
17'h12a9:	data_out=16'h0;
17'h12aa:	data_out=16'h0;
17'h12ab:	data_out=16'h0;
17'h12ac:	data_out=16'h0;
17'h12ad:	data_out=16'h0;
17'h12ae:	data_out=16'h0;
17'h12af:	data_out=16'h0;
17'h12b0:	data_out=16'h0;
17'h12b1:	data_out=16'h0;
17'h12b2:	data_out=16'h0;
17'h12b3:	data_out=16'h0;
17'h12b4:	data_out=16'h0;
17'h12b5:	data_out=16'h0;
17'h12b6:	data_out=16'h0;
17'h12b7:	data_out=16'h0;
17'h12b8:	data_out=16'h0;
17'h12b9:	data_out=16'h0;
17'h12ba:	data_out=16'h0;
17'h12bb:	data_out=16'h0;
17'h12bc:	data_out=16'h0;
17'h12bd:	data_out=16'h0;
17'h12be:	data_out=16'h0;
17'h12bf:	data_out=16'h0;
17'h12c0:	data_out=16'h0;
17'h12c1:	data_out=16'h0;
17'h12c2:	data_out=16'h0;
17'h12c3:	data_out=16'h0;
17'h12c4:	data_out=16'h0;
17'h12c5:	data_out=16'h0;
17'h12c6:	data_out=16'h0;
17'h12c7:	data_out=16'h0;
17'h12c8:	data_out=16'h0;
17'h12c9:	data_out=16'h0;
17'h12ca:	data_out=16'h0;
17'h12cb:	data_out=16'h0;
17'h12cc:	data_out=16'h0;
17'h12cd:	data_out=16'h0;
17'h12ce:	data_out=16'h0;
17'h12cf:	data_out=16'h0;
17'h12d0:	data_out=16'h0;
17'h12d1:	data_out=16'h0;
17'h12d2:	data_out=16'h0;
17'h12d3:	data_out=16'h0;
17'h12d4:	data_out=16'h0;
17'h12d5:	data_out=16'h0;
17'h12d6:	data_out=16'h0;
17'h12d7:	data_out=16'h0;
17'h12d8:	data_out=16'h0;
17'h12d9:	data_out=16'h0;
17'h12da:	data_out=16'h0;
17'h12db:	data_out=16'h0;
17'h12dc:	data_out=16'h92;
17'h12dd:	data_out=16'h100;
17'h12de:	data_out=16'hd4;
17'h12df:	data_out=16'h1f;
17'h12e0:	data_out=16'h0;
17'h12e1:	data_out=16'h0;
17'h12e2:	data_out=16'h0;
17'h12e3:	data_out=16'h0;
17'h12e4:	data_out=16'h0;
17'h12e5:	data_out=16'h0;
17'h12e6:	data_out=16'h0;
17'h12e7:	data_out=16'h0;
17'h12e8:	data_out=16'h0;
17'h12e9:	data_out=16'h0;
17'h12ea:	data_out=16'h0;
17'h12eb:	data_out=16'h0;
17'h12ec:	data_out=16'h0;
17'h12ed:	data_out=16'h0;
17'h12ee:	data_out=16'h0;
17'h12ef:	data_out=16'h0;
17'h12f0:	data_out=16'h0;
17'h12f1:	data_out=16'h0;
17'h12f2:	data_out=16'h0;
17'h12f3:	data_out=16'h0;
17'h12f4:	data_out=16'h0;
17'h12f5:	data_out=16'h0;
17'h12f6:	data_out=16'h0;
17'h12f7:	data_out=16'h20;
17'h12f8:	data_out=16'hee;
17'h12f9:	data_out=16'hfe;
17'h12fa:	data_out=16'hfd;
17'h12fb:	data_out=16'h47;
17'h12fc:	data_out=16'h0;
17'h12fd:	data_out=16'h0;
17'h12fe:	data_out=16'h0;
17'h12ff:	data_out=16'h0;
17'h1300:	data_out=16'h0;
17'h1301:	data_out=16'h0;
17'h1302:	data_out=16'h0;
17'h1303:	data_out=16'h0;
17'h1304:	data_out=16'h0;
17'h1305:	data_out=16'h0;
17'h1306:	data_out=16'h0;
17'h1307:	data_out=16'h0;
17'h1308:	data_out=16'h0;
17'h1309:	data_out=16'h0;
17'h130a:	data_out=16'h0;
17'h130b:	data_out=16'h0;
17'h130c:	data_out=16'h0;
17'h130d:	data_out=16'h0;
17'h130e:	data_out=16'h0;
17'h130f:	data_out=16'h0;
17'h1310:	data_out=16'h0;
17'h1311:	data_out=16'h0;
17'h1312:	data_out=16'h0;
17'h1313:	data_out=16'hb;
17'h1314:	data_out=16'hb0;
17'h1315:	data_out=16'hfe;
17'h1316:	data_out=16'hfd;
17'h1317:	data_out=16'h47;
17'h1318:	data_out=16'h0;
17'h1319:	data_out=16'h0;
17'h131a:	data_out=16'h0;
17'h131b:	data_out=16'h0;
17'h131c:	data_out=16'h0;
17'h131d:	data_out=16'h0;
17'h131e:	data_out=16'h0;
17'h131f:	data_out=16'h0;
17'h1320:	data_out=16'h0;
17'h1321:	data_out=16'h0;
17'h1322:	data_out=16'h0;
17'h1323:	data_out=16'h0;
17'h1324:	data_out=16'h0;
17'h1325:	data_out=16'h0;
17'h1326:	data_out=16'h0;
17'h1327:	data_out=16'h0;
17'h1328:	data_out=16'h0;
17'h1329:	data_out=16'h0;
17'h132a:	data_out=16'h0;
17'h132b:	data_out=16'h0;
17'h132c:	data_out=16'h0;
17'h132d:	data_out=16'h0;
17'h132e:	data_out=16'h0;
17'h132f:	data_out=16'h0;
17'h1330:	data_out=16'h91;
17'h1331:	data_out=16'hfe;
17'h1332:	data_out=16'hfd;
17'h1333:	data_out=16'h47;
17'h1334:	data_out=16'h0;
17'h1335:	data_out=16'h0;
17'h1336:	data_out=16'h0;
17'h1337:	data_out=16'h0;
17'h1338:	data_out=16'h0;
17'h1339:	data_out=16'h0;
17'h133a:	data_out=16'h0;
17'h133b:	data_out=16'h0;
17'h133c:	data_out=16'h0;
17'h133d:	data_out=16'h0;
17'h133e:	data_out=16'h0;
17'h133f:	data_out=16'h0;
17'h1340:	data_out=16'h0;
17'h1341:	data_out=16'h0;
17'h1342:	data_out=16'h0;
17'h1343:	data_out=16'h0;
17'h1344:	data_out=16'h0;
17'h1345:	data_out=16'h0;
17'h1346:	data_out=16'h0;
17'h1347:	data_out=16'h0;
17'h1348:	data_out=16'h0;
17'h1349:	data_out=16'h0;
17'h134a:	data_out=16'h0;
17'h134b:	data_out=16'h10;
17'h134c:	data_out=16'hc0;
17'h134d:	data_out=16'hfe;
17'h134e:	data_out=16'hfd;
17'h134f:	data_out=16'h47;
17'h1350:	data_out=16'h0;
17'h1351:	data_out=16'h0;
17'h1352:	data_out=16'h0;
17'h1353:	data_out=16'h0;
17'h1354:	data_out=16'h0;
17'h1355:	data_out=16'h0;
17'h1356:	data_out=16'h0;
17'h1357:	data_out=16'h0;
17'h1358:	data_out=16'h0;
17'h1359:	data_out=16'h0;
17'h135a:	data_out=16'h0;
17'h135b:	data_out=16'h0;
17'h135c:	data_out=16'h0;
17'h135d:	data_out=16'h0;
17'h135e:	data_out=16'h0;
17'h135f:	data_out=16'h0;
17'h1360:	data_out=16'h0;
17'h1361:	data_out=16'h0;
17'h1362:	data_out=16'h0;
17'h1363:	data_out=16'h0;
17'h1364:	data_out=16'h0;
17'h1365:	data_out=16'h0;
17'h1366:	data_out=16'h0;
17'h1367:	data_out=16'h1a;
17'h1368:	data_out=16'hde;
17'h1369:	data_out=16'hfe;
17'h136a:	data_out=16'hfd;
17'h136b:	data_out=16'h7c;
17'h136c:	data_out=16'h1f;
17'h136d:	data_out=16'h0;
17'h136e:	data_out=16'h0;
17'h136f:	data_out=16'h0;
17'h1370:	data_out=16'h0;
17'h1371:	data_out=16'h0;
17'h1372:	data_out=16'h0;
17'h1373:	data_out=16'h0;
17'h1374:	data_out=16'h0;
17'h1375:	data_out=16'h0;
17'h1376:	data_out=16'h0;
17'h1377:	data_out=16'h0;
17'h1378:	data_out=16'h0;
17'h1379:	data_out=16'h0;
17'h137a:	data_out=16'h0;
17'h137b:	data_out=16'h0;
17'h137c:	data_out=16'h0;
17'h137d:	data_out=16'h0;
17'h137e:	data_out=16'h0;
17'h137f:	data_out=16'h0;
17'h1380:	data_out=16'h0;
17'h1381:	data_out=16'h0;
17'h1382:	data_out=16'h0;
17'h1383:	data_out=16'h0;
17'h1384:	data_out=16'h7d;
17'h1385:	data_out=16'hfe;
17'h1386:	data_out=16'hfd;
17'h1387:	data_out=16'hfd;
17'h1388:	data_out=16'h6c;
17'h1389:	data_out=16'h0;
17'h138a:	data_out=16'h0;
17'h138b:	data_out=16'h0;
17'h138c:	data_out=16'h0;
17'h138d:	data_out=16'h0;
17'h138e:	data_out=16'h0;
17'h138f:	data_out=16'h0;
17'h1390:	data_out=16'h0;
17'h1391:	data_out=16'h0;
17'h1392:	data_out=16'h0;
17'h1393:	data_out=16'h0;
17'h1394:	data_out=16'h0;
17'h1395:	data_out=16'h0;
17'h1396:	data_out=16'h0;
17'h1397:	data_out=16'h0;
17'h1398:	data_out=16'h0;
17'h1399:	data_out=16'h0;
17'h139a:	data_out=16'h0;
17'h139b:	data_out=16'h0;
17'h139c:	data_out=16'h0;
17'h139d:	data_out=16'h0;
17'h139e:	data_out=16'h0;
17'h139f:	data_out=16'h0;
17'h13a0:	data_out=16'h0;
17'h13a1:	data_out=16'hfe;
17'h13a2:	data_out=16'hfd;
17'h13a3:	data_out=16'hfd;
17'h13a4:	data_out=16'h6c;
17'h13a5:	data_out=16'h0;
17'h13a6:	data_out=16'h0;
17'h13a7:	data_out=16'h0;
17'h13a8:	data_out=16'h0;
17'h13a9:	data_out=16'h0;
17'h13aa:	data_out=16'h0;
17'h13ab:	data_out=16'h0;
17'h13ac:	data_out=16'h0;
17'h13ad:	data_out=16'h0;
17'h13ae:	data_out=16'h0;
17'h13af:	data_out=16'h0;
17'h13b0:	data_out=16'h0;
17'h13b1:	data_out=16'h0;
17'h13b2:	data_out=16'h0;
17'h13b3:	data_out=16'h0;
17'h13b4:	data_out=16'h0;
17'h13b5:	data_out=16'h0;
17'h13b6:	data_out=16'h0;
17'h13b7:	data_out=16'h0;
17'h13b8:	data_out=16'h0;
17'h13b9:	data_out=16'h0;
17'h13ba:	data_out=16'h0;
17'h13bb:	data_out=16'h0;
17'h13bc:	data_out=16'h0;
17'h13bd:	data_out=16'h100;
17'h13be:	data_out=16'hfe;
17'h13bf:	data_out=16'hfe;
17'h13c0:	data_out=16'h6c;
17'h13c1:	data_out=16'h0;
17'h13c2:	data_out=16'h0;
17'h13c3:	data_out=16'h0;
17'h13c4:	data_out=16'h0;
17'h13c5:	data_out=16'h0;
17'h13c6:	data_out=16'h0;
17'h13c7:	data_out=16'h0;
17'h13c8:	data_out=16'h0;
17'h13c9:	data_out=16'h0;
17'h13ca:	data_out=16'h0;
17'h13cb:	data_out=16'h0;
17'h13cc:	data_out=16'h0;
17'h13cd:	data_out=16'h0;
17'h13ce:	data_out=16'h0;
17'h13cf:	data_out=16'h0;
17'h13d0:	data_out=16'h0;
17'h13d1:	data_out=16'h0;
17'h13d2:	data_out=16'h0;
17'h13d3:	data_out=16'h0;
17'h13d4:	data_out=16'h0;
17'h13d5:	data_out=16'h0;
17'h13d6:	data_out=16'h0;
17'h13d7:	data_out=16'h0;
17'h13d8:	data_out=16'h0;
17'h13d9:	data_out=16'hfe;
17'h13da:	data_out=16'hfd;
17'h13db:	data_out=16'hfd;
17'h13dc:	data_out=16'h6c;
17'h13dd:	data_out=16'h0;
17'h13de:	data_out=16'h0;
17'h13df:	data_out=16'h0;
17'h13e0:	data_out=16'h0;
17'h13e1:	data_out=16'h0;
17'h13e2:	data_out=16'h0;
17'h13e3:	data_out=16'h0;
17'h13e4:	data_out=16'h0;
17'h13e5:	data_out=16'h0;
17'h13e6:	data_out=16'h0;
17'h13e7:	data_out=16'h0;
17'h13e8:	data_out=16'h0;
17'h13e9:	data_out=16'h0;
17'h13ea:	data_out=16'h0;
17'h13eb:	data_out=16'h0;
17'h13ec:	data_out=16'h0;
17'h13ed:	data_out=16'h0;
17'h13ee:	data_out=16'h0;
17'h13ef:	data_out=16'h0;
17'h13f0:	data_out=16'h0;
17'h13f1:	data_out=16'h0;
17'h13f2:	data_out=16'h0;
17'h13f3:	data_out=16'h0;
17'h13f4:	data_out=16'h0;
17'h13f5:	data_out=16'hfe;
17'h13f6:	data_out=16'hfd;
17'h13f7:	data_out=16'hfd;
17'h13f8:	data_out=16'h6c;
17'h13f9:	data_out=16'h0;
17'h13fa:	data_out=16'h0;
17'h13fb:	data_out=16'h0;
17'h13fc:	data_out=16'h0;
17'h13fd:	data_out=16'h0;
17'h13fe:	data_out=16'h0;
17'h13ff:	data_out=16'h0;
17'h1400:	data_out=16'h0;
17'h1401:	data_out=16'h0;
17'h1402:	data_out=16'h0;
17'h1403:	data_out=16'h0;
17'h1404:	data_out=16'h0;
17'h1405:	data_out=16'h0;
17'h1406:	data_out=16'h0;
17'h1407:	data_out=16'h0;
17'h1408:	data_out=16'h0;
17'h1409:	data_out=16'h0;
17'h140a:	data_out=16'h0;
17'h140b:	data_out=16'h0;
17'h140c:	data_out=16'h0;
17'h140d:	data_out=16'h0;
17'h140e:	data_out=16'h0;
17'h140f:	data_out=16'h0;
17'h1410:	data_out=16'h0;
17'h1411:	data_out=16'hfe;
17'h1412:	data_out=16'hfd;
17'h1413:	data_out=16'hfd;
17'h1414:	data_out=16'h6c;
17'h1415:	data_out=16'h0;
17'h1416:	data_out=16'h0;
17'h1417:	data_out=16'h0;
17'h1418:	data_out=16'h0;
17'h1419:	data_out=16'h0;
17'h141a:	data_out=16'h0;
17'h141b:	data_out=16'h0;
17'h141c:	data_out=16'h0;
17'h141d:	data_out=16'h0;
17'h141e:	data_out=16'h0;
17'h141f:	data_out=16'h0;
17'h1420:	data_out=16'h0;
17'h1421:	data_out=16'h0;
17'h1422:	data_out=16'h0;
17'h1423:	data_out=16'h0;
17'h1424:	data_out=16'h0;
17'h1425:	data_out=16'h0;
17'h1426:	data_out=16'h0;
17'h1427:	data_out=16'h0;
17'h1428:	data_out=16'h0;
17'h1429:	data_out=16'h0;
17'h142a:	data_out=16'h0;
17'h142b:	data_out=16'h0;
17'h142c:	data_out=16'h0;
17'h142d:	data_out=16'h100;
17'h142e:	data_out=16'hfe;
17'h142f:	data_out=16'hfe;
17'h1430:	data_out=16'hab;
17'h1431:	data_out=16'h0;
17'h1432:	data_out=16'h0;
17'h1433:	data_out=16'h0;
17'h1434:	data_out=16'h0;
17'h1435:	data_out=16'h0;
17'h1436:	data_out=16'h0;
17'h1437:	data_out=16'h0;
17'h1438:	data_out=16'h0;
17'h1439:	data_out=16'h0;
17'h143a:	data_out=16'h0;
17'h143b:	data_out=16'h0;
17'h143c:	data_out=16'h0;
17'h143d:	data_out=16'h0;
17'h143e:	data_out=16'h0;
17'h143f:	data_out=16'h0;
17'h1440:	data_out=16'h0;
17'h1441:	data_out=16'h0;
17'h1442:	data_out=16'h0;
17'h1443:	data_out=16'h0;
17'h1444:	data_out=16'h0;
17'h1445:	data_out=16'h0;
17'h1446:	data_out=16'h0;
17'h1447:	data_out=16'h0;
17'h1448:	data_out=16'h0;
17'h1449:	data_out=16'hfe;
17'h144a:	data_out=16'hfd;
17'h144b:	data_out=16'hfd;
17'h144c:	data_out=16'hfd;
17'h144d:	data_out=16'h2a;
17'h144e:	data_out=16'h0;
17'h144f:	data_out=16'h0;
17'h1450:	data_out=16'h0;
17'h1451:	data_out=16'h0;
17'h1452:	data_out=16'h0;
17'h1453:	data_out=16'h0;
17'h1454:	data_out=16'h0;
17'h1455:	data_out=16'h0;
17'h1456:	data_out=16'h0;
17'h1457:	data_out=16'h0;
17'h1458:	data_out=16'h0;
17'h1459:	data_out=16'h0;
17'h145a:	data_out=16'h0;
17'h145b:	data_out=16'h0;
17'h145c:	data_out=16'h0;
17'h145d:	data_out=16'h0;
17'h145e:	data_out=16'h0;
17'h145f:	data_out=16'h0;
17'h1460:	data_out=16'h0;
17'h1461:	data_out=16'h0;
17'h1462:	data_out=16'h0;
17'h1463:	data_out=16'h0;
17'h1464:	data_out=16'h0;
17'h1465:	data_out=16'h96;
17'h1466:	data_out=16'hfd;
17'h1467:	data_out=16'hfd;
17'h1468:	data_out=16'hfd;
17'h1469:	data_out=16'h91;
17'h146a:	data_out=16'h0;
17'h146b:	data_out=16'h0;
17'h146c:	data_out=16'h0;
17'h146d:	data_out=16'h0;
17'h146e:	data_out=16'h0;
17'h146f:	data_out=16'h0;
17'h1470:	data_out=16'h0;
17'h1471:	data_out=16'h0;
17'h1472:	data_out=16'h0;
17'h1473:	data_out=16'h0;
17'h1474:	data_out=16'h0;
17'h1475:	data_out=16'h0;
17'h1476:	data_out=16'h0;
17'h1477:	data_out=16'h0;
17'h1478:	data_out=16'h0;
17'h1479:	data_out=16'h0;
17'h147a:	data_out=16'h0;
17'h147b:	data_out=16'h0;
17'h147c:	data_out=16'h0;
17'h147d:	data_out=16'h0;
17'h147e:	data_out=16'h0;
17'h147f:	data_out=16'h0;
17'h1480:	data_out=16'h0;
17'h1481:	data_out=16'h6d;
17'h1482:	data_out=16'hfd;
17'h1483:	data_out=16'hfd;
17'h1484:	data_out=16'hfd;
17'h1485:	data_out=16'h91;
17'h1486:	data_out=16'h0;
17'h1487:	data_out=16'h0;
17'h1488:	data_out=16'h0;
17'h1489:	data_out=16'h0;
17'h148a:	data_out=16'h0;
17'h148b:	data_out=16'h0;
17'h148c:	data_out=16'h0;
17'h148d:	data_out=16'h0;
17'h148e:	data_out=16'h0;
17'h148f:	data_out=16'h0;
17'h1490:	data_out=16'h0;
17'h1491:	data_out=16'h0;
17'h1492:	data_out=16'h0;
17'h1493:	data_out=16'h0;
17'h1494:	data_out=16'h0;
17'h1495:	data_out=16'h0;
17'h1496:	data_out=16'h0;
17'h1497:	data_out=16'h0;
17'h1498:	data_out=16'h0;
17'h1499:	data_out=16'h0;
17'h149a:	data_out=16'h0;
17'h149b:	data_out=16'h0;
17'h149c:	data_out=16'h0;
17'h149d:	data_out=16'h0;
17'h149e:	data_out=16'hdb;
17'h149f:	data_out=16'hfe;
17'h14a0:	data_out=16'hfe;
17'h14a1:	data_out=16'h100;
17'h14a2:	data_out=16'h23;
17'h14a3:	data_out=16'h0;
17'h14a4:	data_out=16'h0;
17'h14a5:	data_out=16'h0;
17'h14a6:	data_out=16'h0;
17'h14a7:	data_out=16'h0;
17'h14a8:	data_out=16'h0;
17'h14a9:	data_out=16'h0;
17'h14aa:	data_out=16'h0;
17'h14ab:	data_out=16'h0;
17'h14ac:	data_out=16'h0;
17'h14ad:	data_out=16'h0;
17'h14ae:	data_out=16'h0;
17'h14af:	data_out=16'h0;
17'h14b0:	data_out=16'h0;
17'h14b1:	data_out=16'h0;
17'h14b2:	data_out=16'h0;
17'h14b3:	data_out=16'h0;
17'h14b4:	data_out=16'h0;
17'h14b5:	data_out=16'h0;
17'h14b6:	data_out=16'h0;
17'h14b7:	data_out=16'h0;
17'h14b8:	data_out=16'h0;
17'h14b9:	data_out=16'h0;
17'h14ba:	data_out=16'hb0;
17'h14bb:	data_out=16'hfd;
17'h14bc:	data_out=16'hfd;
17'h14bd:	data_out=16'hfe;
17'h14be:	data_out=16'h23;
17'h14bf:	data_out=16'h0;
17'h14c0:	data_out=16'h0;
17'h14c1:	data_out=16'h0;
17'h14c2:	data_out=16'h0;
17'h14c3:	data_out=16'h0;
17'h14c4:	data_out=16'h0;
17'h14c5:	data_out=16'h0;
17'h14c6:	data_out=16'h0;
17'h14c7:	data_out=16'h0;
17'h14c8:	data_out=16'h0;
17'h14c9:	data_out=16'h0;
17'h14ca:	data_out=16'h0;
17'h14cb:	data_out=16'h0;
17'h14cc:	data_out=16'h0;
17'h14cd:	data_out=16'h0;
17'h14ce:	data_out=16'h0;
17'h14cf:	data_out=16'h0;
17'h14d0:	data_out=16'h0;
17'h14d1:	data_out=16'h0;
17'h14d2:	data_out=16'h0;
17'h14d3:	data_out=16'h0;
17'h14d4:	data_out=16'h0;
17'h14d5:	data_out=16'h0;
17'h14d6:	data_out=16'h49;
17'h14d7:	data_out=16'hfd;
17'h14d8:	data_out=16'hfd;
17'h14d9:	data_out=16'hfe;
17'h14da:	data_out=16'h23;
17'h14db:	data_out=16'h0;
17'h14dc:	data_out=16'h0;
17'h14dd:	data_out=16'h0;
17'h14de:	data_out=16'h0;
17'h14df:	data_out=16'h0;
17'h14e0:	data_out=16'h0;
17'h14e1:	data_out=16'h0;
17'h14e2:	data_out=16'h0;
17'h14e3:	data_out=16'h0;
17'h14e4:	data_out=16'h0;
17'h14e5:	data_out=16'h0;
17'h14e6:	data_out=16'h0;
17'h14e7:	data_out=16'h0;
17'h14e8:	data_out=16'h0;
17'h14e9:	data_out=16'h0;
17'h14ea:	data_out=16'h0;
17'h14eb:	data_out=16'h0;
17'h14ec:	data_out=16'h0;
17'h14ed:	data_out=16'h0;
17'h14ee:	data_out=16'h0;
17'h14ef:	data_out=16'h0;
17'h14f0:	data_out=16'h0;
17'h14f1:	data_out=16'h0;
17'h14f2:	data_out=16'h1f;
17'h14f3:	data_out=16'hd4;
17'h14f4:	data_out=16'hfd;
17'h14f5:	data_out=16'hfe;
17'h14f6:	data_out=16'h23;
17'h14f7:	data_out=16'h0;
17'h14f8:	data_out=16'h0;
17'h14f9:	data_out=16'h0;
17'h14fa:	data_out=16'h0;
17'h14fb:	data_out=16'h0;
17'h14fc:	data_out=16'h0;
17'h14fd:	data_out=16'h0;
17'h14fe:	data_out=16'h0;
17'h14ff:	data_out=16'h0;
17'h1500:	data_out=16'h0;
17'h1501:	data_out=16'h0;
17'h1502:	data_out=16'h0;
17'h1503:	data_out=16'h0;
17'h1504:	data_out=16'h0;
17'h1505:	data_out=16'h0;
17'h1506:	data_out=16'h0;
17'h1507:	data_out=16'h0;
17'h1508:	data_out=16'h0;
17'h1509:	data_out=16'h0;
17'h150a:	data_out=16'h0;
17'h150b:	data_out=16'h0;
17'h150c:	data_out=16'h0;
17'h150d:	data_out=16'h0;
17'h150e:	data_out=16'h0;
17'h150f:	data_out=16'h0;
17'h1510:	data_out=16'h0;
17'h1511:	data_out=16'h0;
17'h1512:	data_out=16'h0;
17'h1513:	data_out=16'h0;
17'h1514:	data_out=16'h0;
17'h1515:	data_out=16'h0;
17'h1516:	data_out=16'h0;
17'h1517:	data_out=16'h0;
17'h1518:	data_out=16'h0;
17'h1519:	data_out=16'h0;
17'h151a:	data_out=16'h0;
17'h151b:	data_out=16'h0;
17'h151c:	data_out=16'h0;
17'h151d:	data_out=16'h0;
17'h151e:	data_out=16'h0;
17'h151f:	data_out=16'h0;
17'h1520:	data_out=16'h0;
17'h1521:	data_out=16'h0;
17'h1522:	data_out=16'h0;
17'h1523:	data_out=16'h0;
17'h1524:	data_out=16'h0;
17'h1525:	data_out=16'h0;
17'h1526:	data_out=16'h0;
17'h1527:	data_out=16'h0;
17'h1528:	data_out=16'h0;
17'h1529:	data_out=16'h0;
17'h152a:	data_out=16'h0;
17'h152b:	data_out=16'h0;
17'h152c:	data_out=16'h0;
17'h152d:	data_out=16'h0;
17'h152e:	data_out=16'h0;
17'h152f:	data_out=16'h0;
17'h1530:	data_out=16'h0;
17'h1531:	data_out=16'h0;
17'h1532:	data_out=16'h0;
17'h1533:	data_out=16'h0;
17'h1534:	data_out=16'h0;
17'h1535:	data_out=16'h0;
17'h1536:	data_out=16'h0;
17'h1537:	data_out=16'h0;
17'h1538:	data_out=16'h0;
17'h1539:	data_out=16'h0;
17'h153a:	data_out=16'h0;
17'h153b:	data_out=16'h0;
17'h153c:	data_out=16'h0;
17'h153d:	data_out=16'h0;
17'h153e:	data_out=16'h0;
17'h153f:	data_out=16'h0;
17'h1540:	data_out=16'h0;
17'h1541:	data_out=16'h0;
17'h1542:	data_out=16'h0;
17'h1543:	data_out=16'h0;
17'h1544:	data_out=16'h0;
17'h1545:	data_out=16'h0;
17'h1546:	data_out=16'h0;
17'h1547:	data_out=16'h0;
17'h1548:	data_out=16'h0;
17'h1549:	data_out=16'h0;
17'h154a:	data_out=16'h0;
17'h154b:	data_out=16'h0;
17'h154c:	data_out=16'h0;
17'h154d:	data_out=16'h0;
17'h154e:	data_out=16'h0;
17'h154f:	data_out=16'h0;
17'h1550:	data_out=16'h0;
17'h1551:	data_out=16'h0;
17'h1552:	data_out=16'h0;
17'h1553:	data_out=16'h0;
17'h1554:	data_out=16'h0;
17'h1555:	data_out=16'h0;
17'h1556:	data_out=16'h0;
17'h1557:	data_out=16'h0;
17'h1558:	data_out=16'h0;
17'h1559:	data_out=16'h0;
17'h155a:	data_out=16'h0;
17'h155b:	data_out=16'h0;
17'h155c:	data_out=16'h0;
17'h155d:	data_out=16'h0;
17'h155e:	data_out=16'h0;
17'h155f:	data_out=16'h0;
17'h1560:	data_out=16'h0;
17'h1561:	data_out=16'h0;
17'h1562:	data_out=16'h0;
17'h1563:	data_out=16'h0;
17'h1564:	data_out=16'h0;
17'h1565:	data_out=16'h0;
17'h1566:	data_out=16'h0;
17'h1567:	data_out=16'h0;
17'h1568:	data_out=16'h0;
17'h1569:	data_out=16'h0;
17'h156a:	data_out=16'h0;
17'h156b:	data_out=16'h0;
17'h156c:	data_out=16'h0;
17'h156d:	data_out=16'h0;
17'h156e:	data_out=16'h0;
17'h156f:	data_out=16'h0;
17'h1570:	data_out=16'h0;
17'h1571:	data_out=16'h0;
17'h1572:	data_out=16'h0;
17'h1573:	data_out=16'h0;
17'h1574:	data_out=16'h0;
17'h1575:	data_out=16'h0;
17'h1576:	data_out=16'h0;
17'h1577:	data_out=16'h0;
17'h1578:	data_out=16'h0;
17'h1579:	data_out=16'h0;
17'h157a:	data_out=16'h0;
17'h157b:	data_out=16'h0;
17'h157c:	data_out=16'h0;
17'h157d:	data_out=16'h0;
17'h157e:	data_out=16'h0;
17'h157f:	data_out=16'h0;
17'h1580:	data_out=16'h0;
17'h1581:	data_out=16'h0;
17'h1582:	data_out=16'h0;
17'h1583:	data_out=16'h0;
17'h1584:	data_out=16'h0;
17'h1585:	data_out=16'h0;
17'h1586:	data_out=16'h0;
17'h1587:	data_out=16'h0;
17'h1588:	data_out=16'h0;
17'h1589:	data_out=16'h0;
17'h158a:	data_out=16'h0;
17'h158b:	data_out=16'h0;
17'h158c:	data_out=16'h0;
17'h158d:	data_out=16'h0;
17'h158e:	data_out=16'h0;
17'h158f:	data_out=16'h0;
17'h1590:	data_out=16'h0;
17'h1591:	data_out=16'h0;
17'h1592:	data_out=16'h0;
17'h1593:	data_out=16'h0;
17'h1594:	data_out=16'h0;
17'h1595:	data_out=16'h0;
17'h1596:	data_out=16'h0;
17'h1597:	data_out=16'h0;
17'h1598:	data_out=16'h0;
17'h1599:	data_out=16'h0;
17'h159a:	data_out=16'h0;
17'h159b:	data_out=16'h0;
17'h159c:	data_out=16'h0;
17'h159d:	data_out=16'h0;
17'h159e:	data_out=16'h0;
17'h159f:	data_out=16'h0;
17'h15a0:	data_out=16'h0;
17'h15a1:	data_out=16'h0;
17'h15a2:	data_out=16'h0;
17'h15a3:	data_out=16'h0;
17'h15a4:	data_out=16'h0;
17'h15a5:	data_out=16'h0;
17'h15a6:	data_out=16'h0;
17'h15a7:	data_out=16'h0;
17'h15a8:	data_out=16'h0;
17'h15a9:	data_out=16'h0;
17'h15aa:	data_out=16'h0;
17'h15ab:	data_out=16'h0;
17'h15ac:	data_out=16'h0;
17'h15ad:	data_out=16'h0;
17'h15ae:	data_out=16'h0;
17'h15af:	data_out=16'h0;
17'h15b0:	data_out=16'h0;
17'h15b1:	data_out=16'h0;
17'h15b2:	data_out=16'h0;
17'h15b3:	data_out=16'h0;
17'h15b4:	data_out=16'h0;
17'h15b5:	data_out=16'h0;
17'h15b6:	data_out=16'h0;
17'h15b7:	data_out=16'h0;
17'h15b8:	data_out=16'h0;
17'h15b9:	data_out=16'h0;
17'h15ba:	data_out=16'h0;
17'h15bb:	data_out=16'h0;
17'h15bc:	data_out=16'h0;
17'h15bd:	data_out=16'h0;
17'h15be:	data_out=16'h0;
17'h15bf:	data_out=16'h0;
17'h15c0:	data_out=16'h0;
17'h15c1:	data_out=16'h0;
17'h15c2:	data_out=16'h0;
17'h15c3:	data_out=16'h0;
17'h15c4:	data_out=16'h0;
17'h15c5:	data_out=16'h0;
17'h15c6:	data_out=16'h0;
17'h15c7:	data_out=16'h0;
17'h15c8:	data_out=16'h0;
17'h15c9:	data_out=16'h0;
17'h15ca:	data_out=16'h0;
17'h15cb:	data_out=16'h0;
17'h15cc:	data_out=16'h0;
17'h15cd:	data_out=16'h0;
17'h15ce:	data_out=16'h0;
17'h15cf:	data_out=16'h0;
17'h15d0:	data_out=16'h0;
17'h15d1:	data_out=16'h0;
17'h15d2:	data_out=16'h0;
17'h15d3:	data_out=16'h0;
17'h15d4:	data_out=16'h0;
17'h15d5:	data_out=16'h0;
17'h15d6:	data_out=16'h0;
17'h15d7:	data_out=16'h0;
17'h15d8:	data_out=16'h0;
17'h15d9:	data_out=16'h0;
17'h15da:	data_out=16'h0;
17'h15db:	data_out=16'h0;
17'h15dc:	data_out=16'h0;
17'h15dd:	data_out=16'h0;
17'h15de:	data_out=16'h0;
17'h15df:	data_out=16'h0;
17'h15e0:	data_out=16'h0;
17'h15e1:	data_out=16'h0;
17'h15e2:	data_out=16'h0;
17'h15e3:	data_out=16'h0;
17'h15e4:	data_out=16'h0;
17'h15e5:	data_out=16'h0;
17'h15e6:	data_out=16'h0;
17'h15e7:	data_out=16'h0;
17'h15e8:	data_out=16'h0;
17'h15e9:	data_out=16'h0;
17'h15ea:	data_out=16'h0;
17'h15eb:	data_out=16'h0;
17'h15ec:	data_out=16'h0;
17'h15ed:	data_out=16'h0;
17'h15ee:	data_out=16'h0;
17'h15ef:	data_out=16'h0;
17'h15f0:	data_out=16'h0;
17'h15f1:	data_out=16'h0;
17'h15f2:	data_out=16'h0;
17'h15f3:	data_out=16'h0;
17'h15f4:	data_out=16'h0;
17'h15f5:	data_out=16'h0;
17'h15f6:	data_out=16'h0;
17'h15f7:	data_out=16'h0;
17'h15f8:	data_out=16'h0;
17'h15f9:	data_out=16'h0;
17'h15fa:	data_out=16'h0;
17'h15fb:	data_out=16'h0;
17'h15fc:	data_out=16'h0;
17'h15fd:	data_out=16'h0;
17'h15fe:	data_out=16'h0;
17'h15ff:	data_out=16'h0;
17'h1600:	data_out=16'h0;
17'h1601:	data_out=16'h0;
17'h1602:	data_out=16'h0;
17'h1603:	data_out=16'h0;
17'h1604:	data_out=16'h0;
17'h1605:	data_out=16'h0;
17'h1606:	data_out=16'h0;
17'h1607:	data_out=16'h26;
17'h1608:	data_out=16'h2b;
17'h1609:	data_out=16'h69;
17'h160a:	data_out=16'h100;
17'h160b:	data_out=16'hfe;
17'h160c:	data_out=16'hfe;
17'h160d:	data_out=16'hfe;
17'h160e:	data_out=16'hfe;
17'h160f:	data_out=16'hfe;
17'h1610:	data_out=16'haf;
17'h1611:	data_out=16'h6;
17'h1612:	data_out=16'h0;
17'h1613:	data_out=16'h0;
17'h1614:	data_out=16'h0;
17'h1615:	data_out=16'h0;
17'h1616:	data_out=16'h0;
17'h1617:	data_out=16'h0;
17'h1618:	data_out=16'h0;
17'h1619:	data_out=16'h0;
17'h161a:	data_out=16'h0;
17'h161b:	data_out=16'h0;
17'h161c:	data_out=16'h0;
17'h161d:	data_out=16'h0;
17'h161e:	data_out=16'h0;
17'h161f:	data_out=16'h0;
17'h1620:	data_out=16'h0;
17'h1621:	data_out=16'h2b;
17'h1622:	data_out=16'h8c;
17'h1623:	data_out=16'he1;
17'h1624:	data_out=16'he3;
17'h1625:	data_out=16'hfd;
17'h1626:	data_out=16'hfe;
17'h1627:	data_out=16'hfd;
17'h1628:	data_out=16'hfd;
17'h1629:	data_out=16'hfd;
17'h162a:	data_out=16'hfd;
17'h162b:	data_out=16'hfd;
17'h162c:	data_out=16'hfd;
17'h162d:	data_out=16'h9f;
17'h162e:	data_out=16'he;
17'h162f:	data_out=16'h0;
17'h1630:	data_out=16'h0;
17'h1631:	data_out=16'h0;
17'h1632:	data_out=16'h0;
17'h1633:	data_out=16'h0;
17'h1634:	data_out=16'h0;
17'h1635:	data_out=16'h0;
17'h1636:	data_out=16'h0;
17'h1637:	data_out=16'h0;
17'h1638:	data_out=16'h0;
17'h1639:	data_out=16'h0;
17'h163a:	data_out=16'h0;
17'h163b:	data_out=16'h0;
17'h163c:	data_out=16'h0;
17'h163d:	data_out=16'hb3;
17'h163e:	data_out=16'hfd;
17'h163f:	data_out=16'hfd;
17'h1640:	data_out=16'hfd;
17'h1641:	data_out=16'hfd;
17'h1642:	data_out=16'hfe;
17'h1643:	data_out=16'hfd;
17'h1644:	data_out=16'hfd;
17'h1645:	data_out=16'hfd;
17'h1646:	data_out=16'hfd;
17'h1647:	data_out=16'hfd;
17'h1648:	data_out=16'hfd;
17'h1649:	data_out=16'hfd;
17'h164a:	data_out=16'h3b;
17'h164b:	data_out=16'h0;
17'h164c:	data_out=16'h0;
17'h164d:	data_out=16'h0;
17'h164e:	data_out=16'h0;
17'h164f:	data_out=16'h0;
17'h1650:	data_out=16'h0;
17'h1651:	data_out=16'h0;
17'h1652:	data_out=16'h0;
17'h1653:	data_out=16'h0;
17'h1654:	data_out=16'h0;
17'h1655:	data_out=16'h0;
17'h1656:	data_out=16'h0;
17'h1657:	data_out=16'h0;
17'h1658:	data_out=16'h0;
17'h1659:	data_out=16'h6d;
17'h165a:	data_out=16'hfd;
17'h165b:	data_out=16'hfd;
17'h165c:	data_out=16'he7;
17'h165d:	data_out=16'h85;
17'h165e:	data_out=16'h86;
17'h165f:	data_out=16'h85;
17'h1660:	data_out=16'h85;
17'h1661:	data_out=16'hbe;
17'h1662:	data_out=16'hfd;
17'h1663:	data_out=16'hfd;
17'h1664:	data_out=16'hfd;
17'h1665:	data_out=16'hfd;
17'h1666:	data_out=16'h3b;
17'h1667:	data_out=16'h0;
17'h1668:	data_out=16'h0;
17'h1669:	data_out=16'h0;
17'h166a:	data_out=16'h0;
17'h166b:	data_out=16'h0;
17'h166c:	data_out=16'h0;
17'h166d:	data_out=16'h0;
17'h166e:	data_out=16'h0;
17'h166f:	data_out=16'h0;
17'h1670:	data_out=16'h0;
17'h1671:	data_out=16'h0;
17'h1672:	data_out=16'h0;
17'h1673:	data_out=16'h0;
17'h1674:	data_out=16'h0;
17'h1675:	data_out=16'h4;
17'h1676:	data_out=16'h1d;
17'h1677:	data_out=16'h1d;
17'h1678:	data_out=16'h18;
17'h1679:	data_out=16'h0;
17'h167a:	data_out=16'h0;
17'h167b:	data_out=16'h0;
17'h167c:	data_out=16'h0;
17'h167d:	data_out=16'he;
17'h167e:	data_out=16'he3;
17'h167f:	data_out=16'hfd;
17'h1680:	data_out=16'hfd;
17'h1681:	data_out=16'had;
17'h1682:	data_out=16'h7;
17'h1683:	data_out=16'h0;
17'h1684:	data_out=16'h0;
17'h1685:	data_out=16'h0;
17'h1686:	data_out=16'h0;
17'h1687:	data_out=16'h0;
17'h1688:	data_out=16'h0;
17'h1689:	data_out=16'h0;
17'h168a:	data_out=16'h0;
17'h168b:	data_out=16'h0;
17'h168c:	data_out=16'h0;
17'h168d:	data_out=16'h0;
17'h168e:	data_out=16'h0;
17'h168f:	data_out=16'h0;
17'h1690:	data_out=16'h0;
17'h1691:	data_out=16'h0;
17'h1692:	data_out=16'h0;
17'h1693:	data_out=16'h0;
17'h1694:	data_out=16'h0;
17'h1695:	data_out=16'h0;
17'h1696:	data_out=16'h0;
17'h1697:	data_out=16'h0;
17'h1698:	data_out=16'h0;
17'h1699:	data_out=16'h55;
17'h169a:	data_out=16'hf4;
17'h169b:	data_out=16'hfd;
17'h169c:	data_out=16'hfd;
17'h169d:	data_out=16'h91;
17'h169e:	data_out=16'h0;
17'h169f:	data_out=16'h0;
17'h16a0:	data_out=16'h0;
17'h16a1:	data_out=16'h0;
17'h16a2:	data_out=16'h0;
17'h16a3:	data_out=16'h0;
17'h16a4:	data_out=16'h0;
17'h16a5:	data_out=16'h0;
17'h16a6:	data_out=16'h0;
17'h16a7:	data_out=16'h0;
17'h16a8:	data_out=16'h0;
17'h16a9:	data_out=16'h0;
17'h16aa:	data_out=16'h0;
17'h16ab:	data_out=16'h0;
17'h16ac:	data_out=16'h0;
17'h16ad:	data_out=16'h0;
17'h16ae:	data_out=16'h0;
17'h16af:	data_out=16'h0;
17'h16b0:	data_out=16'h0;
17'h16b1:	data_out=16'h0;
17'h16b2:	data_out=16'h0;
17'h16b3:	data_out=16'h0;
17'h16b4:	data_out=16'h58;
17'h16b5:	data_out=16'hbe;
17'h16b6:	data_out=16'hfd;
17'h16b7:	data_out=16'hfd;
17'h16b8:	data_out=16'hfd;
17'h16b9:	data_out=16'he;
17'h16ba:	data_out=16'h0;
17'h16bb:	data_out=16'h0;
17'h16bc:	data_out=16'h0;
17'h16bd:	data_out=16'h0;
17'h16be:	data_out=16'h0;
17'h16bf:	data_out=16'h0;
17'h16c0:	data_out=16'h0;
17'h16c1:	data_out=16'h0;
17'h16c2:	data_out=16'h0;
17'h16c3:	data_out=16'h0;
17'h16c4:	data_out=16'h0;
17'h16c5:	data_out=16'h0;
17'h16c6:	data_out=16'h0;
17'h16c7:	data_out=16'h0;
17'h16c8:	data_out=16'h0;
17'h16c9:	data_out=16'h0;
17'h16ca:	data_out=16'h0;
17'h16cb:	data_out=16'h0;
17'h16cc:	data_out=16'h0;
17'h16cd:	data_out=16'h0;
17'h16ce:	data_out=16'h5b;
17'h16cf:	data_out=16'hd5;
17'h16d0:	data_out=16'hf8;
17'h16d1:	data_out=16'hfd;
17'h16d2:	data_out=16'hfd;
17'h16d3:	data_out=16'hfd;
17'h16d4:	data_out=16'hcd;
17'h16d5:	data_out=16'h9;
17'h16d6:	data_out=16'h0;
17'h16d7:	data_out=16'h0;
17'h16d8:	data_out=16'h0;
17'h16d9:	data_out=16'h0;
17'h16da:	data_out=16'h0;
17'h16db:	data_out=16'h0;
17'h16dc:	data_out=16'h0;
17'h16dd:	data_out=16'h0;
17'h16de:	data_out=16'h0;
17'h16df:	data_out=16'h0;
17'h16e0:	data_out=16'h0;
17'h16e1:	data_out=16'h0;
17'h16e2:	data_out=16'h0;
17'h16e3:	data_out=16'h0;
17'h16e4:	data_out=16'h0;
17'h16e5:	data_out=16'h20;
17'h16e6:	data_out=16'h7d;
17'h16e7:	data_out=16'hc2;
17'h16e8:	data_out=16'hc2;
17'h16e9:	data_out=16'hc2;
17'h16ea:	data_out=16'hfe;
17'h16eb:	data_out=16'hfd;
17'h16ec:	data_out=16'hfd;
17'h16ed:	data_out=16'hfd;
17'h16ee:	data_out=16'hef;
17'h16ef:	data_out=16'h66;
17'h16f0:	data_out=16'h1c;
17'h16f1:	data_out=16'h0;
17'h16f2:	data_out=16'h0;
17'h16f3:	data_out=16'h0;
17'h16f4:	data_out=16'h0;
17'h16f5:	data_out=16'h0;
17'h16f6:	data_out=16'h0;
17'h16f7:	data_out=16'h0;
17'h16f8:	data_out=16'h0;
17'h16f9:	data_out=16'h0;
17'h16fa:	data_out=16'h0;
17'h16fb:	data_out=16'h0;
17'h16fc:	data_out=16'h0;
17'h16fd:	data_out=16'h0;
17'h16fe:	data_out=16'h0;
17'h16ff:	data_out=16'h0;
17'h1700:	data_out=16'h2d;
17'h1701:	data_out=16'hdf;
17'h1702:	data_out=16'hfd;
17'h1703:	data_out=16'hfd;
17'h1704:	data_out=16'hfd;
17'h1705:	data_out=16'hfd;
17'h1706:	data_out=16'hfe;
17'h1707:	data_out=16'hfd;
17'h1708:	data_out=16'hfd;
17'h1709:	data_out=16'hfd;
17'h170a:	data_out=16'hb2;
17'h170b:	data_out=16'h0;
17'h170c:	data_out=16'h0;
17'h170d:	data_out=16'h0;
17'h170e:	data_out=16'h0;
17'h170f:	data_out=16'h0;
17'h1710:	data_out=16'h0;
17'h1711:	data_out=16'h0;
17'h1712:	data_out=16'h0;
17'h1713:	data_out=16'h0;
17'h1714:	data_out=16'h0;
17'h1715:	data_out=16'h0;
17'h1716:	data_out=16'h0;
17'h1717:	data_out=16'h0;
17'h1718:	data_out=16'h0;
17'h1719:	data_out=16'h0;
17'h171a:	data_out=16'h0;
17'h171b:	data_out=16'h0;
17'h171c:	data_out=16'h2d;
17'h171d:	data_out=16'he0;
17'h171e:	data_out=16'hfe;
17'h171f:	data_out=16'hfe;
17'h1720:	data_out=16'hfe;
17'h1721:	data_out=16'hfe;
17'h1722:	data_out=16'h100;
17'h1723:	data_out=16'hfe;
17'h1724:	data_out=16'hfe;
17'h1725:	data_out=16'hfe;
17'h1726:	data_out=16'hfe;
17'h1727:	data_out=16'h4a;
17'h1728:	data_out=16'h0;
17'h1729:	data_out=16'h0;
17'h172a:	data_out=16'h0;
17'h172b:	data_out=16'h0;
17'h172c:	data_out=16'h0;
17'h172d:	data_out=16'h0;
17'h172e:	data_out=16'h0;
17'h172f:	data_out=16'h0;
17'h1730:	data_out=16'h0;
17'h1731:	data_out=16'h0;
17'h1732:	data_out=16'h0;
17'h1733:	data_out=16'h0;
17'h1734:	data_out=16'h0;
17'h1735:	data_out=16'h0;
17'h1736:	data_out=16'h0;
17'h1737:	data_out=16'h0;
17'h1738:	data_out=16'h0;
17'h1739:	data_out=16'h1f;
17'h173a:	data_out=16'h7b;
17'h173b:	data_out=16'h34;
17'h173c:	data_out=16'h2c;
17'h173d:	data_out=16'h2c;
17'h173e:	data_out=16'h2c;
17'h173f:	data_out=16'h2c;
17'h1740:	data_out=16'h90;
17'h1741:	data_out=16'hfd;
17'h1742:	data_out=16'hfd;
17'h1743:	data_out=16'h4a;
17'h1744:	data_out=16'h0;
17'h1745:	data_out=16'h0;
17'h1746:	data_out=16'h0;
17'h1747:	data_out=16'h0;
17'h1748:	data_out=16'h0;
17'h1749:	data_out=16'h0;
17'h174a:	data_out=16'h0;
17'h174b:	data_out=16'h0;
17'h174c:	data_out=16'h0;
17'h174d:	data_out=16'h0;
17'h174e:	data_out=16'h0;
17'h174f:	data_out=16'h0;
17'h1750:	data_out=16'h0;
17'h1751:	data_out=16'h0;
17'h1752:	data_out=16'h0;
17'h1753:	data_out=16'h0;
17'h1754:	data_out=16'h0;
17'h1755:	data_out=16'h0;
17'h1756:	data_out=16'h0;
17'h1757:	data_out=16'h0;
17'h1758:	data_out=16'h0;
17'h1759:	data_out=16'h0;
17'h175a:	data_out=16'h0;
17'h175b:	data_out=16'h0;
17'h175c:	data_out=16'hf;
17'h175d:	data_out=16'hfd;
17'h175e:	data_out=16'hfd;
17'h175f:	data_out=16'h4a;
17'h1760:	data_out=16'h0;
17'h1761:	data_out=16'h0;
17'h1762:	data_out=16'h0;
17'h1763:	data_out=16'h0;
17'h1764:	data_out=16'h0;
17'h1765:	data_out=16'h0;
17'h1766:	data_out=16'h0;
17'h1767:	data_out=16'h0;
17'h1768:	data_out=16'h0;
17'h1769:	data_out=16'h0;
17'h176a:	data_out=16'h0;
17'h176b:	data_out=16'h0;
17'h176c:	data_out=16'h0;
17'h176d:	data_out=16'h0;
17'h176e:	data_out=16'h0;
17'h176f:	data_out=16'h0;
17'h1770:	data_out=16'h0;
17'h1771:	data_out=16'h0;
17'h1772:	data_out=16'h0;
17'h1773:	data_out=16'h0;
17'h1774:	data_out=16'h0;
17'h1775:	data_out=16'h0;
17'h1776:	data_out=16'h0;
17'h1777:	data_out=16'h0;
17'h1778:	data_out=16'h56;
17'h1779:	data_out=16'hfd;
17'h177a:	data_out=16'hfd;
17'h177b:	data_out=16'h4a;
17'h177c:	data_out=16'h0;
17'h177d:	data_out=16'h0;
17'h177e:	data_out=16'h0;
17'h177f:	data_out=16'h0;
17'h1780:	data_out=16'h0;
17'h1781:	data_out=16'h0;
17'h1782:	data_out=16'h0;
17'h1783:	data_out=16'h0;
17'h1784:	data_out=16'h0;
17'h1785:	data_out=16'h0;
17'h1786:	data_out=16'h0;
17'h1787:	data_out=16'h0;
17'h1788:	data_out=16'h0;
17'h1789:	data_out=16'h0;
17'h178a:	data_out=16'h5;
17'h178b:	data_out=16'h4b;
17'h178c:	data_out=16'h9;
17'h178d:	data_out=16'h0;
17'h178e:	data_out=16'h0;
17'h178f:	data_out=16'h0;
17'h1790:	data_out=16'h0;
17'h1791:	data_out=16'h0;
17'h1792:	data_out=16'h0;
17'h1793:	data_out=16'h62;
17'h1794:	data_out=16'hf3;
17'h1795:	data_out=16'hfd;
17'h1796:	data_out=16'hfd;
17'h1797:	data_out=16'h4a;
17'h1798:	data_out=16'h0;
17'h1799:	data_out=16'h0;
17'h179a:	data_out=16'h0;
17'h179b:	data_out=16'h0;
17'h179c:	data_out=16'h0;
17'h179d:	data_out=16'h0;
17'h179e:	data_out=16'h0;
17'h179f:	data_out=16'h0;
17'h17a0:	data_out=16'h0;
17'h17a1:	data_out=16'h0;
17'h17a2:	data_out=16'h0;
17'h17a3:	data_out=16'h0;
17'h17a4:	data_out=16'h0;
17'h17a5:	data_out=16'h3d;
17'h17a6:	data_out=16'hb8;
17'h17a7:	data_out=16'hfd;
17'h17a8:	data_out=16'h1d;
17'h17a9:	data_out=16'h0;
17'h17aa:	data_out=16'h0;
17'h17ab:	data_out=16'h0;
17'h17ac:	data_out=16'h0;
17'h17ad:	data_out=16'h12;
17'h17ae:	data_out=16'h5c;
17'h17af:	data_out=16'hf0;
17'h17b0:	data_out=16'hfd;
17'h17b1:	data_out=16'hfd;
17'h17b2:	data_out=16'hf4;
17'h17b3:	data_out=16'h41;
17'h17b4:	data_out=16'h0;
17'h17b5:	data_out=16'h0;
17'h17b6:	data_out=16'h0;
17'h17b7:	data_out=16'h0;
17'h17b8:	data_out=16'h0;
17'h17b9:	data_out=16'h0;
17'h17ba:	data_out=16'h0;
17'h17bb:	data_out=16'h0;
17'h17bc:	data_out=16'h0;
17'h17bd:	data_out=16'h0;
17'h17be:	data_out=16'h0;
17'h17bf:	data_out=16'h0;
17'h17c0:	data_out=16'h0;
17'h17c1:	data_out=16'hd1;
17'h17c2:	data_out=16'hfd;
17'h17c3:	data_out=16'hfd;
17'h17c4:	data_out=16'h94;
17'h17c5:	data_out=16'h87;
17'h17c6:	data_out=16'h87;
17'h17c7:	data_out=16'h87;
17'h17c8:	data_out=16'h87;
17'h17c9:	data_out=16'hcc;
17'h17ca:	data_out=16'hfe;
17'h17cb:	data_out=16'hfd;
17'h17cc:	data_out=16'hfd;
17'h17cd:	data_out=16'hbd;
17'h17ce:	data_out=16'h53;
17'h17cf:	data_out=16'h0;
17'h17d0:	data_out=16'h0;
17'h17d1:	data_out=16'h0;
17'h17d2:	data_out=16'h0;
17'h17d3:	data_out=16'h0;
17'h17d4:	data_out=16'h0;
17'h17d5:	data_out=16'h0;
17'h17d6:	data_out=16'h0;
17'h17d7:	data_out=16'h0;
17'h17d8:	data_out=16'h0;
17'h17d9:	data_out=16'h0;
17'h17da:	data_out=16'h0;
17'h17db:	data_out=16'h0;
17'h17dc:	data_out=16'h0;
17'h17dd:	data_out=16'hd1;
17'h17de:	data_out=16'hfd;
17'h17df:	data_out=16'hfd;
17'h17e0:	data_out=16'hfd;
17'h17e1:	data_out=16'hfd;
17'h17e2:	data_out=16'hfd;
17'h17e3:	data_out=16'hfd;
17'h17e4:	data_out=16'hfd;
17'h17e5:	data_out=16'hfd;
17'h17e6:	data_out=16'hfe;
17'h17e7:	data_out=16'he7;
17'h17e8:	data_out=16'h9a;
17'h17e9:	data_out=16'h8;
17'h17ea:	data_out=16'h0;
17'h17eb:	data_out=16'h0;
17'h17ec:	data_out=16'h0;
17'h17ed:	data_out=16'h0;
17'h17ee:	data_out=16'h0;
17'h17ef:	data_out=16'h0;
17'h17f0:	data_out=16'h0;
17'h17f1:	data_out=16'h0;
17'h17f2:	data_out=16'h0;
17'h17f3:	data_out=16'h0;
17'h17f4:	data_out=16'h0;
17'h17f5:	data_out=16'h0;
17'h17f6:	data_out=16'h0;
17'h17f7:	data_out=16'h0;
17'h17f8:	data_out=16'h0;
17'h17f9:	data_out=16'h31;
17'h17fa:	data_out=16'h9e;
17'h17fb:	data_out=16'hfd;
17'h17fc:	data_out=16'hfd;
17'h17fd:	data_out=16'hfd;
17'h17fe:	data_out=16'hfd;
17'h17ff:	data_out=16'hfd;
17'h1800:	data_out=16'hda;
17'h1801:	data_out=16'hd0;
17'h1802:	data_out=16'h93;
17'h1803:	data_out=16'h2d;
17'h1804:	data_out=16'h0;
17'h1805:	data_out=16'h0;
17'h1806:	data_out=16'h0;
17'h1807:	data_out=16'h0;
17'h1808:	data_out=16'h0;
17'h1809:	data_out=16'h0;
17'h180a:	data_out=16'h0;
17'h180b:	data_out=16'h0;
17'h180c:	data_out=16'h0;
17'h180d:	data_out=16'h0;
17'h180e:	data_out=16'h0;
17'h180f:	data_out=16'h0;
17'h1810:	data_out=16'h0;
17'h1811:	data_out=16'h0;
17'h1812:	data_out=16'h0;
17'h1813:	data_out=16'h0;
17'h1814:	data_out=16'h0;
17'h1815:	data_out=16'h0;
17'h1816:	data_out=16'h7;
17'h1817:	data_out=16'h67;
17'h1818:	data_out=16'hec;
17'h1819:	data_out=16'hfd;
17'h181a:	data_out=16'had;
17'h181b:	data_out=16'h67;
17'h181c:	data_out=16'h18;
17'h181d:	data_out=16'h0;
17'h181e:	data_out=16'h0;
17'h181f:	data_out=16'h0;
17'h1820:	data_out=16'h0;
17'h1821:	data_out=16'h0;
17'h1822:	data_out=16'h0;
17'h1823:	data_out=16'h0;
17'h1824:	data_out=16'h0;
17'h1825:	data_out=16'h0;
17'h1826:	data_out=16'h0;
17'h1827:	data_out=16'h0;
17'h1828:	data_out=16'h0;
17'h1829:	data_out=16'h0;
17'h182a:	data_out=16'h0;
17'h182b:	data_out=16'h0;
17'h182c:	data_out=16'h0;
17'h182d:	data_out=16'h0;
17'h182e:	data_out=16'h0;
17'h182f:	data_out=16'h0;
17'h1830:	data_out=16'h0;
17'h1831:	data_out=16'h0;
17'h1832:	data_out=16'h0;
17'h1833:	data_out=16'h0;
17'h1834:	data_out=16'h0;
17'h1835:	data_out=16'h0;
17'h1836:	data_out=16'h0;
17'h1837:	data_out=16'h0;
17'h1838:	data_out=16'h0;
17'h1839:	data_out=16'h0;
17'h183a:	data_out=16'h0;
17'h183b:	data_out=16'h0;
17'h183c:	data_out=16'h0;
17'h183d:	data_out=16'h0;
17'h183e:	data_out=16'h0;
17'h183f:	data_out=16'h0;
17'h1840:	data_out=16'h0;
17'h1841:	data_out=16'h0;
17'h1842:	data_out=16'h0;
17'h1843:	data_out=16'h0;
17'h1844:	data_out=16'h0;
17'h1845:	data_out=16'h0;
17'h1846:	data_out=16'h0;
17'h1847:	data_out=16'h0;
17'h1848:	data_out=16'h0;
17'h1849:	data_out=16'h0;
17'h184a:	data_out=16'h0;
17'h184b:	data_out=16'h0;
17'h184c:	data_out=16'h0;
17'h184d:	data_out=16'h0;
17'h184e:	data_out=16'h0;
17'h184f:	data_out=16'h0;
17'h1850:	data_out=16'h0;
17'h1851:	data_out=16'h0;
17'h1852:	data_out=16'h0;
17'h1853:	data_out=16'h0;
17'h1854:	data_out=16'h0;
17'h1855:	data_out=16'h0;
17'h1856:	data_out=16'h0;
17'h1857:	data_out=16'h0;
17'h1858:	data_out=16'h0;
17'h1859:	data_out=16'h0;
17'h185a:	data_out=16'h0;
17'h185b:	data_out=16'h0;
17'h185c:	data_out=16'h0;
17'h185d:	data_out=16'h0;
17'h185e:	data_out=16'h0;
17'h185f:	data_out=16'h0;
17'h1860:	data_out=16'h0;
17'h1861:	data_out=16'h0;
17'h1862:	data_out=16'h0;
17'h1863:	data_out=16'h0;
17'h1864:	data_out=16'h0;
17'h1865:	data_out=16'h0;
17'h1866:	data_out=16'h0;
17'h1867:	data_out=16'h0;
17'h1868:	data_out=16'h0;
17'h1869:	data_out=16'h0;
17'h186a:	data_out=16'h0;
17'h186b:	data_out=16'h0;
17'h186c:	data_out=16'h0;
17'h186d:	data_out=16'h0;
17'h186e:	data_out=16'h0;
17'h186f:	data_out=16'h0;
17'h1870:	data_out=16'h0;
17'h1871:	data_out=16'h0;
17'h1872:	data_out=16'h0;
17'h1873:	data_out=16'h0;
17'h1874:	data_out=16'h0;
17'h1875:	data_out=16'h0;
17'h1876:	data_out=16'h0;
17'h1877:	data_out=16'h0;
17'h1878:	data_out=16'h0;
17'h1879:	data_out=16'h0;
17'h187a:	data_out=16'h0;
17'h187b:	data_out=16'h0;
17'h187c:	data_out=16'h0;
17'h187d:	data_out=16'h0;
17'h187e:	data_out=16'h0;
17'h187f:	data_out=16'h0;
17'h1880:	data_out=16'h0;
17'h1881:	data_out=16'h0;
17'h1882:	data_out=16'h0;
17'h1883:	data_out=16'h0;
17'h1884:	data_out=16'h0;
17'h1885:	data_out=16'h0;
17'h1886:	data_out=16'h0;
17'h1887:	data_out=16'h0;
17'h1888:	data_out=16'h0;
17'h1889:	data_out=16'h0;
17'h188a:	data_out=16'h0;
17'h188b:	data_out=16'h0;
17'h188c:	data_out=16'h0;
17'h188d:	data_out=16'h0;
17'h188e:	data_out=16'h0;
17'h188f:	data_out=16'h0;
17'h1890:	data_out=16'h0;
17'h1891:	data_out=16'h0;
17'h1892:	data_out=16'h0;
17'h1893:	data_out=16'h0;
17'h1894:	data_out=16'h0;
17'h1895:	data_out=16'h0;
17'h1896:	data_out=16'h0;
17'h1897:	data_out=16'h0;
17'h1898:	data_out=16'h0;
17'h1899:	data_out=16'h0;
17'h189a:	data_out=16'h0;
17'h189b:	data_out=16'h0;
17'h189c:	data_out=16'h0;
17'h189d:	data_out=16'h0;
17'h189e:	data_out=16'h0;
17'h189f:	data_out=16'h0;
17'h18a0:	data_out=16'h0;
17'h18a1:	data_out=16'h0;
17'h18a2:	data_out=16'h0;
17'h18a3:	data_out=16'h0;
17'h18a4:	data_out=16'h0;
17'h18a5:	data_out=16'h0;
17'h18a6:	data_out=16'h0;
17'h18a7:	data_out=16'h0;
17'h18a8:	data_out=16'h0;
17'h18a9:	data_out=16'h0;
17'h18aa:	data_out=16'h0;
17'h18ab:	data_out=16'h0;
17'h18ac:	data_out=16'h0;
17'h18ad:	data_out=16'h0;
17'h18ae:	data_out=16'h0;
17'h18af:	data_out=16'h0;
17'h18b0:	data_out=16'h0;
17'h18b1:	data_out=16'h0;
17'h18b2:	data_out=16'h0;
17'h18b3:	data_out=16'h0;
17'h18b4:	data_out=16'h0;
17'h18b5:	data_out=16'h0;
17'h18b6:	data_out=16'h0;
17'h18b7:	data_out=16'h0;
17'h18b8:	data_out=16'h0;
17'h18b9:	data_out=16'h0;
17'h18ba:	data_out=16'h0;
17'h18bb:	data_out=16'h0;
17'h18bc:	data_out=16'h0;
17'h18bd:	data_out=16'h0;
17'h18be:	data_out=16'h0;
17'h18bf:	data_out=16'h0;
17'h18c0:	data_out=16'h0;
17'h18c1:	data_out=16'h0;
17'h18c2:	data_out=16'h0;
17'h18c3:	data_out=16'h0;
17'h18c4:	data_out=16'h0;
17'h18c5:	data_out=16'h0;
17'h18c6:	data_out=16'h0;
17'h18c7:	data_out=16'h0;
17'h18c8:	data_out=16'h0;
17'h18c9:	data_out=16'h0;
17'h18ca:	data_out=16'h0;
17'h18cb:	data_out=16'h0;
17'h18cc:	data_out=16'h0;
17'h18cd:	data_out=16'h0;
17'h18ce:	data_out=16'h0;
17'h18cf:	data_out=16'h0;
17'h18d0:	data_out=16'h0;
17'h18d1:	data_out=16'h0;
17'h18d2:	data_out=16'h0;
17'h18d3:	data_out=16'h0;
17'h18d4:	data_out=16'h0;
17'h18d5:	data_out=16'h0;
17'h18d6:	data_out=16'h0;
17'h18d7:	data_out=16'h0;
17'h18d8:	data_out=16'h0;
17'h18d9:	data_out=16'h0;
17'h18da:	data_out=16'h0;
17'h18db:	data_out=16'h0;
17'h18dc:	data_out=16'h0;
17'h18dd:	data_out=16'h0;
17'h18de:	data_out=16'h0;
17'h18df:	data_out=16'h0;
17'h18e0:	data_out=16'h0;
17'h18e1:	data_out=16'h0;
17'h18e2:	data_out=16'h0;
17'h18e3:	data_out=16'h0;
17'h18e4:	data_out=16'h0;
17'h18e5:	data_out=16'h0;
17'h18e6:	data_out=16'h0;
17'h18e7:	data_out=16'h0;
17'h18e8:	data_out=16'h0;
17'h18e9:	data_out=16'h0;
17'h18ea:	data_out=16'h0;
17'h18eb:	data_out=16'h0;
17'h18ec:	data_out=16'h0;
17'h18ed:	data_out=16'h0;
17'h18ee:	data_out=16'h0;
17'h18ef:	data_out=16'h0;
17'h18f0:	data_out=16'h0;
17'h18f1:	data_out=16'h0;
17'h18f2:	data_out=16'h0;
17'h18f3:	data_out=16'h0;
17'h18f4:	data_out=16'h0;
17'h18f5:	data_out=16'h0;
17'h18f6:	data_out=16'h0;
17'h18f7:	data_out=16'h0;
17'h18f8:	data_out=16'h0;
17'h18f9:	data_out=16'h0;
17'h18fa:	data_out=16'h0;
17'h18fb:	data_out=16'h0;
17'h18fc:	data_out=16'h0;
17'h18fd:	data_out=16'h0;
17'h18fe:	data_out=16'h0;
17'h18ff:	data_out=16'h0;
17'h1900:	data_out=16'h0;
17'h1901:	data_out=16'h0;
17'h1902:	data_out=16'h0;
17'h1903:	data_out=16'h0;
17'h1904:	data_out=16'h0;
17'h1905:	data_out=16'h0;
17'h1906:	data_out=16'h0;
17'h1907:	data_out=16'h0;
17'h1908:	data_out=16'h0;
17'h1909:	data_out=16'h0;
17'h190a:	data_out=16'h0;
17'h190b:	data_out=16'h0;
17'h190c:	data_out=16'h0;
17'h190d:	data_out=16'h0;
17'h190e:	data_out=16'h0;
17'h190f:	data_out=16'h0;
17'h1910:	data_out=16'h0;
17'h1911:	data_out=16'h0;
17'h1912:	data_out=16'h0;
17'h1913:	data_out=16'h0;
17'h1914:	data_out=16'h0;
17'h1915:	data_out=16'h0;
17'h1916:	data_out=16'h0;
17'h1917:	data_out=16'h0;
17'h1918:	data_out=16'h5;
17'h1919:	data_out=16'h3f;
17'h191a:	data_out=16'hc6;
17'h191b:	data_out=16'h0;
17'h191c:	data_out=16'h0;
17'h191d:	data_out=16'h0;
17'h191e:	data_out=16'h0;
17'h191f:	data_out=16'h0;
17'h1920:	data_out=16'h0;
17'h1921:	data_out=16'h0;
17'h1922:	data_out=16'h0;
17'h1923:	data_out=16'h0;
17'h1924:	data_out=16'h0;
17'h1925:	data_out=16'h0;
17'h1926:	data_out=16'h0;
17'h1927:	data_out=16'h0;
17'h1928:	data_out=16'h0;
17'h1929:	data_out=16'h0;
17'h192a:	data_out=16'h0;
17'h192b:	data_out=16'h0;
17'h192c:	data_out=16'h0;
17'h192d:	data_out=16'h0;
17'h192e:	data_out=16'h0;
17'h192f:	data_out=16'h0;
17'h1930:	data_out=16'h0;
17'h1931:	data_out=16'h0;
17'h1932:	data_out=16'h0;
17'h1933:	data_out=16'h0;
17'h1934:	data_out=16'h14;
17'h1935:	data_out=16'hff;
17'h1936:	data_out=16'he7;
17'h1937:	data_out=16'h18;
17'h1938:	data_out=16'h0;
17'h1939:	data_out=16'h0;
17'h193a:	data_out=16'h0;
17'h193b:	data_out=16'h0;
17'h193c:	data_out=16'h0;
17'h193d:	data_out=16'h0;
17'h193e:	data_out=16'h0;
17'h193f:	data_out=16'h0;
17'h1940:	data_out=16'h0;
17'h1941:	data_out=16'h0;
17'h1942:	data_out=16'h0;
17'h1943:	data_out=16'h0;
17'h1944:	data_out=16'h0;
17'h1945:	data_out=16'h0;
17'h1946:	data_out=16'h0;
17'h1947:	data_out=16'h0;
17'h1948:	data_out=16'h0;
17'h1949:	data_out=16'h0;
17'h194a:	data_out=16'h0;
17'h194b:	data_out=16'h0;
17'h194c:	data_out=16'h0;
17'h194d:	data_out=16'h0;
17'h194e:	data_out=16'h0;
17'h194f:	data_out=16'h0;
17'h1950:	data_out=16'h14;
17'h1951:	data_out=16'hff;
17'h1952:	data_out=16'hff;
17'h1953:	data_out=16'h30;
17'h1954:	data_out=16'h0;
17'h1955:	data_out=16'h0;
17'h1956:	data_out=16'h0;
17'h1957:	data_out=16'h0;
17'h1958:	data_out=16'h0;
17'h1959:	data_out=16'h0;
17'h195a:	data_out=16'h0;
17'h195b:	data_out=16'h0;
17'h195c:	data_out=16'h0;
17'h195d:	data_out=16'h0;
17'h195e:	data_out=16'h0;
17'h195f:	data_out=16'h0;
17'h1960:	data_out=16'h0;
17'h1961:	data_out=16'h0;
17'h1962:	data_out=16'h0;
17'h1963:	data_out=16'h0;
17'h1964:	data_out=16'h0;
17'h1965:	data_out=16'h0;
17'h1966:	data_out=16'h0;
17'h1967:	data_out=16'h0;
17'h1968:	data_out=16'h0;
17'h1969:	data_out=16'h0;
17'h196a:	data_out=16'h0;
17'h196b:	data_out=16'h0;
17'h196c:	data_out=16'h14;
17'h196d:	data_out=16'hff;
17'h196e:	data_out=16'h100;
17'h196f:	data_out=16'h30;
17'h1970:	data_out=16'h0;
17'h1971:	data_out=16'h0;
17'h1972:	data_out=16'h0;
17'h1973:	data_out=16'h0;
17'h1974:	data_out=16'h0;
17'h1975:	data_out=16'h0;
17'h1976:	data_out=16'h0;
17'h1977:	data_out=16'h0;
17'h1978:	data_out=16'h0;
17'h1979:	data_out=16'h0;
17'h197a:	data_out=16'h0;
17'h197b:	data_out=16'h0;
17'h197c:	data_out=16'h0;
17'h197d:	data_out=16'h0;
17'h197e:	data_out=16'h0;
17'h197f:	data_out=16'h0;
17'h1980:	data_out=16'h0;
17'h1981:	data_out=16'h0;
17'h1982:	data_out=16'h0;
17'h1983:	data_out=16'h0;
17'h1984:	data_out=16'h0;
17'h1985:	data_out=16'h0;
17'h1986:	data_out=16'h0;
17'h1987:	data_out=16'h0;
17'h1988:	data_out=16'h14;
17'h1989:	data_out=16'hff;
17'h198a:	data_out=16'hff;
17'h198b:	data_out=16'h39;
17'h198c:	data_out=16'h0;
17'h198d:	data_out=16'h0;
17'h198e:	data_out=16'h0;
17'h198f:	data_out=16'h0;
17'h1990:	data_out=16'h0;
17'h1991:	data_out=16'h0;
17'h1992:	data_out=16'h0;
17'h1993:	data_out=16'h0;
17'h1994:	data_out=16'h0;
17'h1995:	data_out=16'h0;
17'h1996:	data_out=16'h0;
17'h1997:	data_out=16'h0;
17'h1998:	data_out=16'h0;
17'h1999:	data_out=16'h0;
17'h199a:	data_out=16'h0;
17'h199b:	data_out=16'h0;
17'h199c:	data_out=16'h0;
17'h199d:	data_out=16'h0;
17'h199e:	data_out=16'h0;
17'h199f:	data_out=16'h0;
17'h19a0:	data_out=16'h0;
17'h19a1:	data_out=16'h0;
17'h19a2:	data_out=16'h0;
17'h19a3:	data_out=16'h0;
17'h19a4:	data_out=16'h14;
17'h19a5:	data_out=16'hff;
17'h19a6:	data_out=16'hff;
17'h19a7:	data_out=16'h6c;
17'h19a8:	data_out=16'h0;
17'h19a9:	data_out=16'h0;
17'h19aa:	data_out=16'h0;
17'h19ab:	data_out=16'h0;
17'h19ac:	data_out=16'h0;
17'h19ad:	data_out=16'h0;
17'h19ae:	data_out=16'h0;
17'h19af:	data_out=16'h0;
17'h19b0:	data_out=16'h0;
17'h19b1:	data_out=16'h0;
17'h19b2:	data_out=16'h0;
17'h19b3:	data_out=16'h0;
17'h19b4:	data_out=16'h0;
17'h19b5:	data_out=16'h0;
17'h19b6:	data_out=16'h0;
17'h19b7:	data_out=16'h0;
17'h19b8:	data_out=16'h0;
17'h19b9:	data_out=16'h0;
17'h19ba:	data_out=16'h0;
17'h19bb:	data_out=16'h0;
17'h19bc:	data_out=16'h0;
17'h19bd:	data_out=16'h0;
17'h19be:	data_out=16'h0;
17'h19bf:	data_out=16'h0;
17'h19c0:	data_out=16'h10;
17'h19c1:	data_out=16'hf0;
17'h19c2:	data_out=16'hff;
17'h19c3:	data_out=16'h90;
17'h19c4:	data_out=16'h0;
17'h19c5:	data_out=16'h0;
17'h19c6:	data_out=16'h0;
17'h19c7:	data_out=16'h0;
17'h19c8:	data_out=16'h0;
17'h19c9:	data_out=16'h0;
17'h19ca:	data_out=16'h0;
17'h19cb:	data_out=16'h0;
17'h19cc:	data_out=16'h0;
17'h19cd:	data_out=16'h0;
17'h19ce:	data_out=16'h0;
17'h19cf:	data_out=16'h0;
17'h19d0:	data_out=16'h0;
17'h19d1:	data_out=16'h0;
17'h19d2:	data_out=16'h0;
17'h19d3:	data_out=16'h0;
17'h19d4:	data_out=16'h0;
17'h19d5:	data_out=16'h0;
17'h19d6:	data_out=16'h0;
17'h19d7:	data_out=16'h0;
17'h19d8:	data_out=16'h0;
17'h19d9:	data_out=16'h0;
17'h19da:	data_out=16'h0;
17'h19db:	data_out=16'h0;
17'h19dc:	data_out=16'h0;
17'h19dd:	data_out=16'hb3;
17'h19de:	data_out=16'hff;
17'h19df:	data_out=16'h90;
17'h19e0:	data_out=16'h0;
17'h19e1:	data_out=16'h0;
17'h19e2:	data_out=16'h0;
17'h19e3:	data_out=16'h0;
17'h19e4:	data_out=16'h0;
17'h19e5:	data_out=16'h0;
17'h19e6:	data_out=16'h0;
17'h19e7:	data_out=16'h0;
17'h19e8:	data_out=16'h0;
17'h19e9:	data_out=16'h0;
17'h19ea:	data_out=16'h0;
17'h19eb:	data_out=16'h0;
17'h19ec:	data_out=16'h0;
17'h19ed:	data_out=16'h0;
17'h19ee:	data_out=16'h0;
17'h19ef:	data_out=16'h0;
17'h19f0:	data_out=16'h0;
17'h19f1:	data_out=16'h0;
17'h19f2:	data_out=16'h0;
17'h19f3:	data_out=16'h0;
17'h19f4:	data_out=16'h0;
17'h19f5:	data_out=16'h0;
17'h19f6:	data_out=16'h0;
17'h19f7:	data_out=16'h0;
17'h19f8:	data_out=16'h0;
17'h19f9:	data_out=16'hb3;
17'h19fa:	data_out=16'hff;
17'h19fb:	data_out=16'h90;
17'h19fc:	data_out=16'h0;
17'h19fd:	data_out=16'h0;
17'h19fe:	data_out=16'h0;
17'h19ff:	data_out=16'h0;
17'h1a00:	data_out=16'h0;
17'h1a01:	data_out=16'h0;
17'h1a02:	data_out=16'h0;
17'h1a03:	data_out=16'h0;
17'h1a04:	data_out=16'h0;
17'h1a05:	data_out=16'h0;
17'h1a06:	data_out=16'h0;
17'h1a07:	data_out=16'h0;
17'h1a08:	data_out=16'h0;
17'h1a09:	data_out=16'h0;
17'h1a0a:	data_out=16'h0;
17'h1a0b:	data_out=16'h0;
17'h1a0c:	data_out=16'h0;
17'h1a0d:	data_out=16'h0;
17'h1a0e:	data_out=16'h0;
17'h1a0f:	data_out=16'h0;
17'h1a10:	data_out=16'h0;
17'h1a11:	data_out=16'h0;
17'h1a12:	data_out=16'h0;
17'h1a13:	data_out=16'h0;
17'h1a14:	data_out=16'h0;
17'h1a15:	data_out=16'hb3;
17'h1a16:	data_out=16'hff;
17'h1a17:	data_out=16'ha3;
17'h1a18:	data_out=16'h0;
17'h1a19:	data_out=16'h0;
17'h1a1a:	data_out=16'h0;
17'h1a1b:	data_out=16'h0;
17'h1a1c:	data_out=16'h0;
17'h1a1d:	data_out=16'h0;
17'h1a1e:	data_out=16'h0;
17'h1a1f:	data_out=16'h0;
17'h1a20:	data_out=16'h0;
17'h1a21:	data_out=16'h0;
17'h1a22:	data_out=16'h0;
17'h1a23:	data_out=16'h0;
17'h1a24:	data_out=16'h0;
17'h1a25:	data_out=16'h0;
17'h1a26:	data_out=16'h0;
17'h1a27:	data_out=16'h0;
17'h1a28:	data_out=16'h0;
17'h1a29:	data_out=16'h0;
17'h1a2a:	data_out=16'h0;
17'h1a2b:	data_out=16'h0;
17'h1a2c:	data_out=16'h0;
17'h1a2d:	data_out=16'h0;
17'h1a2e:	data_out=16'h0;
17'h1a2f:	data_out=16'h0;
17'h1a30:	data_out=16'h0;
17'h1a31:	data_out=16'hb3;
17'h1a32:	data_out=16'hff;
17'h1a33:	data_out=16'hf1;
17'h1a34:	data_out=16'h0;
17'h1a35:	data_out=16'h0;
17'h1a36:	data_out=16'h0;
17'h1a37:	data_out=16'h0;
17'h1a38:	data_out=16'h0;
17'h1a39:	data_out=16'h0;
17'h1a3a:	data_out=16'h0;
17'h1a3b:	data_out=16'h0;
17'h1a3c:	data_out=16'h0;
17'h1a3d:	data_out=16'h0;
17'h1a3e:	data_out=16'h0;
17'h1a3f:	data_out=16'h0;
17'h1a40:	data_out=16'h0;
17'h1a41:	data_out=16'h0;
17'h1a42:	data_out=16'h0;
17'h1a43:	data_out=16'h0;
17'h1a44:	data_out=16'h0;
17'h1a45:	data_out=16'h0;
17'h1a46:	data_out=16'h0;
17'h1a47:	data_out=16'h0;
17'h1a48:	data_out=16'h0;
17'h1a49:	data_out=16'h0;
17'h1a4a:	data_out=16'h0;
17'h1a4b:	data_out=16'h0;
17'h1a4c:	data_out=16'h0;
17'h1a4d:	data_out=16'h71;
17'h1a4e:	data_out=16'hff;
17'h1a4f:	data_out=16'hf1;
17'h1a50:	data_out=16'h0;
17'h1a51:	data_out=16'h0;
17'h1a52:	data_out=16'h0;
17'h1a53:	data_out=16'h0;
17'h1a54:	data_out=16'h0;
17'h1a55:	data_out=16'h0;
17'h1a56:	data_out=16'h0;
17'h1a57:	data_out=16'h0;
17'h1a58:	data_out=16'h0;
17'h1a59:	data_out=16'h0;
17'h1a5a:	data_out=16'h0;
17'h1a5b:	data_out=16'h0;
17'h1a5c:	data_out=16'h0;
17'h1a5d:	data_out=16'h0;
17'h1a5e:	data_out=16'h0;
17'h1a5f:	data_out=16'h0;
17'h1a60:	data_out=16'h0;
17'h1a61:	data_out=16'h0;
17'h1a62:	data_out=16'h0;
17'h1a63:	data_out=16'h0;
17'h1a64:	data_out=16'h0;
17'h1a65:	data_out=16'h0;
17'h1a66:	data_out=16'h0;
17'h1a67:	data_out=16'h0;
17'h1a68:	data_out=16'h0;
17'h1a69:	data_out=16'h53;
17'h1a6a:	data_out=16'hff;
17'h1a6b:	data_out=16'hf6;
17'h1a6c:	data_out=16'h1f;
17'h1a6d:	data_out=16'h0;
17'h1a6e:	data_out=16'h0;
17'h1a6f:	data_out=16'h0;
17'h1a70:	data_out=16'h0;
17'h1a71:	data_out=16'h0;
17'h1a72:	data_out=16'h0;
17'h1a73:	data_out=16'h0;
17'h1a74:	data_out=16'h0;
17'h1a75:	data_out=16'h0;
17'h1a76:	data_out=16'h0;
17'h1a77:	data_out=16'h0;
17'h1a78:	data_out=16'h0;
17'h1a79:	data_out=16'h0;
17'h1a7a:	data_out=16'h0;
17'h1a7b:	data_out=16'h0;
17'h1a7c:	data_out=16'h0;
17'h1a7d:	data_out=16'h0;
17'h1a7e:	data_out=16'h0;
17'h1a7f:	data_out=16'h0;
17'h1a80:	data_out=16'h0;
17'h1a81:	data_out=16'h0;
17'h1a82:	data_out=16'h0;
17'h1a83:	data_out=16'h0;
17'h1a84:	data_out=16'h0;
17'h1a85:	data_out=16'h4f;
17'h1a86:	data_out=16'hff;
17'h1a87:	data_out=16'hf7;
17'h1a88:	data_out=16'h26;
17'h1a89:	data_out=16'h0;
17'h1a8a:	data_out=16'h0;
17'h1a8b:	data_out=16'h0;
17'h1a8c:	data_out=16'h0;
17'h1a8d:	data_out=16'h0;
17'h1a8e:	data_out=16'h0;
17'h1a8f:	data_out=16'h0;
17'h1a90:	data_out=16'h0;
17'h1a91:	data_out=16'h0;
17'h1a92:	data_out=16'h0;
17'h1a93:	data_out=16'h0;
17'h1a94:	data_out=16'h0;
17'h1a95:	data_out=16'h0;
17'h1a96:	data_out=16'h0;
17'h1a97:	data_out=16'h0;
17'h1a98:	data_out=16'h0;
17'h1a99:	data_out=16'h0;
17'h1a9a:	data_out=16'h0;
17'h1a9b:	data_out=16'h0;
17'h1a9c:	data_out=16'h0;
17'h1a9d:	data_out=16'h0;
17'h1a9e:	data_out=16'h0;
17'h1a9f:	data_out=16'h0;
17'h1aa0:	data_out=16'h0;
17'h1aa1:	data_out=16'h0;
17'h1aa2:	data_out=16'hd7;
17'h1aa3:	data_out=16'hff;
17'h1aa4:	data_out=16'h97;
17'h1aa5:	data_out=16'h0;
17'h1aa6:	data_out=16'h0;
17'h1aa7:	data_out=16'h0;
17'h1aa8:	data_out=16'h0;
17'h1aa9:	data_out=16'h0;
17'h1aaa:	data_out=16'h0;
17'h1aab:	data_out=16'h0;
17'h1aac:	data_out=16'h0;
17'h1aad:	data_out=16'h0;
17'h1aae:	data_out=16'h0;
17'h1aaf:	data_out=16'h0;
17'h1ab0:	data_out=16'h0;
17'h1ab1:	data_out=16'h0;
17'h1ab2:	data_out=16'h0;
17'h1ab3:	data_out=16'h0;
17'h1ab4:	data_out=16'h0;
17'h1ab5:	data_out=16'h0;
17'h1ab6:	data_out=16'h0;
17'h1ab7:	data_out=16'h0;
17'h1ab8:	data_out=16'h0;
17'h1ab9:	data_out=16'h0;
17'h1aba:	data_out=16'h0;
17'h1abb:	data_out=16'h0;
17'h1abc:	data_out=16'h0;
17'h1abd:	data_out=16'h0;
17'h1abe:	data_out=16'h91;
17'h1abf:	data_out=16'hf2;
17'h1ac0:	data_out=16'h8;
17'h1ac1:	data_out=16'h0;
17'h1ac2:	data_out=16'h0;
17'h1ac3:	data_out=16'h0;
17'h1ac4:	data_out=16'h0;
17'h1ac5:	data_out=16'h0;
17'h1ac6:	data_out=16'h0;
17'h1ac7:	data_out=16'h0;
17'h1ac8:	data_out=16'h0;
17'h1ac9:	data_out=16'h0;
17'h1aca:	data_out=16'h0;
17'h1acb:	data_out=16'h0;
17'h1acc:	data_out=16'h0;
17'h1acd:	data_out=16'h0;
17'h1ace:	data_out=16'h0;
17'h1acf:	data_out=16'h0;
17'h1ad0:	data_out=16'h0;
17'h1ad1:	data_out=16'h0;
17'h1ad2:	data_out=16'h0;
17'h1ad3:	data_out=16'h0;
17'h1ad4:	data_out=16'h0;
17'h1ad5:	data_out=16'h0;
17'h1ad6:	data_out=16'h0;
17'h1ad7:	data_out=16'h0;
17'h1ad8:	data_out=16'h0;
17'h1ad9:	data_out=16'h0;
17'h1ada:	data_out=16'h91;
17'h1adb:	data_out=16'hf1;
17'h1adc:	data_out=16'h2;
17'h1add:	data_out=16'h0;
17'h1ade:	data_out=16'h0;
17'h1adf:	data_out=16'h0;
17'h1ae0:	data_out=16'h0;
17'h1ae1:	data_out=16'h0;
17'h1ae2:	data_out=16'h0;
17'h1ae3:	data_out=16'h0;
17'h1ae4:	data_out=16'h0;
17'h1ae5:	data_out=16'h0;
17'h1ae6:	data_out=16'h0;
17'h1ae7:	data_out=16'h0;
17'h1ae8:	data_out=16'h0;
17'h1ae9:	data_out=16'h0;
17'h1aea:	data_out=16'h0;
17'h1aeb:	data_out=16'h0;
17'h1aec:	data_out=16'h0;
17'h1aed:	data_out=16'h0;
17'h1aee:	data_out=16'h0;
17'h1aef:	data_out=16'h0;
17'h1af0:	data_out=16'h0;
17'h1af1:	data_out=16'h0;
17'h1af2:	data_out=16'h0;
17'h1af3:	data_out=16'h0;
17'h1af4:	data_out=16'h0;
17'h1af5:	data_out=16'h0;
17'h1af6:	data_out=16'h91;
17'h1af7:	data_out=16'hff;
17'h1af8:	data_out=16'h52;
17'h1af9:	data_out=16'h0;
17'h1afa:	data_out=16'h0;
17'h1afb:	data_out=16'h0;
17'h1afc:	data_out=16'h0;
17'h1afd:	data_out=16'h0;
17'h1afe:	data_out=16'h0;
17'h1aff:	data_out=16'h0;
17'h1b00:	data_out=16'h0;
17'h1b01:	data_out=16'h0;
17'h1b02:	data_out=16'h0;
17'h1b03:	data_out=16'h0;
17'h1b04:	data_out=16'h0;
17'h1b05:	data_out=16'h0;
17'h1b06:	data_out=16'h0;
17'h1b07:	data_out=16'h0;
17'h1b08:	data_out=16'h0;
17'h1b09:	data_out=16'h0;
17'h1b0a:	data_out=16'h0;
17'h1b0b:	data_out=16'h0;
17'h1b0c:	data_out=16'h0;
17'h1b0d:	data_out=16'h0;
17'h1b0e:	data_out=16'h0;
17'h1b0f:	data_out=16'h0;
17'h1b10:	data_out=16'h0;
17'h1b11:	data_out=16'h0;
17'h1b12:	data_out=16'he7;
17'h1b13:	data_out=16'hf8;
17'h1b14:	data_out=16'h28;
17'h1b15:	data_out=16'h0;
17'h1b16:	data_out=16'h0;
17'h1b17:	data_out=16'h0;
17'h1b18:	data_out=16'h0;
17'h1b19:	data_out=16'h0;
17'h1b1a:	data_out=16'h0;
17'h1b1b:	data_out=16'h0;
17'h1b1c:	data_out=16'h0;
17'h1b1d:	data_out=16'h0;
17'h1b1e:	data_out=16'h0;
17'h1b1f:	data_out=16'h0;
17'h1b20:	data_out=16'h0;
17'h1b21:	data_out=16'h0;
17'h1b22:	data_out=16'h0;
17'h1b23:	data_out=16'h0;
17'h1b24:	data_out=16'h0;
17'h1b25:	data_out=16'h0;
17'h1b26:	data_out=16'h0;
17'h1b27:	data_out=16'h0;
17'h1b28:	data_out=16'h0;
17'h1b29:	data_out=16'h0;
17'h1b2a:	data_out=16'h0;
17'h1b2b:	data_out=16'h0;
17'h1b2c:	data_out=16'h0;
17'h1b2d:	data_out=16'h0;
17'h1b2e:	data_out=16'ha9;
17'h1b2f:	data_out=16'hd2;
17'h1b30:	data_out=16'h1f;
17'h1b31:	data_out=16'h0;
17'h1b32:	data_out=16'h0;
17'h1b33:	data_out=16'h0;
17'h1b34:	data_out=16'h0;
17'h1b35:	data_out=16'h0;
17'h1b36:	data_out=16'h0;
17'h1b37:	data_out=16'h0;
17'h1b38:	data_out=16'h0;
17'h1b39:	data_out=16'h0;
17'h1b3a:	data_out=16'h0;
17'h1b3b:	data_out=16'h0;
17'h1b3c:	data_out=16'h0;
17'h1b3d:	data_out=16'h0;
17'h1b3e:	data_out=16'h0;
17'h1b3f:	data_out=16'h0;
17'h1b40:	data_out=16'h0;
17'h1b41:	data_out=16'h0;
17'h1b42:	data_out=16'h0;
17'h1b43:	data_out=16'h0;
17'h1b44:	data_out=16'h0;
17'h1b45:	data_out=16'h0;
17'h1b46:	data_out=16'h0;
17'h1b47:	data_out=16'h0;
17'h1b48:	data_out=16'h0;
17'h1b49:	data_out=16'h0;
17'h1b4a:	data_out=16'h0;
17'h1b4b:	data_out=16'h0;
17'h1b4c:	data_out=16'h0;
17'h1b4d:	data_out=16'h0;
17'h1b4e:	data_out=16'h0;
17'h1b4f:	data_out=16'h0;
17'h1b50:	data_out=16'h0;
17'h1b51:	data_out=16'h0;
17'h1b52:	data_out=16'h0;
17'h1b53:	data_out=16'h0;
17'h1b54:	data_out=16'h0;
17'h1b55:	data_out=16'h0;
17'h1b56:	data_out=16'h0;
17'h1b57:	data_out=16'h0;
17'h1b58:	data_out=16'h0;
17'h1b59:	data_out=16'h0;
17'h1b5a:	data_out=16'h0;
17'h1b5b:	data_out=16'h0;
17'h1b5c:	data_out=16'h0;
17'h1b5d:	data_out=16'h0;
17'h1b5e:	data_out=16'h0;
17'h1b5f:	data_out=16'h0;
17'h1b60:	data_out=16'h0;
17'h1b61:	data_out=16'h0;
17'h1b62:	data_out=16'h0;
17'h1b63:	data_out=16'h0;
17'h1b64:	data_out=16'h0;
17'h1b65:	data_out=16'h0;
17'h1b66:	data_out=16'h0;
17'h1b67:	data_out=16'h0;
17'h1b68:	data_out=16'h0;
17'h1b69:	data_out=16'h0;
17'h1b6a:	data_out=16'h0;
17'h1b6b:	data_out=16'h0;
17'h1b6c:	data_out=16'h0;
17'h1b6d:	data_out=16'h0;
17'h1b6e:	data_out=16'h0;
17'h1b6f:	data_out=16'h0;
17'h1b70:	data_out=16'h0;
17'h1b71:	data_out=16'h0;
17'h1b72:	data_out=16'h0;
17'h1b73:	data_out=16'h0;
17'h1b74:	data_out=16'h0;
17'h1b75:	data_out=16'h0;
17'h1b76:	data_out=16'h0;
17'h1b77:	data_out=16'h0;
17'h1b78:	data_out=16'h0;
17'h1b79:	data_out=16'h0;
17'h1b7a:	data_out=16'h0;
17'h1b7b:	data_out=16'h0;
17'h1b7c:	data_out=16'h0;
17'h1b7d:	data_out=16'h0;
17'h1b7e:	data_out=16'h0;
17'h1b7f:	data_out=16'h0;
17'h1b80:	data_out=16'h0;
17'h1b81:	data_out=16'h0;
17'h1b82:	data_out=16'h0;
17'h1b83:	data_out=16'h0;
17'h1b84:	data_out=16'h0;
17'h1b85:	data_out=16'h0;
17'h1b86:	data_out=16'h0;
17'h1b87:	data_out=16'h0;
17'h1b88:	data_out=16'h0;
17'h1b89:	data_out=16'h0;
17'h1b8a:	data_out=16'h0;
17'h1b8b:	data_out=16'h0;
17'h1b8c:	data_out=16'h0;
17'h1b8d:	data_out=16'h0;
17'h1b8e:	data_out=16'h0;
17'h1b8f:	data_out=16'h0;
17'h1b90:	data_out=16'h0;
17'h1b91:	data_out=16'h0;
17'h1b92:	data_out=16'h0;
17'h1b93:	data_out=16'h0;
17'h1b94:	data_out=16'h0;
17'h1b95:	data_out=16'h0;
17'h1b96:	data_out=16'h0;
17'h1b97:	data_out=16'h0;
17'h1b98:	data_out=16'h0;
17'h1b99:	data_out=16'h0;
17'h1b9a:	data_out=16'h0;
17'h1b9b:	data_out=16'h0;
17'h1b9c:	data_out=16'h0;
17'h1b9d:	data_out=16'h0;
17'h1b9e:	data_out=16'h0;
17'h1b9f:	data_out=16'h0;
17'h1ba0:	data_out=16'h0;
17'h1ba1:	data_out=16'h0;
17'h1ba2:	data_out=16'h0;
17'h1ba3:	data_out=16'h0;
17'h1ba4:	data_out=16'h0;
17'h1ba5:	data_out=16'h0;
17'h1ba6:	data_out=16'h0;
17'h1ba7:	data_out=16'h0;
17'h1ba8:	data_out=16'h0;
17'h1ba9:	data_out=16'h0;
17'h1baa:	data_out=16'h0;
17'h1bab:	data_out=16'h0;
17'h1bac:	data_out=16'h0;
17'h1bad:	data_out=16'h0;
17'h1bae:	data_out=16'h0;
17'h1baf:	data_out=16'h0;
17'h1bb0:	data_out=16'h0;
17'h1bb1:	data_out=16'h0;
17'h1bb2:	data_out=16'h0;
17'h1bb3:	data_out=16'h0;
17'h1bb4:	data_out=16'h0;
17'h1bb5:	data_out=16'h0;
17'h1bb6:	data_out=16'h0;
17'h1bb7:	data_out=16'h0;
17'h1bb8:	data_out=16'h0;
17'h1bb9:	data_out=16'h0;
17'h1bba:	data_out=16'h0;
17'h1bbb:	data_out=16'h0;
17'h1bbc:	data_out=16'h0;
17'h1bbd:	data_out=16'h0;
17'h1bbe:	data_out=16'h0;
17'h1bbf:	data_out=16'h0;
17'h1bc0:	data_out=16'h0;
17'h1bc1:	data_out=16'h0;
17'h1bc2:	data_out=16'h0;
17'h1bc3:	data_out=16'h0;
17'h1bc4:	data_out=16'h0;
17'h1bc5:	data_out=16'h0;
17'h1bc6:	data_out=16'h0;
17'h1bc7:	data_out=16'h0;
17'h1bc8:	data_out=16'h0;
17'h1bc9:	data_out=16'h0;
17'h1bca:	data_out=16'h0;
17'h1bcb:	data_out=16'h0;
17'h1bcc:	data_out=16'h0;
17'h1bcd:	data_out=16'h0;
17'h1bce:	data_out=16'h0;
17'h1bcf:	data_out=16'h0;
17'h1bd0:	data_out=16'h0;
17'h1bd1:	data_out=16'h0;
17'h1bd2:	data_out=16'h0;
17'h1bd3:	data_out=16'h0;
17'h1bd4:	data_out=16'h0;
17'h1bd5:	data_out=16'h0;
17'h1bd6:	data_out=16'h0;
17'h1bd7:	data_out=16'h0;
17'h1bd8:	data_out=16'h0;
17'h1bd9:	data_out=16'h0;
17'h1bda:	data_out=16'h0;
17'h1bdb:	data_out=16'h0;
17'h1bdc:	data_out=16'h0;
17'h1bdd:	data_out=16'h0;
17'h1bde:	data_out=16'h0;
17'h1bdf:	data_out=16'h0;
17'h1be0:	data_out=16'h0;
17'h1be1:	data_out=16'h0;
17'h1be2:	data_out=16'h0;
17'h1be3:	data_out=16'h0;
17'h1be4:	data_out=16'h0;
17'h1be5:	data_out=16'h0;
17'h1be6:	data_out=16'h0;
17'h1be7:	data_out=16'h0;
17'h1be8:	data_out=16'h0;
17'h1be9:	data_out=16'h0;
17'h1bea:	data_out=16'h0;
17'h1beb:	data_out=16'h0;
17'h1bec:	data_out=16'h0;
17'h1bed:	data_out=16'h0;
17'h1bee:	data_out=16'h0;
17'h1bef:	data_out=16'h0;
17'h1bf0:	data_out=16'h0;
17'h1bf1:	data_out=16'h0;
17'h1bf2:	data_out=16'h0;
17'h1bf3:	data_out=16'h0;
17'h1bf4:	data_out=16'h0;
17'h1bf5:	data_out=16'h0;
17'h1bf6:	data_out=16'h0;
17'h1bf7:	data_out=16'h0;
17'h1bf8:	data_out=16'h0;
17'h1bf9:	data_out=16'h0;
17'h1bfa:	data_out=16'h0;
17'h1bfb:	data_out=16'h0;
17'h1bfc:	data_out=16'h0;
17'h1bfd:	data_out=16'h0;
17'h1bfe:	data_out=16'h0;
17'h1bff:	data_out=16'h0;
17'h1c00:	data_out=16'h0;
17'h1c01:	data_out=16'h0;
17'h1c02:	data_out=16'h0;
17'h1c03:	data_out=16'h0;
17'h1c04:	data_out=16'h0;
17'h1c05:	data_out=16'h0;
17'h1c06:	data_out=16'h0;
17'h1c07:	data_out=16'h0;
17'h1c08:	data_out=16'h0;
17'h1c09:	data_out=16'h0;
17'h1c0a:	data_out=16'h0;
17'h1c0b:	data_out=16'h0;
17'h1c0c:	data_out=16'h0;
17'h1c0d:	data_out=16'h0;
17'h1c0e:	data_out=16'h0;
17'h1c0f:	data_out=16'h0;
17'h1c10:	data_out=16'h0;
17'h1c11:	data_out=16'h0;
17'h1c12:	data_out=16'h0;
17'h1c13:	data_out=16'h0;
17'h1c14:	data_out=16'h0;
17'h1c15:	data_out=16'h0;
17'h1c16:	data_out=16'hbe;
17'h1c17:	data_out=16'hbf;
17'h1c18:	data_out=16'h0;
17'h1c19:	data_out=16'h0;
17'h1c1a:	data_out=16'h0;
17'h1c1b:	data_out=16'h0;
17'h1c1c:	data_out=16'h0;
17'h1c1d:	data_out=16'h0;
17'h1c1e:	data_out=16'h0;
17'h1c1f:	data_out=16'h0;
17'h1c20:	data_out=16'h0;
17'h1c21:	data_out=16'h0;
17'h1c22:	data_out=16'h0;
17'h1c23:	data_out=16'h0;
17'h1c24:	data_out=16'h0;
17'h1c25:	data_out=16'h0;
17'h1c26:	data_out=16'h0;
17'h1c27:	data_out=16'h0;
17'h1c28:	data_out=16'h0;
17'h1c29:	data_out=16'h0;
17'h1c2a:	data_out=16'h0;
17'h1c2b:	data_out=16'h0;
17'h1c2c:	data_out=16'h0;
17'h1c2d:	data_out=16'h0;
17'h1c2e:	data_out=16'h0;
17'h1c2f:	data_out=16'h0;
17'h1c30:	data_out=16'h0;
17'h1c31:	data_out=16'h90;
17'h1c32:	data_out=16'hf8;
17'h1c33:	data_out=16'h9a;
17'h1c34:	data_out=16'h0;
17'h1c35:	data_out=16'h0;
17'h1c36:	data_out=16'h0;
17'h1c37:	data_out=16'h0;
17'h1c38:	data_out=16'h0;
17'h1c39:	data_out=16'h0;
17'h1c3a:	data_out=16'h0;
17'h1c3b:	data_out=16'h0;
17'h1c3c:	data_out=16'h0;
17'h1c3d:	data_out=16'h0;
17'h1c3e:	data_out=16'h0;
17'h1c3f:	data_out=16'h0;
17'h1c40:	data_out=16'h0;
17'h1c41:	data_out=16'h0;
17'h1c42:	data_out=16'h0;
17'h1c43:	data_out=16'h0;
17'h1c44:	data_out=16'h0;
17'h1c45:	data_out=16'h0;
17'h1c46:	data_out=16'h0;
17'h1c47:	data_out=16'h0;
17'h1c48:	data_out=16'h0;
17'h1c49:	data_out=16'h0;
17'h1c4a:	data_out=16'h0;
17'h1c4b:	data_out=16'h0;
17'h1c4c:	data_out=16'h89;
17'h1c4d:	data_out=16'hf8;
17'h1c4e:	data_out=16'hf3;
17'h1c4f:	data_out=16'h56;
17'h1c50:	data_out=16'h0;
17'h1c51:	data_out=16'h0;
17'h1c52:	data_out=16'h0;
17'h1c53:	data_out=16'h0;
17'h1c54:	data_out=16'h0;
17'h1c55:	data_out=16'h0;
17'h1c56:	data_out=16'h0;
17'h1c57:	data_out=16'h0;
17'h1c58:	data_out=16'h0;
17'h1c59:	data_out=16'h0;
17'h1c5a:	data_out=16'h0;
17'h1c5b:	data_out=16'h0;
17'h1c5c:	data_out=16'h0;
17'h1c5d:	data_out=16'h0;
17'h1c5e:	data_out=16'h0;
17'h1c5f:	data_out=16'h0;
17'h1c60:	data_out=16'h0;
17'h1c61:	data_out=16'h0;
17'h1c62:	data_out=16'h0;
17'h1c63:	data_out=16'h0;
17'h1c64:	data_out=16'h0;
17'h1c65:	data_out=16'h0;
17'h1c66:	data_out=16'h0;
17'h1c67:	data_out=16'h0;
17'h1c68:	data_out=16'hc1;
17'h1c69:	data_out=16'hfd;
17'h1c6a:	data_out=16'hbc;
17'h1c6b:	data_out=16'h0;
17'h1c6c:	data_out=16'h0;
17'h1c6d:	data_out=16'h0;
17'h1c6e:	data_out=16'h0;
17'h1c6f:	data_out=16'h0;
17'h1c70:	data_out=16'h0;
17'h1c71:	data_out=16'h0;
17'h1c72:	data_out=16'h0;
17'h1c73:	data_out=16'h0;
17'h1c74:	data_out=16'h0;
17'h1c75:	data_out=16'h0;
17'h1c76:	data_out=16'h0;
17'h1c77:	data_out=16'h0;
17'h1c78:	data_out=16'h0;
17'h1c79:	data_out=16'h0;
17'h1c7a:	data_out=16'h0;
17'h1c7b:	data_out=16'h0;
17'h1c7c:	data_out=16'h3e;
17'h1c7d:	data_out=16'hba;
17'h1c7e:	data_out=16'h12;
17'h1c7f:	data_out=16'h0;
17'h1c80:	data_out=16'h0;
17'h1c81:	data_out=16'h0;
17'h1c82:	data_out=16'h0;
17'h1c83:	data_out=16'h59;
17'h1c84:	data_out=16'hed;
17'h1c85:	data_out=16'hda;
17'h1c86:	data_out=16'h2f;
17'h1c87:	data_out=16'h0;
17'h1c88:	data_out=16'h0;
17'h1c89:	data_out=16'h0;
17'h1c8a:	data_out=16'h0;
17'h1c8b:	data_out=16'h0;
17'h1c8c:	data_out=16'h0;
17'h1c8d:	data_out=16'h0;
17'h1c8e:	data_out=16'h0;
17'h1c8f:	data_out=16'h0;
17'h1c90:	data_out=16'h0;
17'h1c91:	data_out=16'h0;
17'h1c92:	data_out=16'h0;
17'h1c93:	data_out=16'h0;
17'h1c94:	data_out=16'h0;
17'h1c95:	data_out=16'h0;
17'h1c96:	data_out=16'h0;
17'h1c97:	data_out=16'h0;
17'h1c98:	data_out=16'hd9;
17'h1c99:	data_out=16'hfe;
17'h1c9a:	data_out=16'h3c;
17'h1c9b:	data_out=16'h0;
17'h1c9c:	data_out=16'h0;
17'h1c9d:	data_out=16'h0;
17'h1c9e:	data_out=16'h0;
17'h1c9f:	data_out=16'hd5;
17'h1ca0:	data_out=16'h100;
17'h1ca1:	data_out=16'h51;
17'h1ca2:	data_out=16'h0;
17'h1ca3:	data_out=16'h0;
17'h1ca4:	data_out=16'h0;
17'h1ca5:	data_out=16'h0;
17'h1ca6:	data_out=16'h0;
17'h1ca7:	data_out=16'h0;
17'h1ca8:	data_out=16'h0;
17'h1ca9:	data_out=16'h0;
17'h1caa:	data_out=16'h0;
17'h1cab:	data_out=16'h0;
17'h1cac:	data_out=16'h0;
17'h1cad:	data_out=16'h0;
17'h1cae:	data_out=16'h0;
17'h1caf:	data_out=16'h0;
17'h1cb0:	data_out=16'h0;
17'h1cb1:	data_out=16'h0;
17'h1cb2:	data_out=16'h0;
17'h1cb3:	data_out=16'h0;
17'h1cb4:	data_out=16'hcf;
17'h1cb5:	data_out=16'hfd;
17'h1cb6:	data_out=16'h44;
17'h1cb7:	data_out=16'h0;
17'h1cb8:	data_out=16'h0;
17'h1cb9:	data_out=16'h0;
17'h1cba:	data_out=16'h30;
17'h1cbb:	data_out=16'hf3;
17'h1cbc:	data_out=16'hfe;
17'h1cbd:	data_out=16'h59;
17'h1cbe:	data_out=16'h0;
17'h1cbf:	data_out=16'h0;
17'h1cc0:	data_out=16'h0;
17'h1cc1:	data_out=16'h0;
17'h1cc2:	data_out=16'h0;
17'h1cc3:	data_out=16'h0;
17'h1cc4:	data_out=16'h0;
17'h1cc5:	data_out=16'h0;
17'h1cc6:	data_out=16'h0;
17'h1cc7:	data_out=16'h0;
17'h1cc8:	data_out=16'h0;
17'h1cc9:	data_out=16'h0;
17'h1cca:	data_out=16'h0;
17'h1ccb:	data_out=16'h0;
17'h1ccc:	data_out=16'h0;
17'h1ccd:	data_out=16'h0;
17'h1cce:	data_out=16'h0;
17'h1ccf:	data_out=16'h84;
17'h1cd0:	data_out=16'hfc;
17'h1cd1:	data_out=16'hd5;
17'h1cd2:	data_out=16'h15;
17'h1cd3:	data_out=16'h0;
17'h1cd4:	data_out=16'h0;
17'h1cd5:	data_out=16'hb;
17'h1cd6:	data_out=16'ha8;
17'h1cd7:	data_out=16'hfd;
17'h1cd8:	data_out=16'hc6;
17'h1cd9:	data_out=16'h5;
17'h1cda:	data_out=16'h0;
17'h1cdb:	data_out=16'h0;
17'h1cdc:	data_out=16'h0;
17'h1cdd:	data_out=16'h0;
17'h1cde:	data_out=16'h0;
17'h1cdf:	data_out=16'h0;
17'h1ce0:	data_out=16'h0;
17'h1ce1:	data_out=16'h0;
17'h1ce2:	data_out=16'h0;
17'h1ce3:	data_out=16'h0;
17'h1ce4:	data_out=16'h0;
17'h1ce5:	data_out=16'h0;
17'h1ce6:	data_out=16'h0;
17'h1ce7:	data_out=16'h0;
17'h1ce8:	data_out=16'h0;
17'h1ce9:	data_out=16'h0;
17'h1cea:	data_out=16'h1d;
17'h1ceb:	data_out=16'he9;
17'h1cec:	data_out=16'hf8;
17'h1ced:	data_out=16'h3f;
17'h1cee:	data_out=16'h0;
17'h1cef:	data_out=16'h0;
17'h1cf0:	data_out=16'h0;
17'h1cf1:	data_out=16'h9a;
17'h1cf2:	data_out=16'hfd;
17'h1cf3:	data_out=16'he3;
17'h1cf4:	data_out=16'h0;
17'h1cf5:	data_out=16'h0;
17'h1cf6:	data_out=16'h0;
17'h1cf7:	data_out=16'h0;
17'h1cf8:	data_out=16'h0;
17'h1cf9:	data_out=16'h0;
17'h1cfa:	data_out=16'h0;
17'h1cfb:	data_out=16'h0;
17'h1cfc:	data_out=16'h0;
17'h1cfd:	data_out=16'h0;
17'h1cfe:	data_out=16'h0;
17'h1cff:	data_out=16'h0;
17'h1d00:	data_out=16'h0;
17'h1d01:	data_out=16'h0;
17'h1d02:	data_out=16'h0;
17'h1d03:	data_out=16'h0;
17'h1d04:	data_out=16'h0;
17'h1d05:	data_out=16'h2d;
17'h1d06:	data_out=16'hdc;
17'h1d07:	data_out=16'hfd;
17'h1d08:	data_out=16'h90;
17'h1d09:	data_out=16'h0;
17'h1d0a:	data_out=16'h0;
17'h1d0b:	data_out=16'h0;
17'h1d0c:	data_out=16'h74;
17'h1d0d:	data_out=16'hfa;
17'h1d0e:	data_out=16'hfd;
17'h1d0f:	data_out=16'h67;
17'h1d10:	data_out=16'h0;
17'h1d11:	data_out=16'h0;
17'h1d12:	data_out=16'h0;
17'h1d13:	data_out=16'h0;
17'h1d14:	data_out=16'h0;
17'h1d15:	data_out=16'h0;
17'h1d16:	data_out=16'h0;
17'h1d17:	data_out=16'h0;
17'h1d18:	data_out=16'h0;
17'h1d19:	data_out=16'h0;
17'h1d1a:	data_out=16'h0;
17'h1d1b:	data_out=16'h0;
17'h1d1c:	data_out=16'h0;
17'h1d1d:	data_out=16'h0;
17'h1d1e:	data_out=16'h0;
17'h1d1f:	data_out=16'h4;
17'h1d20:	data_out=16'h60;
17'h1d21:	data_out=16'hfe;
17'h1d22:	data_out=16'h100;
17'h1d23:	data_out=16'hfe;
17'h1d24:	data_out=16'hc9;
17'h1d25:	data_out=16'h7a;
17'h1d26:	data_out=16'h7;
17'h1d27:	data_out=16'h19;
17'h1d28:	data_out=16'hca;
17'h1d29:	data_out=16'hfb;
17'h1d2a:	data_out=16'h9f;
17'h1d2b:	data_out=16'h0;
17'h1d2c:	data_out=16'h0;
17'h1d2d:	data_out=16'h0;
17'h1d2e:	data_out=16'h0;
17'h1d2f:	data_out=16'h0;
17'h1d30:	data_out=16'h0;
17'h1d31:	data_out=16'h0;
17'h1d32:	data_out=16'h0;
17'h1d33:	data_out=16'h0;
17'h1d34:	data_out=16'h0;
17'h1d35:	data_out=16'h0;
17'h1d36:	data_out=16'h0;
17'h1d37:	data_out=16'h0;
17'h1d38:	data_out=16'h0;
17'h1d39:	data_out=16'h0;
17'h1d3a:	data_out=16'h0;
17'h1d3b:	data_out=16'h5c;
17'h1d3c:	data_out=16'hfd;
17'h1d3d:	data_out=16'hfd;
17'h1d3e:	data_out=16'hfe;
17'h1d3f:	data_out=16'hda;
17'h1d40:	data_out=16'hfd;
17'h1d41:	data_out=16'hfd;
17'h1d42:	data_out=16'hc9;
17'h1d43:	data_out=16'he4;
17'h1d44:	data_out=16'hfd;
17'h1d45:	data_out=16'he8;
17'h1d46:	data_out=16'h0;
17'h1d47:	data_out=16'h0;
17'h1d48:	data_out=16'h0;
17'h1d49:	data_out=16'h0;
17'h1d4a:	data_out=16'h0;
17'h1d4b:	data_out=16'h0;
17'h1d4c:	data_out=16'h0;
17'h1d4d:	data_out=16'h0;
17'h1d4e:	data_out=16'h0;
17'h1d4f:	data_out=16'h0;
17'h1d50:	data_out=16'h0;
17'h1d51:	data_out=16'h0;
17'h1d52:	data_out=16'h0;
17'h1d53:	data_out=16'h0;
17'h1d54:	data_out=16'h0;
17'h1d55:	data_out=16'h0;
17'h1d56:	data_out=16'h57;
17'h1d57:	data_out=16'hfc;
17'h1d58:	data_out=16'hf8;
17'h1d59:	data_out=16'he8;
17'h1d5a:	data_out=16'h41;
17'h1d5b:	data_out=16'h30;
17'h1d5c:	data_out=16'hbe;
17'h1d5d:	data_out=16'hfd;
17'h1d5e:	data_out=16'hfd;
17'h1d5f:	data_out=16'hfe;
17'h1d60:	data_out=16'hfd;
17'h1d61:	data_out=16'hfc;
17'h1d62:	data_out=16'he4;
17'h1d63:	data_out=16'h23;
17'h1d64:	data_out=16'h0;
17'h1d65:	data_out=16'h0;
17'h1d66:	data_out=16'h0;
17'h1d67:	data_out=16'h0;
17'h1d68:	data_out=16'h0;
17'h1d69:	data_out=16'h0;
17'h1d6a:	data_out=16'h0;
17'h1d6b:	data_out=16'h0;
17'h1d6c:	data_out=16'h0;
17'h1d6d:	data_out=16'h0;
17'h1d6e:	data_out=16'h0;
17'h1d6f:	data_out=16'h0;
17'h1d70:	data_out=16'h0;
17'h1d71:	data_out=16'h0;
17'h1d72:	data_out=16'hbf;
17'h1d73:	data_out=16'hde;
17'h1d74:	data_out=16'h62;
17'h1d75:	data_out=16'h0;
17'h1d76:	data_out=16'h0;
17'h1d77:	data_out=16'h0;
17'h1d78:	data_out=16'h2a;
17'h1d79:	data_out=16'hc5;
17'h1d7a:	data_out=16'hfd;
17'h1d7b:	data_out=16'hfe;
17'h1d7c:	data_out=16'hfd;
17'h1d7d:	data_out=16'hfd;
17'h1d7e:	data_out=16'ha3;
17'h1d7f:	data_out=16'h0;
17'h1d80:	data_out=16'h0;
17'h1d81:	data_out=16'h0;
17'h1d82:	data_out=16'h0;
17'h1d83:	data_out=16'h0;
17'h1d84:	data_out=16'h0;
17'h1d85:	data_out=16'h0;
17'h1d86:	data_out=16'h0;
17'h1d87:	data_out=16'h0;
17'h1d88:	data_out=16'h0;
17'h1d89:	data_out=16'h0;
17'h1d8a:	data_out=16'h0;
17'h1d8b:	data_out=16'h0;
17'h1d8c:	data_out=16'h0;
17'h1d8d:	data_out=16'h0;
17'h1d8e:	data_out=16'h6f;
17'h1d8f:	data_out=16'h1d;
17'h1d90:	data_out=16'h0;
17'h1d91:	data_out=16'h0;
17'h1d92:	data_out=16'h0;
17'h1d93:	data_out=16'h0;
17'h1d94:	data_out=16'h3e;
17'h1d95:	data_out=16'hf0;
17'h1d96:	data_out=16'hfd;
17'h1d97:	data_out=16'h56;
17'h1d98:	data_out=16'h2a;
17'h1d99:	data_out=16'h2a;
17'h1d9a:	data_out=16'he;
17'h1d9b:	data_out=16'h0;
17'h1d9c:	data_out=16'h0;
17'h1d9d:	data_out=16'h0;
17'h1d9e:	data_out=16'h0;
17'h1d9f:	data_out=16'h0;
17'h1da0:	data_out=16'h0;
17'h1da1:	data_out=16'h0;
17'h1da2:	data_out=16'h0;
17'h1da3:	data_out=16'h0;
17'h1da4:	data_out=16'h0;
17'h1da5:	data_out=16'h0;
17'h1da6:	data_out=16'h0;
17'h1da7:	data_out=16'h0;
17'h1da8:	data_out=16'h0;
17'h1da9:	data_out=16'h0;
17'h1daa:	data_out=16'h0;
17'h1dab:	data_out=16'h0;
17'h1dac:	data_out=16'h0;
17'h1dad:	data_out=16'h0;
17'h1dae:	data_out=16'h0;
17'h1daf:	data_out=16'hf;
17'h1db0:	data_out=16'h95;
17'h1db1:	data_out=16'hfe;
17'h1db2:	data_out=16'hdb;
17'h1db3:	data_out=16'h0;
17'h1db4:	data_out=16'h0;
17'h1db5:	data_out=16'h0;
17'h1db6:	data_out=16'h0;
17'h1db7:	data_out=16'h0;
17'h1db8:	data_out=16'h0;
17'h1db9:	data_out=16'h0;
17'h1dba:	data_out=16'h0;
17'h1dbb:	data_out=16'h0;
17'h1dbc:	data_out=16'h0;
17'h1dbd:	data_out=16'h0;
17'h1dbe:	data_out=16'h0;
17'h1dbf:	data_out=16'h0;
17'h1dc0:	data_out=16'h0;
17'h1dc1:	data_out=16'h0;
17'h1dc2:	data_out=16'h0;
17'h1dc3:	data_out=16'h0;
17'h1dc4:	data_out=16'h0;
17'h1dc5:	data_out=16'h0;
17'h1dc6:	data_out=16'h0;
17'h1dc7:	data_out=16'h0;
17'h1dc8:	data_out=16'h0;
17'h1dc9:	data_out=16'h0;
17'h1dca:	data_out=16'h0;
17'h1dcb:	data_out=16'h79;
17'h1dcc:	data_out=16'hfd;
17'h1dcd:	data_out=16'he8;
17'h1dce:	data_out=16'h1c;
17'h1dcf:	data_out=16'h0;
17'h1dd0:	data_out=16'h0;
17'h1dd1:	data_out=16'h0;
17'h1dd2:	data_out=16'h0;
17'h1dd3:	data_out=16'h0;
17'h1dd4:	data_out=16'h0;
17'h1dd5:	data_out=16'h0;
17'h1dd6:	data_out=16'h0;
17'h1dd7:	data_out=16'h0;
17'h1dd8:	data_out=16'h0;
17'h1dd9:	data_out=16'h0;
17'h1dda:	data_out=16'h0;
17'h1ddb:	data_out=16'h0;
17'h1ddc:	data_out=16'h0;
17'h1ddd:	data_out=16'h0;
17'h1dde:	data_out=16'h0;
17'h1ddf:	data_out=16'h0;
17'h1de0:	data_out=16'h0;
17'h1de1:	data_out=16'h0;
17'h1de2:	data_out=16'h0;
17'h1de3:	data_out=16'h0;
17'h1de4:	data_out=16'h0;
17'h1de5:	data_out=16'h0;
17'h1de6:	data_out=16'h1f;
17'h1de7:	data_out=16'hde;
17'h1de8:	data_out=16'hfc;
17'h1de9:	data_out=16'h82;
17'h1dea:	data_out=16'h0;
17'h1deb:	data_out=16'h0;
17'h1dec:	data_out=16'h0;
17'h1ded:	data_out=16'h0;
17'h1dee:	data_out=16'h0;
17'h1def:	data_out=16'h0;
17'h1df0:	data_out=16'h0;
17'h1df1:	data_out=16'h0;
17'h1df2:	data_out=16'h0;
17'h1df3:	data_out=16'h0;
17'h1df4:	data_out=16'h0;
17'h1df5:	data_out=16'h0;
17'h1df6:	data_out=16'h0;
17'h1df7:	data_out=16'h0;
17'h1df8:	data_out=16'h0;
17'h1df9:	data_out=16'h0;
17'h1dfa:	data_out=16'h0;
17'h1dfb:	data_out=16'h0;
17'h1dfc:	data_out=16'h0;
17'h1dfd:	data_out=16'h0;
17'h1dfe:	data_out=16'h0;
17'h1dff:	data_out=16'h0;
17'h1e00:	data_out=16'h0;
17'h1e01:	data_out=16'h0;
17'h1e02:	data_out=16'hdb;
17'h1e03:	data_out=16'hfd;
17'h1e04:	data_out=16'ha1;
17'h1e05:	data_out=16'h0;
17'h1e06:	data_out=16'h0;
17'h1e07:	data_out=16'h0;
17'h1e08:	data_out=16'h0;
17'h1e09:	data_out=16'h0;
17'h1e0a:	data_out=16'h0;
17'h1e0b:	data_out=16'h0;
17'h1e0c:	data_out=16'h0;
17'h1e0d:	data_out=16'h0;
17'h1e0e:	data_out=16'h0;
17'h1e0f:	data_out=16'h0;
17'h1e10:	data_out=16'h0;
17'h1e11:	data_out=16'h0;
17'h1e12:	data_out=16'h0;
17'h1e13:	data_out=16'h0;
17'h1e14:	data_out=16'h0;
17'h1e15:	data_out=16'h0;
17'h1e16:	data_out=16'h0;
17'h1e17:	data_out=16'h0;
17'h1e18:	data_out=16'h0;
17'h1e19:	data_out=16'h0;
17'h1e1a:	data_out=16'h0;
17'h1e1b:	data_out=16'h0;
17'h1e1c:	data_out=16'h0;
17'h1e1d:	data_out=16'h0;
17'h1e1e:	data_out=16'h7a;
17'h1e1f:	data_out=16'hfd;
17'h1e20:	data_out=16'h52;
17'h1e21:	data_out=16'h0;
17'h1e22:	data_out=16'h0;
17'h1e23:	data_out=16'h0;
17'h1e24:	data_out=16'h0;
17'h1e25:	data_out=16'h0;
17'h1e26:	data_out=16'h0;
17'h1e27:	data_out=16'h0;
17'h1e28:	data_out=16'h0;
17'h1e29:	data_out=16'h0;
17'h1e2a:	data_out=16'h0;
17'h1e2b:	data_out=16'h0;
17'h1e2c:	data_out=16'h0;
17'h1e2d:	data_out=16'h0;
17'h1e2e:	data_out=16'h0;
17'h1e2f:	data_out=16'h0;
17'h1e30:	data_out=16'h0;
17'h1e31:	data_out=16'h0;
17'h1e32:	data_out=16'h0;
17'h1e33:	data_out=16'h0;
17'h1e34:	data_out=16'h0;
17'h1e35:	data_out=16'h0;
17'h1e36:	data_out=16'h0;
17'h1e37:	data_out=16'h0;
17'h1e38:	data_out=16'h0;
17'h1e39:	data_out=16'h0;
17'h1e3a:	data_out=16'h0;
17'h1e3b:	data_out=16'h0;
17'h1e3c:	data_out=16'h0;
17'h1e3d:	data_out=16'h0;
17'h1e3e:	data_out=16'h0;
17'h1e3f:	data_out=16'h0;
17'h1e40:	data_out=16'h0;
17'h1e41:	data_out=16'h0;
17'h1e42:	data_out=16'h0;
17'h1e43:	data_out=16'h0;
17'h1e44:	data_out=16'h0;
17'h1e45:	data_out=16'h0;
17'h1e46:	data_out=16'h0;
17'h1e47:	data_out=16'h0;
17'h1e48:	data_out=16'h0;
17'h1e49:	data_out=16'h0;
17'h1e4a:	data_out=16'h0;
17'h1e4b:	data_out=16'h0;
17'h1e4c:	data_out=16'h0;
17'h1e4d:	data_out=16'h0;
17'h1e4e:	data_out=16'h0;
17'h1e4f:	data_out=16'h0;
17'h1e50:	data_out=16'h0;
17'h1e51:	data_out=16'h0;
17'h1e52:	data_out=16'h0;
17'h1e53:	data_out=16'h0;
17'h1e54:	data_out=16'h0;
17'h1e55:	data_out=16'h0;
17'h1e56:	data_out=16'h0;
17'h1e57:	data_out=16'h0;
17'h1e58:	data_out=16'h0;
17'h1e59:	data_out=16'h0;
17'h1e5a:	data_out=16'h0;
17'h1e5b:	data_out=16'h0;
17'h1e5c:	data_out=16'h0;
17'h1e5d:	data_out=16'h0;
17'h1e5e:	data_out=16'h0;
17'h1e5f:	data_out=16'h0;
17'h1e60:	data_out=16'h0;
17'h1e61:	data_out=16'h0;
17'h1e62:	data_out=16'h0;
17'h1e63:	data_out=16'h0;
17'h1e64:	data_out=16'h0;
17'h1e65:	data_out=16'h0;
17'h1e66:	data_out=16'h0;
17'h1e67:	data_out=16'h0;
17'h1e68:	data_out=16'h0;
17'h1e69:	data_out=16'h0;
17'h1e6a:	data_out=16'h0;
17'h1e6b:	data_out=16'h0;
17'h1e6c:	data_out=16'h0;
17'h1e6d:	data_out=16'h0;
17'h1e6e:	data_out=16'h0;
17'h1e6f:	data_out=16'h0;
17'h1e70:	data_out=16'h0;
17'h1e71:	data_out=16'h0;
17'h1e72:	data_out=16'h0;
17'h1e73:	data_out=16'h0;
17'h1e74:	data_out=16'h0;
17'h1e75:	data_out=16'h0;
17'h1e76:	data_out=16'h0;
17'h1e77:	data_out=16'h0;
17'h1e78:	data_out=16'h0;
17'h1e79:	data_out=16'h0;
17'h1e7a:	data_out=16'h0;
17'h1e7b:	data_out=16'h0;
17'h1e7c:	data_out=16'h0;
17'h1e7d:	data_out=16'h0;
17'h1e7e:	data_out=16'h0;
17'h1e7f:	data_out=16'h0;
17'h1e80:	data_out=16'h0;
17'h1e81:	data_out=16'h0;
17'h1e82:	data_out=16'h0;
17'h1e83:	data_out=16'h0;
17'h1e84:	data_out=16'h0;
17'h1e85:	data_out=16'h0;
17'h1e86:	data_out=16'h0;
17'h1e87:	data_out=16'h0;
17'h1e88:	data_out=16'h0;
17'h1e89:	data_out=16'h0;
17'h1e8a:	data_out=16'h0;
17'h1e8b:	data_out=16'h0;
17'h1e8c:	data_out=16'h0;
17'h1e8d:	data_out=16'h0;
17'h1e8e:	data_out=16'h0;
17'h1e8f:	data_out=16'h0;
17'h1e90:	data_out=16'h0;
17'h1e91:	data_out=16'h0;
17'h1e92:	data_out=16'h0;
17'h1e93:	data_out=16'h0;
17'h1e94:	data_out=16'h0;
17'h1e95:	data_out=16'h0;
17'h1e96:	data_out=16'h0;
17'h1e97:	data_out=16'h0;
17'h1e98:	data_out=16'h0;
17'h1e99:	data_out=16'h0;
17'h1e9a:	data_out=16'h0;
17'h1e9b:	data_out=16'h0;
17'h1e9c:	data_out=16'h0;
17'h1e9d:	data_out=16'h0;
17'h1e9e:	data_out=16'h0;
		default: #7 data_out=32'hFFFF;
	endcase
end
endmodule

module ReadOnlyMemory_WIH(output reg [15:0] data_out, input [16:0] address);
always@(address)begin
	case(address) 
    17'h0:	data_out=16'h0;
17'h1:	data_out=16'h2;
17'h2:	data_out=16'h8006;
17'h3:	data_out=16'h8008;
17'h4:	data_out=16'h9;
17'h5:	data_out=16'h0;
17'h6:	data_out=16'h8004;
17'h7:	data_out=16'h8009;
17'h8:	data_out=16'h5;
17'h9:	data_out=16'h8004;
17'ha:	data_out=16'h8003;
17'hb:	data_out=16'h2;
17'hc:	data_out=16'h4;
17'hd:	data_out=16'h8;
17'he:	data_out=16'h8009;
17'hf:	data_out=16'h8009;
17'h10:	data_out=16'h3;
17'h11:	data_out=16'h8002;
17'h12:	data_out=16'h2;
17'h13:	data_out=16'h8004;
17'h14:	data_out=16'h8008;
17'h15:	data_out=16'h8003;
17'h16:	data_out=16'h5;
17'h17:	data_out=16'h0;
17'h18:	data_out=16'h8007;
17'h19:	data_out=16'h4;
17'h1a:	data_out=16'h8;
17'h1b:	data_out=16'h8001;
17'h1c:	data_out=16'h8004;
17'h1d:	data_out=16'h8004;
17'h1e:	data_out=16'h8003;
17'h1f:	data_out=16'h6;
17'h20:	data_out=16'h7;
17'h21:	data_out=16'h8000;
17'h22:	data_out=16'h7;
17'h23:	data_out=16'h7;
17'h24:	data_out=16'h8009;
17'h25:	data_out=16'h8006;
17'h26:	data_out=16'h7;
17'h27:	data_out=16'h5;
17'h28:	data_out=16'h8002;
17'h29:	data_out=16'h8005;
17'h2a:	data_out=16'h8002;
17'h2b:	data_out=16'h8007;
17'h2c:	data_out=16'h8007;
17'h2d:	data_out=16'h8002;
17'h2e:	data_out=16'h8007;
17'h2f:	data_out=16'h5;
17'h30:	data_out=16'h5;
17'h31:	data_out=16'h5;
17'h32:	data_out=16'h8008;
17'h33:	data_out=16'h7;
17'h34:	data_out=16'h8008;
17'h35:	data_out=16'h6;
17'h36:	data_out=16'h8002;
17'h37:	data_out=16'h8006;
17'h38:	data_out=16'h1;
17'h39:	data_out=16'h8003;
17'h3a:	data_out=16'h3;
17'h3b:	data_out=16'h7;
17'h3c:	data_out=16'h2;
17'h3d:	data_out=16'h9;
17'h3e:	data_out=16'h3;
17'h3f:	data_out=16'h8001;
17'h40:	data_out=16'h8001;
17'h41:	data_out=16'h1;
17'h42:	data_out=16'h8003;
17'h43:	data_out=16'h8000;
17'h44:	data_out=16'h4;
17'h45:	data_out=16'h8005;
17'h46:	data_out=16'h8005;
17'h47:	data_out=16'h8007;
17'h48:	data_out=16'h8001;
17'h49:	data_out=16'h2;
17'h4a:	data_out=16'h8005;
17'h4b:	data_out=16'h1;
17'h4c:	data_out=16'h9;
17'h4d:	data_out=16'h8003;
17'h4e:	data_out=16'h8003;
17'h4f:	data_out=16'h5;
17'h50:	data_out=16'h8007;
17'h51:	data_out=16'h8002;
17'h52:	data_out=16'h3;
17'h53:	data_out=16'h8006;
17'h54:	data_out=16'h8004;
17'h55:	data_out=16'h8009;
17'h56:	data_out=16'h8002;
17'h57:	data_out=16'h6;
17'h58:	data_out=16'h8003;
17'h59:	data_out=16'h8009;
17'h5a:	data_out=16'h4;
17'h5b:	data_out=16'h8;
17'h5c:	data_out=16'h8009;
17'h5d:	data_out=16'h8002;
17'h5e:	data_out=16'h8001;
17'h5f:	data_out=16'h8000;
17'h60:	data_out=16'h8;
17'h61:	data_out=16'h5;
17'h62:	data_out=16'h8;
17'h63:	data_out=16'h3;
17'h64:	data_out=16'h9;
17'h65:	data_out=16'h8006;
17'h66:	data_out=16'h5;
17'h67:	data_out=16'h8002;
17'h68:	data_out=16'h5;
17'h69:	data_out=16'h9;
17'h6a:	data_out=16'h8;
17'h6b:	data_out=16'h4;
17'h6c:	data_out=16'h8003;
17'h6d:	data_out=16'h8004;
17'h6e:	data_out=16'h0;
17'h6f:	data_out=16'h8001;
17'h70:	data_out=16'h4;
17'h71:	data_out=16'h8006;
17'h72:	data_out=16'h2;
17'h73:	data_out=16'h9;
17'h74:	data_out=16'h8006;
17'h75:	data_out=16'h8009;
17'h76:	data_out=16'h6;
17'h77:	data_out=16'h1;
17'h78:	data_out=16'h8008;
17'h79:	data_out=16'h1;
17'h7a:	data_out=16'h8000;
17'h7b:	data_out=16'h8008;
17'h7c:	data_out=16'h8;
17'h7d:	data_out=16'h7;
17'h7e:	data_out=16'h1;
17'h7f:	data_out=16'h7;
17'h80:	data_out=16'h3;
17'h81:	data_out=16'h8000;
17'h82:	data_out=16'h1;
17'h83:	data_out=16'h2;
17'h84:	data_out=16'h3;
17'h85:	data_out=16'h8004;
17'h86:	data_out=16'h8009;
17'h87:	data_out=16'h8001;
17'h88:	data_out=16'h8004;
17'h89:	data_out=16'h9;
17'h8a:	data_out=16'h8006;
17'h8b:	data_out=16'h2;
17'h8c:	data_out=16'h8004;
17'h8d:	data_out=16'h3;
17'h8e:	data_out=16'h8008;
17'h8f:	data_out=16'h8;
17'h90:	data_out=16'h6;
17'h91:	data_out=16'h4;
17'h92:	data_out=16'h8;
17'h93:	data_out=16'h8008;
17'h94:	data_out=16'h4;
17'h95:	data_out=16'h5;
17'h96:	data_out=16'h1;
17'h97:	data_out=16'h5;
17'h98:	data_out=16'h8004;
17'h99:	data_out=16'h8008;
17'h9a:	data_out=16'h6;
17'h9b:	data_out=16'h8005;
17'h9c:	data_out=16'h9;
17'h9d:	data_out=16'h8003;
17'h9e:	data_out=16'h8007;
17'h9f:	data_out=16'h2;
17'ha0:	data_out=16'h6;
17'ha1:	data_out=16'h3;
17'ha2:	data_out=16'h8004;
17'ha3:	data_out=16'h8000;
17'ha4:	data_out=16'h8;
17'ha5:	data_out=16'h8004;
17'ha6:	data_out=16'h8;
17'ha7:	data_out=16'h8005;
17'ha8:	data_out=16'h8005;
17'ha9:	data_out=16'h8007;
17'haa:	data_out=16'h7;
17'hab:	data_out=16'h0;
17'hac:	data_out=16'h6;
17'had:	data_out=16'h8;
17'hae:	data_out=16'h8001;
17'haf:	data_out=16'h3;
17'hb0:	data_out=16'h3;
17'hb1:	data_out=16'h8002;
17'hb2:	data_out=16'h4;
17'hb3:	data_out=16'h8002;
17'hb4:	data_out=16'h8007;
17'hb5:	data_out=16'h8004;
17'hb6:	data_out=16'h8007;
17'hb7:	data_out=16'h8001;
17'hb8:	data_out=16'h8003;
17'hb9:	data_out=16'h8;
17'hba:	data_out=16'h3;
17'hbb:	data_out=16'h8004;
17'hbc:	data_out=16'h8004;
17'hbd:	data_out=16'h5;
17'hbe:	data_out=16'h8;
17'hbf:	data_out=16'h8007;
17'hc0:	data_out=16'h8001;
17'hc1:	data_out=16'h8006;
17'hc2:	data_out=16'h2;
17'hc3:	data_out=16'h8002;
17'hc4:	data_out=16'h8001;
17'hc5:	data_out=16'h1;
17'hc6:	data_out=16'h3;
17'hc7:	data_out=16'h4;
17'hc8:	data_out=16'h3;
17'hc9:	data_out=16'h8000;
17'hca:	data_out=16'h8005;
17'hcb:	data_out=16'h8001;
17'hcc:	data_out=16'h8001;
17'hcd:	data_out=16'h3;
17'hce:	data_out=16'h8007;
17'hcf:	data_out=16'h8008;
17'hd0:	data_out=16'h8008;
17'hd1:	data_out=16'h5;
17'hd2:	data_out=16'h8001;
17'hd3:	data_out=16'h8006;
17'hd4:	data_out=16'h8008;
17'hd5:	data_out=16'h1;
17'hd6:	data_out=16'h2;
17'hd7:	data_out=16'h8002;
17'hd8:	data_out=16'h0;
17'hd9:	data_out=16'h8004;
17'hda:	data_out=16'h4;
17'hdb:	data_out=16'h5;
17'hdc:	data_out=16'h8008;
17'hdd:	data_out=16'h3;
17'hde:	data_out=16'h7;
17'hdf:	data_out=16'h0;
17'he0:	data_out=16'h6;
17'he1:	data_out=16'h8001;
17'he2:	data_out=16'h8;
17'he3:	data_out=16'h8004;
17'he4:	data_out=16'h8009;
17'he5:	data_out=16'h1;
17'he6:	data_out=16'h8009;
17'he7:	data_out=16'h3;
17'he8:	data_out=16'h8008;
17'he9:	data_out=16'h8005;
17'hea:	data_out=16'h8008;
17'heb:	data_out=16'h8000;
17'hec:	data_out=16'h7;
17'hed:	data_out=16'h8006;
17'hee:	data_out=16'h1;
17'hef:	data_out=16'h8;
17'hf0:	data_out=16'h9;
17'hf1:	data_out=16'h8009;
17'hf2:	data_out=16'h8007;
17'hf3:	data_out=16'h8008;
17'hf4:	data_out=16'h2;
17'hf5:	data_out=16'h5;
17'hf6:	data_out=16'h8001;
17'hf7:	data_out=16'h8007;
17'hf8:	data_out=16'h8008;
17'hf9:	data_out=16'h8006;
17'hfa:	data_out=16'h7;
17'hfb:	data_out=16'h8007;
17'hfc:	data_out=16'h6;
17'hfd:	data_out=16'h4;
17'hfe:	data_out=16'h3;
17'hff:	data_out=16'h2;
17'h100:	data_out=16'h8005;
17'h101:	data_out=16'h1;
17'h102:	data_out=16'h8;
17'h103:	data_out=16'h8005;
17'h104:	data_out=16'h8007;
17'h105:	data_out=16'h8;
17'h106:	data_out=16'h7;
17'h107:	data_out=16'h8006;
17'h108:	data_out=16'h8006;
17'h109:	data_out=16'h8;
17'h10a:	data_out=16'h3;
17'h10b:	data_out=16'h8009;
17'h10c:	data_out=16'h8007;
17'h10d:	data_out=16'h8004;
17'h10e:	data_out=16'h9;
17'h10f:	data_out=16'h8007;
17'h110:	data_out=16'h8004;
17'h111:	data_out=16'h8007;
17'h112:	data_out=16'h8007;
17'h113:	data_out=16'h7;
17'h114:	data_out=16'h6;
17'h115:	data_out=16'h2;
17'h116:	data_out=16'h9;
17'h117:	data_out=16'h7;
17'h118:	data_out=16'h5;
17'h119:	data_out=16'h6;
17'h11a:	data_out=16'h8009;
17'h11b:	data_out=16'h1;
17'h11c:	data_out=16'h1;
17'h11d:	data_out=16'h3;
17'h11e:	data_out=16'h8006;
17'h11f:	data_out=16'h5;
17'h120:	data_out=16'h8005;
17'h121:	data_out=16'h8007;
17'h122:	data_out=16'h8009;
17'h123:	data_out=16'h8003;
17'h124:	data_out=16'h8008;
17'h125:	data_out=16'h7;
17'h126:	data_out=16'h0;
17'h127:	data_out=16'h8005;
17'h128:	data_out=16'h6;
17'h129:	data_out=16'h8005;
17'h12a:	data_out=16'h8005;
17'h12b:	data_out=16'h8;
17'h12c:	data_out=16'h8001;
17'h12d:	data_out=16'h8006;
17'h12e:	data_out=16'h8009;
17'h12f:	data_out=16'h5;
17'h130:	data_out=16'h8004;
17'h131:	data_out=16'h8006;
17'h132:	data_out=16'h2;
17'h133:	data_out=16'h8006;
17'h134:	data_out=16'h5;
17'h135:	data_out=16'h2;
17'h136:	data_out=16'h8008;
17'h137:	data_out=16'h0;
17'h138:	data_out=16'h8001;
17'h139:	data_out=16'h8008;
17'h13a:	data_out=16'h8008;
17'h13b:	data_out=16'h8009;
17'h13c:	data_out=16'h4;
17'h13d:	data_out=16'h8004;
17'h13e:	data_out=16'h6;
17'h13f:	data_out=16'h7;
17'h140:	data_out=16'h8002;
17'h141:	data_out=16'h6;
17'h142:	data_out=16'h8005;
17'h143:	data_out=16'h8001;
17'h144:	data_out=16'h4;
17'h145:	data_out=16'h5;
17'h146:	data_out=16'h3;
17'h147:	data_out=16'h0;
17'h148:	data_out=16'h8;
17'h149:	data_out=16'h7;
17'h14a:	data_out=16'h8001;
17'h14b:	data_out=16'h8001;
17'h14c:	data_out=16'h8007;
17'h14d:	data_out=16'h8001;
17'h14e:	data_out=16'h8006;
17'h14f:	data_out=16'h8002;
17'h150:	data_out=16'h3;
17'h151:	data_out=16'h5;
17'h152:	data_out=16'h1;
17'h153:	data_out=16'h8002;
17'h154:	data_out=16'h8002;
17'h155:	data_out=16'h2;
17'h156:	data_out=16'h8;
17'h157:	data_out=16'h6;
17'h158:	data_out=16'h3;
17'h159:	data_out=16'h8009;
17'h15a:	data_out=16'h7;
17'h15b:	data_out=16'h8003;
17'h15c:	data_out=16'h8004;
17'h15d:	data_out=16'h3;
17'h15e:	data_out=16'h8005;
17'h15f:	data_out=16'h3;
17'h160:	data_out=16'h0;
17'h161:	data_out=16'h8000;
17'h162:	data_out=16'h8006;
17'h163:	data_out=16'h8005;
17'h164:	data_out=16'h8005;
17'h165:	data_out=16'h6;
17'h166:	data_out=16'h4;
17'h167:	data_out=16'h8005;
17'h168:	data_out=16'h4;
17'h169:	data_out=16'h8007;
17'h16a:	data_out=16'h3;
17'h16b:	data_out=16'h6;
17'h16c:	data_out=16'h2;
17'h16d:	data_out=16'h6;
17'h16e:	data_out=16'h8005;
17'h16f:	data_out=16'h8005;
17'h170:	data_out=16'h2;
17'h171:	data_out=16'h5;
17'h172:	data_out=16'h3;
17'h173:	data_out=16'h8009;
17'h174:	data_out=16'h8003;
17'h175:	data_out=16'h1;
17'h176:	data_out=16'h6;
17'h177:	data_out=16'h9;
17'h178:	data_out=16'h2;
17'h179:	data_out=16'h4;
17'h17a:	data_out=16'h8003;
17'h17b:	data_out=16'h7;
17'h17c:	data_out=16'h8002;
17'h17d:	data_out=16'h1;
17'h17e:	data_out=16'h1;
17'h17f:	data_out=16'h7;
17'h180:	data_out=16'h8008;
17'h181:	data_out=16'h4;
17'h182:	data_out=16'h8007;
17'h183:	data_out=16'h8003;
17'h184:	data_out=16'h0;
17'h185:	data_out=16'h6;
17'h186:	data_out=16'h1;
17'h187:	data_out=16'h8005;
17'h188:	data_out=16'h8;
17'h189:	data_out=16'h8006;
17'h18a:	data_out=16'h8008;
17'h18b:	data_out=16'h1;
17'h18c:	data_out=16'h9;
17'h18d:	data_out=16'h8004;
17'h18e:	data_out=16'h6;
17'h18f:	data_out=16'h2;
17'h190:	data_out=16'h8009;
17'h191:	data_out=16'h8001;
17'h192:	data_out=16'h2;
17'h193:	data_out=16'h8003;
17'h194:	data_out=16'h8008;
17'h195:	data_out=16'h8001;
17'h196:	data_out=16'h8003;
17'h197:	data_out=16'h2;
17'h198:	data_out=16'h8006;
17'h199:	data_out=16'h3;
17'h19a:	data_out=16'h0;
17'h19b:	data_out=16'h1;
17'h19c:	data_out=16'h8005;
17'h19d:	data_out=16'h8008;
17'h19e:	data_out=16'h8001;
17'h19f:	data_out=16'h8004;
17'h1a0:	data_out=16'h5;
17'h1a1:	data_out=16'h1;
17'h1a2:	data_out=16'h2;
17'h1a3:	data_out=16'h8004;
17'h1a4:	data_out=16'h8002;
17'h1a5:	data_out=16'h8007;
17'h1a6:	data_out=16'h0;
17'h1a7:	data_out=16'h8003;
17'h1a8:	data_out=16'h8004;
17'h1a9:	data_out=16'h1;
17'h1aa:	data_out=16'h7;
17'h1ab:	data_out=16'h8004;
17'h1ac:	data_out=16'h6;
17'h1ad:	data_out=16'h4;
17'h1ae:	data_out=16'h7;
17'h1af:	data_out=16'h6;
17'h1b0:	data_out=16'h8006;
17'h1b1:	data_out=16'h8000;
17'h1b2:	data_out=16'h8006;
17'h1b3:	data_out=16'h8005;
17'h1b4:	data_out=16'h8;
17'h1b5:	data_out=16'h0;
17'h1b6:	data_out=16'h6;
17'h1b7:	data_out=16'h8007;
17'h1b8:	data_out=16'h8007;
17'h1b9:	data_out=16'h8003;
17'h1ba:	data_out=16'h3;
17'h1bb:	data_out=16'h8003;
17'h1bc:	data_out=16'h8002;
17'h1bd:	data_out=16'h8007;
17'h1be:	data_out=16'h2;
17'h1bf:	data_out=16'h8006;
17'h1c0:	data_out=16'h4;
17'h1c1:	data_out=16'h8005;
17'h1c2:	data_out=16'h8001;
17'h1c3:	data_out=16'h8008;
17'h1c4:	data_out=16'h8003;
17'h1c5:	data_out=16'h9;
17'h1c6:	data_out=16'h8002;
17'h1c7:	data_out=16'h3;
17'h1c8:	data_out=16'h1;
17'h1c9:	data_out=16'h8004;
17'h1ca:	data_out=16'h8;
17'h1cb:	data_out=16'h8003;
17'h1cc:	data_out=16'h9;
17'h1cd:	data_out=16'h6;
17'h1ce:	data_out=16'h8006;
17'h1cf:	data_out=16'h8007;
17'h1d0:	data_out=16'h8004;
17'h1d1:	data_out=16'h8002;
17'h1d2:	data_out=16'h8003;
17'h1d3:	data_out=16'h8005;
17'h1d4:	data_out=16'h7;
17'h1d5:	data_out=16'h8006;
17'h1d6:	data_out=16'h8003;
17'h1d7:	data_out=16'h8009;
17'h1d8:	data_out=16'h0;
17'h1d9:	data_out=16'h9;
17'h1da:	data_out=16'h8002;
17'h1db:	data_out=16'h8;
17'h1dc:	data_out=16'h8007;
17'h1dd:	data_out=16'h8009;
17'h1de:	data_out=16'h8008;
17'h1df:	data_out=16'h6;
17'h1e0:	data_out=16'h8005;
17'h1e1:	data_out=16'h0;
17'h1e2:	data_out=16'h7;
17'h1e3:	data_out=16'h2;
17'h1e4:	data_out=16'h8000;
17'h1e5:	data_out=16'h8004;
17'h1e6:	data_out=16'h8005;
17'h1e7:	data_out=16'h8009;
17'h1e8:	data_out=16'h1;
17'h1e9:	data_out=16'h8006;
17'h1ea:	data_out=16'h8002;
17'h1eb:	data_out=16'h1;
17'h1ec:	data_out=16'h8009;
17'h1ed:	data_out=16'h1;
17'h1ee:	data_out=16'h4;
17'h1ef:	data_out=16'h8004;
17'h1f0:	data_out=16'h8;
17'h1f1:	data_out=16'h8008;
17'h1f2:	data_out=16'h0;
17'h1f3:	data_out=16'h6;
17'h1f4:	data_out=16'h8005;
17'h1f5:	data_out=16'h6;
17'h1f6:	data_out=16'h6;
17'h1f7:	data_out=16'h5;
17'h1f8:	data_out=16'h6;
17'h1f9:	data_out=16'h8006;
17'h1fa:	data_out=16'h3;
17'h1fb:	data_out=16'h8;
17'h1fc:	data_out=16'h8005;
17'h1fd:	data_out=16'h4;
17'h1fe:	data_out=16'h5;
17'h1ff:	data_out=16'h8001;
17'h200:	data_out=16'h8004;
17'h201:	data_out=16'h3;
17'h202:	data_out=16'h8008;
17'h203:	data_out=16'h4;
17'h204:	data_out=16'h8;
17'h205:	data_out=16'h8004;
17'h206:	data_out=16'h5;
17'h207:	data_out=16'h0;
17'h208:	data_out=16'h8000;
17'h209:	data_out=16'h8007;
17'h20a:	data_out=16'h8008;
17'h20b:	data_out=16'h8000;
17'h20c:	data_out=16'h4;
17'h20d:	data_out=16'h5;
17'h20e:	data_out=16'h5;
17'h20f:	data_out=16'h3;
17'h210:	data_out=16'h6;
17'h211:	data_out=16'h8004;
17'h212:	data_out=16'h8001;
17'h213:	data_out=16'h8008;
17'h214:	data_out=16'h8007;
17'h215:	data_out=16'h8004;
17'h216:	data_out=16'h5;
17'h217:	data_out=16'h8;
17'h218:	data_out=16'h8000;
17'h219:	data_out=16'h8001;
17'h21a:	data_out=16'h7;
17'h21b:	data_out=16'h3;
17'h21c:	data_out=16'h8006;
17'h21d:	data_out=16'h3;
17'h21e:	data_out=16'h8007;
17'h21f:	data_out=16'h8001;
17'h220:	data_out=16'h8004;
17'h221:	data_out=16'h8006;
17'h222:	data_out=16'h8005;
17'h223:	data_out=16'h8005;
17'h224:	data_out=16'h8001;
17'h225:	data_out=16'h8;
17'h226:	data_out=16'h4;
17'h227:	data_out=16'h8;
17'h228:	data_out=16'h8007;
17'h229:	data_out=16'h5;
17'h22a:	data_out=16'h8001;
17'h22b:	data_out=16'h6;
17'h22c:	data_out=16'h1;
17'h22d:	data_out=16'h8006;
17'h22e:	data_out=16'h8000;
17'h22f:	data_out=16'h8002;
17'h230:	data_out=16'h8000;
17'h231:	data_out=16'h8;
17'h232:	data_out=16'h8001;
17'h233:	data_out=16'h2;
17'h234:	data_out=16'h8005;
17'h235:	data_out=16'h8005;
17'h236:	data_out=16'h1;
17'h237:	data_out=16'h4;
17'h238:	data_out=16'h4;
17'h239:	data_out=16'h8001;
17'h23a:	data_out=16'h8002;
17'h23b:	data_out=16'h7;
17'h23c:	data_out=16'h8007;
17'h23d:	data_out=16'h1;
17'h23e:	data_out=16'h8003;
17'h23f:	data_out=16'h8002;
17'h240:	data_out=16'h4;
17'h241:	data_out=16'h1;
17'h242:	data_out=16'h1;
17'h243:	data_out=16'h8006;
17'h244:	data_out=16'h0;
17'h245:	data_out=16'h8004;
17'h246:	data_out=16'h8007;
17'h247:	data_out=16'h2;
17'h248:	data_out=16'h8008;
17'h249:	data_out=16'h1;
17'h24a:	data_out=16'h8001;
17'h24b:	data_out=16'h2;
17'h24c:	data_out=16'h4;
17'h24d:	data_out=16'h8;
17'h24e:	data_out=16'h8009;
17'h24f:	data_out=16'h8005;
17'h250:	data_out=16'h7;
17'h251:	data_out=16'h8001;
17'h252:	data_out=16'h6;
17'h253:	data_out=16'h8007;
17'h254:	data_out=16'h3;
17'h255:	data_out=16'h8002;
17'h256:	data_out=16'h6;
17'h257:	data_out=16'h8002;
17'h258:	data_out=16'h6;
17'h259:	data_out=16'h8005;
17'h25a:	data_out=16'h8004;
17'h25b:	data_out=16'h8;
17'h25c:	data_out=16'h5;
17'h25d:	data_out=16'h2;
17'h25e:	data_out=16'h8003;
17'h25f:	data_out=16'h8000;
17'h260:	data_out=16'h8006;
17'h261:	data_out=16'h7;
17'h262:	data_out=16'h3;
17'h263:	data_out=16'h3;
17'h264:	data_out=16'h8006;
17'h265:	data_out=16'h5;
17'h266:	data_out=16'h8003;
17'h267:	data_out=16'h8005;
17'h268:	data_out=16'h8004;
17'h269:	data_out=16'h5;
17'h26a:	data_out=16'h6;
17'h26b:	data_out=16'h8009;
17'h26c:	data_out=16'h3;
17'h26d:	data_out=16'h6;
17'h26e:	data_out=16'h8005;
17'h26f:	data_out=16'h1;
17'h270:	data_out=16'h8004;
17'h271:	data_out=16'h8008;
17'h272:	data_out=16'h3;
17'h273:	data_out=16'h8;
17'h274:	data_out=16'h8001;
17'h275:	data_out=16'h8000;
17'h276:	data_out=16'h8003;
17'h277:	data_out=16'h8003;
17'h278:	data_out=16'h4;
17'h279:	data_out=16'h2;
17'h27a:	data_out=16'h8004;
17'h27b:	data_out=16'h8000;
17'h27c:	data_out=16'h8005;
17'h27d:	data_out=16'h1;
17'h27e:	data_out=16'h9;
17'h27f:	data_out=16'h8002;
17'h280:	data_out=16'h8001;
17'h281:	data_out=16'h2;
17'h282:	data_out=16'h8008;
17'h283:	data_out=16'h2;
17'h284:	data_out=16'h8002;
17'h285:	data_out=16'h8002;
17'h286:	data_out=16'h6;
17'h287:	data_out=16'h3;
17'h288:	data_out=16'h8007;
17'h289:	data_out=16'h3;
17'h28a:	data_out=16'h3;
17'h28b:	data_out=16'h6;
17'h28c:	data_out=16'h1;
17'h28d:	data_out=16'h8;
17'h28e:	data_out=16'h8002;
17'h28f:	data_out=16'h6;
17'h290:	data_out=16'h9;
17'h291:	data_out=16'h8008;
17'h292:	data_out=16'h5;
17'h293:	data_out=16'h8001;
17'h294:	data_out=16'h1;
17'h295:	data_out=16'h8007;
17'h296:	data_out=16'h5;
17'h297:	data_out=16'h8004;
17'h298:	data_out=16'h4;
17'h299:	data_out=16'h8009;
17'h29a:	data_out=16'h5;
17'h29b:	data_out=16'h8;
17'h29c:	data_out=16'h2;
17'h29d:	data_out=16'h4;
17'h29e:	data_out=16'h8004;
17'h29f:	data_out=16'h8009;
17'h2a0:	data_out=16'h8003;
17'h2a1:	data_out=16'h8002;
17'h2a2:	data_out=16'h3;
17'h2a3:	data_out=16'h4;
17'h2a4:	data_out=16'h4;
17'h2a5:	data_out=16'h8000;
17'h2a6:	data_out=16'h8002;
17'h2a7:	data_out=16'h7;
17'h2a8:	data_out=16'h8006;
17'h2a9:	data_out=16'h8008;
17'h2aa:	data_out=16'h4;
17'h2ab:	data_out=16'h4;
17'h2ac:	data_out=16'h8;
17'h2ad:	data_out=16'h8008;
17'h2ae:	data_out=16'h1;
17'h2af:	data_out=16'h8;
17'h2b0:	data_out=16'h8007;
17'h2b1:	data_out=16'h8003;
17'h2b2:	data_out=16'h8002;
17'h2b3:	data_out=16'h3;
17'h2b4:	data_out=16'h8001;
17'h2b5:	data_out=16'h8006;
17'h2b6:	data_out=16'h8;
17'h2b7:	data_out=16'h8006;
17'h2b8:	data_out=16'h8006;
17'h2b9:	data_out=16'h3;
17'h2ba:	data_out=16'h8007;
17'h2bb:	data_out=16'h4;
17'h2bc:	data_out=16'h8002;
17'h2bd:	data_out=16'h8002;
17'h2be:	data_out=16'h5;
17'h2bf:	data_out=16'h4;
17'h2c0:	data_out=16'h5;
17'h2c1:	data_out=16'h8002;
17'h2c2:	data_out=16'h8001;
17'h2c3:	data_out=16'h0;
17'h2c4:	data_out=16'h7;
17'h2c5:	data_out=16'h6;
17'h2c6:	data_out=16'h8002;
17'h2c7:	data_out=16'h8008;
17'h2c8:	data_out=16'h7;
17'h2c9:	data_out=16'h8008;
17'h2ca:	data_out=16'h5;
17'h2cb:	data_out=16'h6;
17'h2cc:	data_out=16'h8006;
17'h2cd:	data_out=16'h8003;
17'h2ce:	data_out=16'h5;
17'h2cf:	data_out=16'h8004;
17'h2d0:	data_out=16'h3;
17'h2d1:	data_out=16'h8006;
17'h2d2:	data_out=16'h8;
17'h2d3:	data_out=16'h8007;
17'h2d4:	data_out=16'h8004;
17'h2d5:	data_out=16'h7;
17'h2d6:	data_out=16'h8004;
17'h2d7:	data_out=16'h8001;
17'h2d8:	data_out=16'h0;
17'h2d9:	data_out=16'h8002;
17'h2da:	data_out=16'h8005;
17'h2db:	data_out=16'h7;
17'h2dc:	data_out=16'h5;
17'h2dd:	data_out=16'h9;
17'h2de:	data_out=16'h2;
17'h2df:	data_out=16'h1;
17'h2e0:	data_out=16'h8002;
17'h2e1:	data_out=16'h8008;
17'h2e2:	data_out=16'h8008;
17'h2e3:	data_out=16'h8004;
17'h2e4:	data_out=16'h7;
17'h2e5:	data_out=16'h8001;
17'h2e6:	data_out=16'h8003;
17'h2e7:	data_out=16'h4;
17'h2e8:	data_out=16'h1;
17'h2e9:	data_out=16'h8007;
17'h2ea:	data_out=16'h1;
17'h2eb:	data_out=16'h4;
17'h2ec:	data_out=16'h8001;
17'h2ed:	data_out=16'h8003;
17'h2ee:	data_out=16'h9;
17'h2ef:	data_out=16'h8007;
17'h2f0:	data_out=16'h8000;
17'h2f1:	data_out=16'h8;
17'h2f2:	data_out=16'h8005;
17'h2f3:	data_out=16'h5;
17'h2f4:	data_out=16'h5;
17'h2f5:	data_out=16'h1;
17'h2f6:	data_out=16'h8005;
17'h2f7:	data_out=16'h8004;
17'h2f8:	data_out=16'h8;
17'h2f9:	data_out=16'h8001;
17'h2fa:	data_out=16'h8005;
17'h2fb:	data_out=16'h4;
17'h2fc:	data_out=16'h8001;
17'h2fd:	data_out=16'h6;
17'h2fe:	data_out=16'h8004;
17'h2ff:	data_out=16'h6;
17'h300:	data_out=16'h7;
17'h301:	data_out=16'h8003;
17'h302:	data_out=16'h8007;
17'h303:	data_out=16'h5;
17'h304:	data_out=16'h5;
17'h305:	data_out=16'h8000;
17'h306:	data_out=16'h0;
17'h307:	data_out=16'h8004;
17'h308:	data_out=16'h2;
17'h309:	data_out=16'h8008;
17'h30a:	data_out=16'h8009;
17'h30b:	data_out=16'h8008;
17'h30c:	data_out=16'h8002;
17'h30d:	data_out=16'h9;
17'h30e:	data_out=16'h8006;
17'h30f:	data_out=16'h7;
17'h310:	data_out=16'h7;
17'h311:	data_out=16'h8002;
17'h312:	data_out=16'h3;
17'h313:	data_out=16'h3;
17'h314:	data_out=16'h8;
17'h315:	data_out=16'h7;
17'h316:	data_out=16'h9;
17'h317:	data_out=16'h6;
17'h318:	data_out=16'h8003;
17'h319:	data_out=16'h8006;
17'h31a:	data_out=16'h1;
17'h31b:	data_out=16'h5;
17'h31c:	data_out=16'h8009;
17'h31d:	data_out=16'h6;
17'h31e:	data_out=16'h2;
17'h31f:	data_out=16'h8;
17'h320:	data_out=16'h8007;
17'h321:	data_out=16'h4;
17'h322:	data_out=16'h3;
17'h323:	data_out=16'h7;
17'h324:	data_out=16'h8005;
17'h325:	data_out=16'h8006;
17'h326:	data_out=16'h8005;
17'h327:	data_out=16'h6;
17'h328:	data_out=16'h8004;
17'h329:	data_out=16'h8005;
17'h32a:	data_out=16'h7;
17'h32b:	data_out=16'h3;
17'h32c:	data_out=16'h8006;
17'h32d:	data_out=16'h8008;
17'h32e:	data_out=16'h1;
17'h32f:	data_out=16'h8007;
17'h330:	data_out=16'h8001;
17'h331:	data_out=16'h8005;
17'h332:	data_out=16'h5;
17'h333:	data_out=16'h8002;
17'h334:	data_out=16'h8007;
17'h335:	data_out=16'h5;
17'h336:	data_out=16'h8005;
17'h337:	data_out=16'h8001;
17'h338:	data_out=16'h9;
17'h339:	data_out=16'h5;
17'h33a:	data_out=16'h8005;
17'h33b:	data_out=16'h8009;
17'h33c:	data_out=16'h2;
17'h33d:	data_out=16'h6;
17'h33e:	data_out=16'h8;
17'h33f:	data_out=16'h4;
17'h340:	data_out=16'h2;
17'h341:	data_out=16'h2;
17'h342:	data_out=16'h2;
17'h343:	data_out=16'h5;
17'h344:	data_out=16'h6;
17'h345:	data_out=16'h6;
17'h346:	data_out=16'h2;
17'h347:	data_out=16'h8008;
17'h348:	data_out=16'h8008;
17'h349:	data_out=16'h8001;
17'h34a:	data_out=16'h4;
17'h34b:	data_out=16'h8005;
17'h34c:	data_out=16'h8000;
17'h34d:	data_out=16'h8004;
17'h34e:	data_out=16'h8003;
17'h34f:	data_out=16'h8;
17'h350:	data_out=16'h8000;
17'h351:	data_out=16'h8007;
17'h352:	data_out=16'h8003;
17'h353:	data_out=16'h2;
17'h354:	data_out=16'h7;
17'h355:	data_out=16'h1;
17'h356:	data_out=16'h8008;
17'h357:	data_out=16'h7;
17'h358:	data_out=16'h8003;
17'h359:	data_out=16'h8004;
17'h35a:	data_out=16'h7;
17'h35b:	data_out=16'h8;
17'h35c:	data_out=16'h8006;
17'h35d:	data_out=16'h6;
17'h35e:	data_out=16'h3;
17'h35f:	data_out=16'h4;
17'h360:	data_out=16'h8001;
17'h361:	data_out=16'h8004;
17'h362:	data_out=16'h0;
17'h363:	data_out=16'h8005;
17'h364:	data_out=16'h8007;
17'h365:	data_out=16'h8007;
17'h366:	data_out=16'h8004;
17'h367:	data_out=16'h8006;
17'h368:	data_out=16'h1;
17'h369:	data_out=16'h8008;
17'h36a:	data_out=16'h8002;
17'h36b:	data_out=16'h8008;
17'h36c:	data_out=16'h8003;
17'h36d:	data_out=16'h5;
17'h36e:	data_out=16'h9;
17'h36f:	data_out=16'h6;
17'h370:	data_out=16'h7;
17'h371:	data_out=16'h8004;
17'h372:	data_out=16'h8002;
17'h373:	data_out=16'h5;
17'h374:	data_out=16'h6;
17'h375:	data_out=16'h8001;
17'h376:	data_out=16'h3;
17'h377:	data_out=16'h8006;
17'h378:	data_out=16'h5;
17'h379:	data_out=16'h1;
17'h37a:	data_out=16'h8008;
17'h37b:	data_out=16'h7;
17'h37c:	data_out=16'h8003;
17'h37d:	data_out=16'h4;
17'h37e:	data_out=16'h3;
17'h37f:	data_out=16'h5;
17'h380:	data_out=16'h8009;
17'h381:	data_out=16'h8006;
17'h382:	data_out=16'h9;
17'h383:	data_out=16'h8006;
17'h384:	data_out=16'h8004;
17'h385:	data_out=16'h8004;
17'h386:	data_out=16'h8003;
17'h387:	data_out=16'h6;
17'h388:	data_out=16'h8003;
17'h389:	data_out=16'h5;
17'h38a:	data_out=16'h7;
17'h38b:	data_out=16'h3;
17'h38c:	data_out=16'h0;
17'h38d:	data_out=16'h7;
17'h38e:	data_out=16'h8001;
17'h38f:	data_out=16'h8002;
17'h390:	data_out=16'h8006;
17'h391:	data_out=16'h7;
17'h392:	data_out=16'h8006;
17'h393:	data_out=16'h9;
17'h394:	data_out=16'h8003;
17'h395:	data_out=16'h6;
17'h396:	data_out=16'h8006;
17'h397:	data_out=16'h8008;
17'h398:	data_out=16'h8003;
17'h399:	data_out=16'h8005;
17'h39a:	data_out=16'h9;
17'h39b:	data_out=16'h3;
17'h39c:	data_out=16'h9;
17'h39d:	data_out=16'h2;
17'h39e:	data_out=16'h8001;
17'h39f:	data_out=16'h8009;
17'h3a0:	data_out=16'h5;
17'h3a1:	data_out=16'h8001;
17'h3a2:	data_out=16'h8006;
17'h3a3:	data_out=16'h8008;
17'h3a4:	data_out=16'h4;
17'h3a5:	data_out=16'h0;
17'h3a6:	data_out=16'h7;
17'h3a7:	data_out=16'h8008;
17'h3a8:	data_out=16'h8004;
17'h3a9:	data_out=16'h5;
17'h3aa:	data_out=16'h4;
17'h3ab:	data_out=16'h6;
17'h3ac:	data_out=16'h2;
17'h3ad:	data_out=16'h8005;
17'h3ae:	data_out=16'h8006;
17'h3af:	data_out=16'h5;
17'h3b0:	data_out=16'h8008;
17'h3b1:	data_out=16'h8003;
17'h3b2:	data_out=16'h5;
17'h3b3:	data_out=16'h8002;
17'h3b4:	data_out=16'h8007;
17'h3b5:	data_out=16'h7;
17'h3b6:	data_out=16'h8000;
17'h3b7:	data_out=16'h8000;
17'h3b8:	data_out=16'h8007;
17'h3b9:	data_out=16'h8000;
17'h3ba:	data_out=16'h8006;
17'h3bb:	data_out=16'h8007;
17'h3bc:	data_out=16'h8007;
17'h3bd:	data_out=16'h2;
17'h3be:	data_out=16'h8007;
17'h3bf:	data_out=16'h7;
17'h3c0:	data_out=16'h8009;
17'h3c1:	data_out=16'h8004;
17'h3c2:	data_out=16'h8;
17'h3c3:	data_out=16'h5;
17'h3c4:	data_out=16'h6;
17'h3c5:	data_out=16'h6;
17'h3c6:	data_out=16'h6;
17'h3c7:	data_out=16'h8007;
17'h3c8:	data_out=16'h1;
17'h3c9:	data_out=16'h2;
17'h3ca:	data_out=16'h8;
17'h3cb:	data_out=16'h8006;
17'h3cc:	data_out=16'h5;
17'h3cd:	data_out=16'h8007;
17'h3ce:	data_out=16'h8;
17'h3cf:	data_out=16'h7;
17'h3d0:	data_out=16'h8001;
17'h3d1:	data_out=16'h3;
17'h3d2:	data_out=16'h8004;
17'h3d3:	data_out=16'h1;
17'h3d4:	data_out=16'h2;
17'h3d5:	data_out=16'h5;
17'h3d6:	data_out=16'h8008;
17'h3d7:	data_out=16'h4;
17'h3d8:	data_out=16'h8005;
17'h3d9:	data_out=16'h8005;
17'h3da:	data_out=16'h6;
17'h3db:	data_out=16'h8003;
17'h3dc:	data_out=16'h6;
17'h3dd:	data_out=16'h8;
17'h3de:	data_out=16'h8005;
17'h3df:	data_out=16'h6;
17'h3e0:	data_out=16'h8004;
17'h3e1:	data_out=16'h8006;
17'h3e2:	data_out=16'h2;
17'h3e3:	data_out=16'h8008;
17'h3e4:	data_out=16'h9;
17'h3e5:	data_out=16'h8001;
17'h3e6:	data_out=16'h8005;
17'h3e7:	data_out=16'h1;
17'h3e8:	data_out=16'h8008;
17'h3e9:	data_out=16'h8007;
17'h3ea:	data_out=16'h4;
17'h3eb:	data_out=16'h6;
17'h3ec:	data_out=16'h8005;
17'h3ed:	data_out=16'h3;
17'h3ee:	data_out=16'h4;
17'h3ef:	data_out=16'h3;
17'h3f0:	data_out=16'h8003;
17'h3f1:	data_out=16'h9;
17'h3f2:	data_out=16'h8005;
17'h3f3:	data_out=16'h8;
17'h3f4:	data_out=16'h5;
17'h3f5:	data_out=16'h8004;
17'h3f6:	data_out=16'h3;
17'h3f7:	data_out=16'h9;
17'h3f8:	data_out=16'h0;
17'h3f9:	data_out=16'h8000;
17'h3fa:	data_out=16'h8003;
17'h3fb:	data_out=16'h8003;
17'h3fc:	data_out=16'h8001;
17'h3fd:	data_out=16'h1;
17'h3fe:	data_out=16'h8006;
17'h3ff:	data_out=16'h4;
17'h400:	data_out=16'h4;
17'h401:	data_out=16'h5;
17'h402:	data_out=16'h5;
17'h403:	data_out=16'h4;
17'h404:	data_out=16'h8005;
17'h405:	data_out=16'h8009;
17'h406:	data_out=16'h8005;
17'h407:	data_out=16'h8005;
17'h408:	data_out=16'h8007;
17'h409:	data_out=16'h8;
17'h40a:	data_out=16'h8008;
17'h40b:	data_out=16'h8003;
17'h40c:	data_out=16'h2;
17'h40d:	data_out=16'h5;
17'h40e:	data_out=16'h8009;
17'h40f:	data_out=16'h8;
17'h410:	data_out=16'h5;
17'h411:	data_out=16'h8004;
17'h412:	data_out=16'h7;
17'h413:	data_out=16'h0;
17'h414:	data_out=16'h1;
17'h415:	data_out=16'h1;
17'h416:	data_out=16'h0;
17'h417:	data_out=16'h8008;
17'h418:	data_out=16'h8008;
17'h419:	data_out=16'h6;
17'h41a:	data_out=16'h8002;
17'h41b:	data_out=16'h8000;
17'h41c:	data_out=16'h8001;
17'h41d:	data_out=16'h1;
17'h41e:	data_out=16'h8005;
17'h41f:	data_out=16'h8006;
17'h420:	data_out=16'h8004;
17'h421:	data_out=16'h8009;
17'h422:	data_out=16'h6;
17'h423:	data_out=16'h8000;
17'h424:	data_out=16'h8009;
17'h425:	data_out=16'h8007;
17'h426:	data_out=16'h4;
17'h427:	data_out=16'h8006;
17'h428:	data_out=16'h8008;
17'h429:	data_out=16'h6;
17'h42a:	data_out=16'h8000;
17'h42b:	data_out=16'h3;
17'h42c:	data_out=16'h2;
17'h42d:	data_out=16'h0;
17'h42e:	data_out=16'h2;
17'h42f:	data_out=16'h8002;
17'h430:	data_out=16'h5;
17'h431:	data_out=16'h0;
17'h432:	data_out=16'h7;
17'h433:	data_out=16'h8003;
17'h434:	data_out=16'h8008;
17'h435:	data_out=16'h8002;
17'h436:	data_out=16'h8001;
17'h437:	data_out=16'h8007;
17'h438:	data_out=16'h8004;
17'h439:	data_out=16'h6;
17'h43a:	data_out=16'h2;
17'h43b:	data_out=16'h3;
17'h43c:	data_out=16'h8002;
17'h43d:	data_out=16'h6;
17'h43e:	data_out=16'h6;
17'h43f:	data_out=16'h3;
17'h440:	data_out=16'h6;
17'h441:	data_out=16'h3;
17'h442:	data_out=16'h8006;
17'h443:	data_out=16'h6;
17'h444:	data_out=16'h5;
17'h445:	data_out=16'h7;
17'h446:	data_out=16'h9;
17'h447:	data_out=16'h6;
17'h448:	data_out=16'h4;
17'h449:	data_out=16'h8000;
17'h44a:	data_out=16'h0;
17'h44b:	data_out=16'h8004;
17'h44c:	data_out=16'h8009;
17'h44d:	data_out=16'h8007;
17'h44e:	data_out=16'h3;
17'h44f:	data_out=16'h5;
17'h450:	data_out=16'h3;
17'h451:	data_out=16'h1;
17'h452:	data_out=16'h8006;
17'h453:	data_out=16'h4;
17'h454:	data_out=16'h8;
17'h455:	data_out=16'h1;
17'h456:	data_out=16'h6;
17'h457:	data_out=16'h8005;
17'h458:	data_out=16'h8002;
17'h459:	data_out=16'h8001;
17'h45a:	data_out=16'h7;
17'h45b:	data_out=16'h5;
17'h45c:	data_out=16'h8005;
17'h45d:	data_out=16'h4;
17'h45e:	data_out=16'h8001;
17'h45f:	data_out=16'h8008;
17'h460:	data_out=16'h8002;
17'h461:	data_out=16'h2;
17'h462:	data_out=16'h8;
17'h463:	data_out=16'h8006;
17'h464:	data_out=16'h8000;
17'h465:	data_out=16'h7;
17'h466:	data_out=16'h8009;
17'h467:	data_out=16'h8006;
17'h468:	data_out=16'h8002;
17'h469:	data_out=16'h0;
17'h46a:	data_out=16'h0;
17'h46b:	data_out=16'h8002;
17'h46c:	data_out=16'h3;
17'h46d:	data_out=16'h8006;
17'h46e:	data_out=16'h8006;
17'h46f:	data_out=16'h8003;
17'h470:	data_out=16'h4;
17'h471:	data_out=16'h8003;
17'h472:	data_out=16'h8008;
17'h473:	data_out=16'h3;
17'h474:	data_out=16'h8;
17'h475:	data_out=16'h7;
17'h476:	data_out=16'h7;
17'h477:	data_out=16'h8003;
17'h478:	data_out=16'h8004;
17'h479:	data_out=16'h5;
17'h47a:	data_out=16'h8007;
17'h47b:	data_out=16'h1;
17'h47c:	data_out=16'h0;
17'h47d:	data_out=16'h0;
17'h47e:	data_out=16'h2;
17'h47f:	data_out=16'h8;
17'h480:	data_out=16'h8007;
17'h481:	data_out=16'h1;
17'h482:	data_out=16'h8007;
17'h483:	data_out=16'h2;
17'h484:	data_out=16'h8001;
17'h485:	data_out=16'h8007;
17'h486:	data_out=16'h5;
17'h487:	data_out=16'h6;
17'h488:	data_out=16'h2;
17'h489:	data_out=16'h8004;
17'h48a:	data_out=16'h8005;
17'h48b:	data_out=16'h8004;
17'h48c:	data_out=16'h8001;
17'h48d:	data_out=16'h8001;
17'h48e:	data_out=16'h2;
17'h48f:	data_out=16'h8006;
17'h490:	data_out=16'h5;
17'h491:	data_out=16'h3;
17'h492:	data_out=16'h7;
17'h493:	data_out=16'h4;
17'h494:	data_out=16'h1;
17'h495:	data_out=16'h5;
17'h496:	data_out=16'h8008;
17'h497:	data_out=16'h6;
17'h498:	data_out=16'h1;
17'h499:	data_out=16'h8006;
17'h49a:	data_out=16'h8002;
17'h49b:	data_out=16'h8008;
17'h49c:	data_out=16'h3;
17'h49d:	data_out=16'h9;
17'h49e:	data_out=16'h8009;
17'h49f:	data_out=16'h5;
17'h4a0:	data_out=16'h1;
17'h4a1:	data_out=16'h8007;
17'h4a2:	data_out=16'h8003;
17'h4a3:	data_out=16'h9;
17'h4a4:	data_out=16'h8006;
17'h4a5:	data_out=16'h8007;
17'h4a6:	data_out=16'h6;
17'h4a7:	data_out=16'h6;
17'h4a8:	data_out=16'h8002;
17'h4a9:	data_out=16'h8008;
17'h4aa:	data_out=16'h8007;
17'h4ab:	data_out=16'h7;
17'h4ac:	data_out=16'h0;
17'h4ad:	data_out=16'h4;
17'h4ae:	data_out=16'h8008;
17'h4af:	data_out=16'h8003;
17'h4b0:	data_out=16'h8002;
17'h4b1:	data_out=16'h7;
17'h4b2:	data_out=16'h8009;
17'h4b3:	data_out=16'h8;
17'h4b4:	data_out=16'h3;
17'h4b5:	data_out=16'h8008;
17'h4b6:	data_out=16'h5;
17'h4b7:	data_out=16'h8005;
17'h4b8:	data_out=16'h8005;
17'h4b9:	data_out=16'h8007;
17'h4ba:	data_out=16'h8003;
17'h4bb:	data_out=16'h7;
17'h4bc:	data_out=16'h8007;
17'h4bd:	data_out=16'h8003;
17'h4be:	data_out=16'h3;
17'h4bf:	data_out=16'h3;
17'h4c0:	data_out=16'h8001;
17'h4c1:	data_out=16'h8009;
17'h4c2:	data_out=16'h3;
17'h4c3:	data_out=16'h2;
17'h4c4:	data_out=16'h8006;
17'h4c5:	data_out=16'h8000;
17'h4c6:	data_out=16'h8001;
17'h4c7:	data_out=16'h1;
17'h4c8:	data_out=16'h1;
17'h4c9:	data_out=16'h2;
17'h4ca:	data_out=16'h8001;
17'h4cb:	data_out=16'h8007;
17'h4cc:	data_out=16'h8003;
17'h4cd:	data_out=16'h8000;
17'h4ce:	data_out=16'h8002;
17'h4cf:	data_out=16'h4;
17'h4d0:	data_out=16'h8002;
17'h4d1:	data_out=16'h8001;
17'h4d2:	data_out=16'h3;
17'h4d3:	data_out=16'h8008;
17'h4d4:	data_out=16'h1;
17'h4d5:	data_out=16'h8001;
17'h4d6:	data_out=16'h8003;
17'h4d7:	data_out=16'h5;
17'h4d8:	data_out=16'h1;
17'h4d9:	data_out=16'h3;
17'h4da:	data_out=16'h3;
17'h4db:	data_out=16'h4;
17'h4dc:	data_out=16'h8009;
17'h4dd:	data_out=16'h8003;
17'h4de:	data_out=16'h8002;
17'h4df:	data_out=16'h8001;
17'h4e0:	data_out=16'h8002;
17'h4e1:	data_out=16'h8008;
17'h4e2:	data_out=16'h8008;
17'h4e3:	data_out=16'h1;
17'h4e4:	data_out=16'h1;
17'h4e5:	data_out=16'h1;
17'h4e6:	data_out=16'h8007;
17'h4e7:	data_out=16'h8007;
17'h4e8:	data_out=16'h8007;
17'h4e9:	data_out=16'h1;
17'h4ea:	data_out=16'h8005;
17'h4eb:	data_out=16'h8001;
17'h4ec:	data_out=16'h8009;
17'h4ed:	data_out=16'h2;
17'h4ee:	data_out=16'h8006;
17'h4ef:	data_out=16'h8002;
17'h4f0:	data_out=16'h8008;
17'h4f1:	data_out=16'h7;
17'h4f2:	data_out=16'h8000;
17'h4f3:	data_out=16'h2;
17'h4f4:	data_out=16'h8004;
17'h4f5:	data_out=16'h6;
17'h4f6:	data_out=16'h8002;
17'h4f7:	data_out=16'h7;
17'h4f8:	data_out=16'h8001;
17'h4f9:	data_out=16'h8008;
17'h4fa:	data_out=16'h1;
17'h4fb:	data_out=16'h8001;
17'h4fc:	data_out=16'h8002;
17'h4fd:	data_out=16'h8;
17'h4fe:	data_out=16'h7;
17'h4ff:	data_out=16'h5;
17'h500:	data_out=16'h9;
17'h501:	data_out=16'h9;
17'h502:	data_out=16'h8004;
17'h503:	data_out=16'h0;
17'h504:	data_out=16'h0;
17'h505:	data_out=16'h8002;
17'h506:	data_out=16'h2;
17'h507:	data_out=16'h3;
17'h508:	data_out=16'h8;
17'h509:	data_out=16'h6;
17'h50a:	data_out=16'h8007;
17'h50b:	data_out=16'h9;
17'h50c:	data_out=16'h8001;
17'h50d:	data_out=16'h8004;
17'h50e:	data_out=16'h8002;
17'h50f:	data_out=16'h1;
17'h510:	data_out=16'h8006;
17'h511:	data_out=16'h7;
17'h512:	data_out=16'h8007;
17'h513:	data_out=16'h8001;
17'h514:	data_out=16'h3;
17'h515:	data_out=16'h0;
17'h516:	data_out=16'h8003;
17'h517:	data_out=16'h8006;
17'h518:	data_out=16'h1;
17'h519:	data_out=16'h7;
17'h51a:	data_out=16'h2;
17'h51b:	data_out=16'h8;
17'h51c:	data_out=16'h6;
17'h51d:	data_out=16'h0;
17'h51e:	data_out=16'h3;
17'h51f:	data_out=16'h5;
17'h520:	data_out=16'h8000;
17'h521:	data_out=16'h8;
17'h522:	data_out=16'h8004;
17'h523:	data_out=16'h8009;
17'h524:	data_out=16'h8003;
17'h525:	data_out=16'h7;
17'h526:	data_out=16'h3;
17'h527:	data_out=16'h8003;
17'h528:	data_out=16'h4;
17'h529:	data_out=16'h5;
17'h52a:	data_out=16'h8004;
17'h52b:	data_out=16'h8006;
17'h52c:	data_out=16'h8008;
17'h52d:	data_out=16'h4;
17'h52e:	data_out=16'h4;
17'h52f:	data_out=16'h8005;
17'h530:	data_out=16'h1;
17'h531:	data_out=16'h7;
17'h532:	data_out=16'h3;
17'h533:	data_out=16'h8004;
17'h534:	data_out=16'h8002;
17'h535:	data_out=16'h9;
17'h536:	data_out=16'h8002;
17'h537:	data_out=16'h8;
17'h538:	data_out=16'h6;
17'h539:	data_out=16'h8009;
17'h53a:	data_out=16'h7;
17'h53b:	data_out=16'h3;
17'h53c:	data_out=16'h1;
17'h53d:	data_out=16'h1;
17'h53e:	data_out=16'h8001;
17'h53f:	data_out=16'h8008;
17'h540:	data_out=16'h0;
17'h541:	data_out=16'h4;
17'h542:	data_out=16'h8008;
17'h543:	data_out=16'h7;
17'h544:	data_out=16'h2;
17'h545:	data_out=16'h4;
17'h546:	data_out=16'h8006;
17'h547:	data_out=16'h8003;
17'h548:	data_out=16'h8001;
17'h549:	data_out=16'h8000;
17'h54a:	data_out=16'h0;
17'h54b:	data_out=16'h0;
17'h54c:	data_out=16'h8006;
17'h54d:	data_out=16'h8005;
17'h54e:	data_out=16'h4;
17'h54f:	data_out=16'h4;
17'h550:	data_out=16'h8007;
17'h551:	data_out=16'h8002;
17'h552:	data_out=16'h8009;
17'h553:	data_out=16'h8000;
17'h554:	data_out=16'h8003;
17'h555:	data_out=16'h8002;
17'h556:	data_out=16'h8002;
17'h557:	data_out=16'h8006;
17'h558:	data_out=16'h8001;
17'h559:	data_out=16'h8004;
17'h55a:	data_out=16'h6;
17'h55b:	data_out=16'h9;
17'h55c:	data_out=16'h6;
17'h55d:	data_out=16'h8004;
17'h55e:	data_out=16'h8009;
17'h55f:	data_out=16'h8003;
17'h560:	data_out=16'h8;
17'h561:	data_out=16'h8008;
17'h562:	data_out=16'h8005;
17'h563:	data_out=16'h1;
17'h564:	data_out=16'h5;
17'h565:	data_out=16'h8002;
17'h566:	data_out=16'h7;
17'h567:	data_out=16'h8004;
17'h568:	data_out=16'h7;
17'h569:	data_out=16'h8002;
17'h56a:	data_out=16'h5;
17'h56b:	data_out=16'h8008;
17'h56c:	data_out=16'h3;
17'h56d:	data_out=16'h8000;
17'h56e:	data_out=16'h6;
17'h56f:	data_out=16'h5;
17'h570:	data_out=16'h6;
17'h571:	data_out=16'h6;
17'h572:	data_out=16'h8005;
17'h573:	data_out=16'h8006;
17'h574:	data_out=16'h8005;
17'h575:	data_out=16'h3;
17'h576:	data_out=16'h8002;
17'h577:	data_out=16'h3;
17'h578:	data_out=16'h8;
17'h579:	data_out=16'h8005;
17'h57a:	data_out=16'h3;
17'h57b:	data_out=16'h5;
17'h57c:	data_out=16'h8000;
17'h57d:	data_out=16'h3;
17'h57e:	data_out=16'h8007;
17'h57f:	data_out=16'h8001;
17'h580:	data_out=16'h5;
17'h581:	data_out=16'h8003;
17'h582:	data_out=16'h9;
17'h583:	data_out=16'h1;
17'h584:	data_out=16'h4;
17'h585:	data_out=16'h7;
17'h586:	data_out=16'h6;
17'h587:	data_out=16'h2;
17'h588:	data_out=16'h8004;
17'h589:	data_out=16'h1;
17'h58a:	data_out=16'h3;
17'h58b:	data_out=16'h8;
17'h58c:	data_out=16'h8008;
17'h58d:	data_out=16'h8000;
17'h58e:	data_out=16'h3;
17'h58f:	data_out=16'h7;
17'h590:	data_out=16'h8004;
17'h591:	data_out=16'h7;
17'h592:	data_out=16'h8007;
17'h593:	data_out=16'h0;
17'h594:	data_out=16'h1;
17'h595:	data_out=16'h8000;
17'h596:	data_out=16'h8006;
17'h597:	data_out=16'h8000;
17'h598:	data_out=16'h4;
17'h599:	data_out=16'h6;
17'h59a:	data_out=16'h8004;
17'h59b:	data_out=16'h8006;
17'h59c:	data_out=16'h8000;
17'h59d:	data_out=16'h8002;
17'h59e:	data_out=16'h2;
17'h59f:	data_out=16'h8005;
17'h5a0:	data_out=16'h4;
17'h5a1:	data_out=16'h2;
17'h5a2:	data_out=16'h5;
17'h5a3:	data_out=16'h8001;
17'h5a4:	data_out=16'h8000;
17'h5a5:	data_out=16'h2;
17'h5a6:	data_out=16'h8008;
17'h5a7:	data_out=16'h5;
17'h5a8:	data_out=16'h8006;
17'h5a9:	data_out=16'h5;
17'h5aa:	data_out=16'h3;
17'h5ab:	data_out=16'h8005;
17'h5ac:	data_out=16'h8004;
17'h5ad:	data_out=16'h8003;
17'h5ae:	data_out=16'h8007;
17'h5af:	data_out=16'h1;
17'h5b0:	data_out=16'h8004;
17'h5b1:	data_out=16'h8006;
17'h5b2:	data_out=16'h8008;
17'h5b3:	data_out=16'h6;
17'h5b4:	data_out=16'h3;
17'h5b5:	data_out=16'h8004;
17'h5b6:	data_out=16'h8004;
17'h5b7:	data_out=16'h8002;
17'h5b8:	data_out=16'h8007;
17'h5b9:	data_out=16'h1;
17'h5ba:	data_out=16'h1;
17'h5bb:	data_out=16'h2;
17'h5bc:	data_out=16'h8;
17'h5bd:	data_out=16'h8005;
17'h5be:	data_out=16'h6;
17'h5bf:	data_out=16'h3;
17'h5c0:	data_out=16'h6;
17'h5c1:	data_out=16'h2;
17'h5c2:	data_out=16'h8007;
17'h5c3:	data_out=16'h8004;
17'h5c4:	data_out=16'h8005;
17'h5c5:	data_out=16'h8006;
17'h5c6:	data_out=16'h8008;
17'h5c7:	data_out=16'h8002;
17'h5c8:	data_out=16'h8;
17'h5c9:	data_out=16'h4;
17'h5ca:	data_out=16'h2;
17'h5cb:	data_out=16'h8005;
17'h5cc:	data_out=16'h8007;
17'h5cd:	data_out=16'h4;
17'h5ce:	data_out=16'h5;
17'h5cf:	data_out=16'h8003;
17'h5d0:	data_out=16'h7;
17'h5d1:	data_out=16'h7;
17'h5d2:	data_out=16'h8006;
17'h5d3:	data_out=16'h1;
17'h5d4:	data_out=16'h8006;
17'h5d5:	data_out=16'h8001;
17'h5d6:	data_out=16'h8;
17'h5d7:	data_out=16'h8005;
17'h5d8:	data_out=16'h8009;
17'h5d9:	data_out=16'h1;
17'h5da:	data_out=16'h6;
17'h5db:	data_out=16'h8;
17'h5dc:	data_out=16'h5;
17'h5dd:	data_out=16'h3;
17'h5de:	data_out=16'h2;
17'h5df:	data_out=16'h1;
17'h5e0:	data_out=16'h8004;
17'h5e1:	data_out=16'h3;
17'h5e2:	data_out=16'h7;
17'h5e3:	data_out=16'h0;
17'h5e4:	data_out=16'h7;
17'h5e5:	data_out=16'h8;
17'h5e6:	data_out=16'h7;
17'h5e7:	data_out=16'h6;
17'h5e8:	data_out=16'h3;
17'h5e9:	data_out=16'h0;
17'h5ea:	data_out=16'h8008;
17'h5eb:	data_out=16'h5;
17'h5ec:	data_out=16'h8006;
17'h5ed:	data_out=16'h7;
17'h5ee:	data_out=16'h8007;
17'h5ef:	data_out=16'h8008;
17'h5f0:	data_out=16'h4;
17'h5f1:	data_out=16'h8004;
17'h5f2:	data_out=16'h3;
17'h5f3:	data_out=16'h7;
17'h5f4:	data_out=16'h4;
17'h5f5:	data_out=16'h2;
17'h5f6:	data_out=16'h8007;
17'h5f7:	data_out=16'h4;
17'h5f8:	data_out=16'h8006;
17'h5f9:	data_out=16'h8;
17'h5fa:	data_out=16'h3;
17'h5fb:	data_out=16'h8;
17'h5fc:	data_out=16'h2;
17'h5fd:	data_out=16'h8005;
17'h5fe:	data_out=16'h8000;
17'h5ff:	data_out=16'h8;
17'h600:	data_out=16'h4f;
17'h601:	data_out=16'h59;
17'h602:	data_out=16'hf;
17'h603:	data_out=16'h4c;
17'h604:	data_out=16'h56;
17'h605:	data_out=16'h55;
17'h606:	data_out=16'h8000;
17'h607:	data_out=16'h8002;
17'h608:	data_out=16'h4a;
17'h609:	data_out=16'h801c;
17'h60a:	data_out=16'h6f;
17'h60b:	data_out=16'h40;
17'h60c:	data_out=16'h4a;
17'h60d:	data_out=16'h13;
17'h60e:	data_out=16'h8004;
17'h60f:	data_out=16'h800c;
17'h610:	data_out=16'hd;
17'h611:	data_out=16'h5f;
17'h612:	data_out=16'h8032;
17'h613:	data_out=16'h51;
17'h614:	data_out=16'ha;
17'h615:	data_out=16'h19;
17'h616:	data_out=16'h2f;
17'h617:	data_out=16'h1d;
17'h618:	data_out=16'h8006;
17'h619:	data_out=16'h22;
17'h61a:	data_out=16'h75;
17'h61b:	data_out=16'h56;
17'h61c:	data_out=16'h59;
17'h61d:	data_out=16'h69;
17'h61e:	data_out=16'h9;
17'h61f:	data_out=16'h8026;
17'h620:	data_out=16'h54;
17'h621:	data_out=16'h8001;
17'h622:	data_out=16'h8003;
17'h623:	data_out=16'h0;
17'h624:	data_out=16'h1;
17'h625:	data_out=16'h6;
17'h626:	data_out=16'h15;
17'h627:	data_out=16'h60;
17'h628:	data_out=16'h3;
17'h629:	data_out=16'h27;
17'h62a:	data_out=16'h800f;
17'h62b:	data_out=16'h1f;
17'h62c:	data_out=16'h3e;
17'h62d:	data_out=16'h79;
17'h62e:	data_out=16'h800a;
17'h62f:	data_out=16'h52;
17'h630:	data_out=16'ha7;
17'h631:	data_out=16'h65;
17'h632:	data_out=16'hb3;
17'h633:	data_out=16'h7;
17'h634:	data_out=16'h4f;
17'h635:	data_out=16'h6e;
17'h636:	data_out=16'h29;
17'h637:	data_out=16'hd;
17'h638:	data_out=16'h49;
17'h639:	data_out=16'h800e;
17'h63a:	data_out=16'h8044;
17'h63b:	data_out=16'h4f;
17'h63c:	data_out=16'h5f;
17'h63d:	data_out=16'h3c;
17'h63e:	data_out=16'h8006;
17'h63f:	data_out=16'h75;
17'h640:	data_out=16'h12;
17'h641:	data_out=16'h33;
17'h642:	data_out=16'h8c;
17'h643:	data_out=16'h17;
17'h644:	data_out=16'h68;
17'h645:	data_out=16'he;
17'h646:	data_out=16'h3b;
17'h647:	data_out=16'h8032;
17'h648:	data_out=16'h801a;
17'h649:	data_out=16'h9;
17'h64a:	data_out=16'h10;
17'h64b:	data_out=16'h84;
17'h64c:	data_out=16'h3;
17'h64d:	data_out=16'h10;
17'h64e:	data_out=16'h33;
17'h64f:	data_out=16'h9;
17'h650:	data_out=16'h8003;
17'h651:	data_out=16'h2c;
17'h652:	data_out=16'h800a;
17'h653:	data_out=16'h62;
17'h654:	data_out=16'h68;
17'h655:	data_out=16'h30;
17'h656:	data_out=16'h8009;
17'h657:	data_out=16'h8024;
17'h658:	data_out=16'h39;
17'h659:	data_out=16'h1d;
17'h65a:	data_out=16'h46;
17'h65b:	data_out=16'h64;
17'h65c:	data_out=16'h4a;
17'h65d:	data_out=16'h51;
17'h65e:	data_out=16'h71;
17'h65f:	data_out=16'h2;
17'h660:	data_out=16'h29;
17'h661:	data_out=16'h84;
17'h662:	data_out=16'h17;
17'h663:	data_out=16'h13;
17'h664:	data_out=16'h27;
17'h665:	data_out=16'h49;
17'h666:	data_out=16'h19;
17'h667:	data_out=16'h8011;
17'h668:	data_out=16'ha;
17'h669:	data_out=16'h3c;
17'h66a:	data_out=16'h8;
17'h66b:	data_out=16'h5c;
17'h66c:	data_out=16'h5e;
17'h66d:	data_out=16'h3;
17'h66e:	data_out=16'h6;
17'h66f:	data_out=16'h6c;
17'h670:	data_out=16'h8007;
17'h671:	data_out=16'h8046;
17'h672:	data_out=16'h60;
17'h673:	data_out=16'h5c;
17'h674:	data_out=16'ha5;
17'h675:	data_out=16'h8e;
17'h676:	data_out=16'hf;
17'h677:	data_out=16'h23;
17'h678:	data_out=16'hd;
17'h679:	data_out=16'h8005;
17'h67a:	data_out=16'hd;
17'h67b:	data_out=16'h6;
17'h67c:	data_out=16'h8016;
17'h67d:	data_out=16'h8005;
17'h67e:	data_out=16'h8008;
17'h67f:	data_out=16'h8006;
17'h680:	data_out=16'hc9;
17'h681:	data_out=16'h105;
17'h682:	data_out=16'h33;
17'h683:	data_out=16'ha3;
17'h684:	data_out=16'hd1;
17'h685:	data_out=16'he3;
17'h686:	data_out=16'h800b;
17'h687:	data_out=16'h8009;
17'h688:	data_out=16'hb6;
17'h689:	data_out=16'h8039;
17'h68a:	data_out=16'h105;
17'h68b:	data_out=16'h9f;
17'h68c:	data_out=16'h92;
17'h68d:	data_out=16'h42;
17'h68e:	data_out=16'h13;
17'h68f:	data_out=16'h25;
17'h690:	data_out=16'h37;
17'h691:	data_out=16'heb;
17'h692:	data_out=16'h805f;
17'h693:	data_out=16'hcc;
17'h694:	data_out=16'h2c;
17'h695:	data_out=16'h63;
17'h696:	data_out=16'h9c;
17'h697:	data_out=16'h55;
17'h698:	data_out=16'h15;
17'h699:	data_out=16'h6f;
17'h69a:	data_out=16'hfd;
17'h69b:	data_out=16'hd0;
17'h69c:	data_out=16'h10d;
17'h69d:	data_out=16'hfa;
17'h69e:	data_out=16'h36;
17'h69f:	data_out=16'h804e;
17'h6a0:	data_out=16'he4;
17'h6a1:	data_out=16'h11;
17'h6a2:	data_out=16'hc;
17'h6a3:	data_out=16'h8010;
17'h6a4:	data_out=16'h8006;
17'h6a5:	data_out=16'h9;
17'h6a6:	data_out=16'h50;
17'h6a7:	data_out=16'hec;
17'h6a8:	data_out=16'h16;
17'h6a9:	data_out=16'h58;
17'h6aa:	data_out=16'h8016;
17'h6ab:	data_out=16'h76;
17'h6ac:	data_out=16'h8b;
17'h6ad:	data_out=16'hf9;
17'h6ae:	data_out=16'h8003;
17'h6af:	data_out=16'hfb;
17'h6b0:	data_out=16'h178;
17'h6b1:	data_out=16'h113;
17'h6b2:	data_out=16'h196;
17'h6b3:	data_out=16'h13;
17'h6b4:	data_out=16'hc1;
17'h6b5:	data_out=16'h100;
17'h6b6:	data_out=16'h5f;
17'h6b7:	data_out=16'h37;
17'h6b8:	data_out=16'hf7;
17'h6b9:	data_out=16'h24;
17'h6ba:	data_out=16'h808a;
17'h6bb:	data_out=16'hca;
17'h6bc:	data_out=16'hf3;
17'h6bd:	data_out=16'h9e;
17'h6be:	data_out=16'h13;
17'h6bf:	data_out=16'h124;
17'h6c0:	data_out=16'h2f;
17'h6c1:	data_out=16'h96;
17'h6c2:	data_out=16'h11b;
17'h6c3:	data_out=16'h25;
17'h6c4:	data_out=16'hd9;
17'h6c5:	data_out=16'h56;
17'h6c6:	data_out=16'h94;
17'h6c7:	data_out=16'h8077;
17'h6c8:	data_out=16'h8041;
17'h6c9:	data_out=16'h8005;
17'h6ca:	data_out=16'h32;
17'h6cb:	data_out=16'h104;
17'h6cc:	data_out=16'h8008;
17'h6cd:	data_out=16'h1a;
17'h6ce:	data_out=16'h7e;
17'h6cf:	data_out=16'h1a;
17'h6d0:	data_out=16'hd;
17'h6d1:	data_out=16'h93;
17'h6d2:	data_out=16'h1;
17'h6d3:	data_out=16'h11f;
17'h6d4:	data_out=16'hf7;
17'h6d5:	data_out=16'h6b;
17'h6d6:	data_out=16'h8000;
17'h6d7:	data_out=16'h8045;
17'h6d8:	data_out=16'h87;
17'h6d9:	data_out=16'h52;
17'h6da:	data_out=16'ha3;
17'h6db:	data_out=16'h104;
17'h6dc:	data_out=16'hb8;
17'h6dd:	data_out=16'hbc;
17'h6de:	data_out=16'h12f;
17'h6df:	data_out=16'h1c;
17'h6e0:	data_out=16'h69;
17'h6e1:	data_out=16'h140;
17'h6e2:	data_out=16'h42;
17'h6e3:	data_out=16'h39;
17'h6e4:	data_out=16'h69;
17'h6e5:	data_out=16'h96;
17'h6e6:	data_out=16'h56;
17'h6e7:	data_out=16'h8018;
17'h6e8:	data_out=16'ha;
17'h6e9:	data_out=16'ha1;
17'h6ea:	data_out=16'hc;
17'h6eb:	data_out=16'hfa;
17'h6ec:	data_out=16'hfa;
17'h6ed:	data_out=16'h20;
17'h6ee:	data_out=16'h4;
17'h6ef:	data_out=16'h127;
17'h6f0:	data_out=16'h12;
17'h6f1:	data_out=16'h80a4;
17'h6f2:	data_out=16'hfc;
17'h6f3:	data_out=16'hdd;
17'h6f4:	data_out=16'h17b;
17'h6f5:	data_out=16'h154;
17'h6f6:	data_out=16'h2a;
17'h6f7:	data_out=16'h4e;
17'h6f8:	data_out=16'h3b;
17'h6f9:	data_out=16'hc;
17'h6fa:	data_out=16'h33;
17'h6fb:	data_out=16'h12;
17'h6fc:	data_out=16'h802d;
17'h6fd:	data_out=16'h8011;
17'h6fe:	data_out=16'ha;
17'h6ff:	data_out=16'h17;
17'h700:	data_out=16'h2d;
17'h701:	data_out=16'h33;
17'h702:	data_out=16'h10;
17'h703:	data_out=16'h9;
17'h704:	data_out=16'ha;
17'h705:	data_out=16'h21;
17'h706:	data_out=16'h8007;
17'h707:	data_out=16'h5;
17'h708:	data_out=16'h28;
17'h709:	data_out=16'h1b;
17'h70a:	data_out=16'h29;
17'h70b:	data_out=16'h8004;
17'h70c:	data_out=16'h8010;
17'h70d:	data_out=16'h19;
17'h70e:	data_out=16'h8001;
17'h70f:	data_out=16'h3b;
17'h710:	data_out=16'h8000;
17'h711:	data_out=16'h32;
17'h712:	data_out=16'h7;
17'h713:	data_out=16'h32;
17'h714:	data_out=16'h14;
17'h715:	data_out=16'h37;
17'h716:	data_out=16'h44;
17'h717:	data_out=16'h1b;
17'h718:	data_out=16'h1d;
17'h719:	data_out=16'h14;
17'h71a:	data_out=16'h8001;
17'h71b:	data_out=16'h27;
17'h71c:	data_out=16'h41;
17'h71d:	data_out=16'h2f;
17'h71e:	data_out=16'h31;
17'h71f:	data_out=16'h1;
17'h720:	data_out=16'h32;
17'h721:	data_out=16'h7;
17'h722:	data_out=16'h4;
17'h723:	data_out=16'h8007;
17'h724:	data_out=16'h800b;
17'h725:	data_out=16'h3;
17'h726:	data_out=16'h22;
17'h727:	data_out=16'h2a;
17'h728:	data_out=16'h6;
17'h729:	data_out=16'h8001;
17'h72a:	data_out=16'h16;
17'h72b:	data_out=16'h19;
17'h72c:	data_out=16'h11;
17'h72d:	data_out=16'h8013;
17'h72e:	data_out=16'h16;
17'h72f:	data_out=16'h3c;
17'h730:	data_out=16'ha;
17'h731:	data_out=16'h36;
17'h732:	data_out=16'h14;
17'h733:	data_out=16'h14;
17'h734:	data_out=16'h1a;
17'h735:	data_out=16'h8;
17'h736:	data_out=16'h5;
17'h737:	data_out=16'h16;
17'h738:	data_out=16'h59;
17'h739:	data_out=16'h33;
17'h73a:	data_out=16'h1;
17'h73b:	data_out=16'h30;
17'h73c:	data_out=16'h16;
17'h73d:	data_out=16'h36;
17'h73e:	data_out=16'h4;
17'h73f:	data_out=16'h1a;
17'h740:	data_out=16'h8003;
17'h741:	data_out=16'h23;
17'h742:	data_out=16'h8008;
17'h743:	data_out=16'h8005;
17'h744:	data_out=16'he;
17'h745:	data_out=16'h37;
17'h746:	data_out=16'h13;
17'h747:	data_out=16'h8000;
17'h748:	data_out=16'h3;
17'h749:	data_out=16'h8011;
17'h74a:	data_out=16'h8003;
17'h74b:	data_out=16'h801c;
17'h74c:	data_out=16'h8008;
17'h74d:	data_out=16'he;
17'h74e:	data_out=16'h16;
17'h74f:	data_out=16'h8009;
17'h750:	data_out=16'h8002;
17'h751:	data_out=16'h41;
17'h752:	data_out=16'h1;
17'h753:	data_out=16'h3c;
17'h754:	data_out=16'h2b;
17'h755:	data_out=16'h10;
17'h756:	data_out=16'hf;
17'h757:	data_out=16'h4;
17'h758:	data_out=16'h8;
17'h759:	data_out=16'h7;
17'h75a:	data_out=16'h17;
17'h75b:	data_out=16'h2c;
17'h75c:	data_out=16'hc;
17'h75d:	data_out=16'h11;
17'h75e:	data_out=16'h2c;
17'h75f:	data_out=16'h19;
17'h760:	data_out=16'h25;
17'h761:	data_out=16'h39;
17'h762:	data_out=16'h16;
17'h763:	data_out=16'h13;
17'h764:	data_out=16'hd;
17'h765:	data_out=16'hd;
17'h766:	data_out=16'h5;
17'h767:	data_out=16'hf;
17'h768:	data_out=16'h8002;
17'h769:	data_out=16'h1c;
17'h76a:	data_out=16'h1;
17'h76b:	data_out=16'h31;
17'h76c:	data_out=16'h1b;
17'h76d:	data_out=16'h13;
17'h76e:	data_out=16'ha;
17'h76f:	data_out=16'h3e;
17'h770:	data_out=16'hd;
17'h771:	data_out=16'h6;
17'h772:	data_out=16'h2c;
17'h773:	data_out=16'h2b;
17'h774:	data_out=16'hc;
17'h775:	data_out=16'h2e;
17'h776:	data_out=16'h1d;
17'h777:	data_out=16'h800d;
17'h778:	data_out=16'h21;
17'h779:	data_out=16'he;
17'h77a:	data_out=16'h1f;
17'h77b:	data_out=16'hc;
17'h77c:	data_out=16'h8006;
17'h77d:	data_out=16'h3;
17'h77e:	data_out=16'he;
17'h77f:	data_out=16'h9;
17'h780:	data_out=16'h1;
17'h781:	data_out=16'h7;
17'h782:	data_out=16'h4;
17'h783:	data_out=16'h6;
17'h784:	data_out=16'h3;
17'h785:	data_out=16'h8006;
17'h786:	data_out=16'h5;
17'h787:	data_out=16'h5;
17'h788:	data_out=16'h6;
17'h789:	data_out=16'ha;
17'h78a:	data_out=16'h8006;
17'h78b:	data_out=16'h8005;
17'h78c:	data_out=16'h8005;
17'h78d:	data_out=16'h8;
17'h78e:	data_out=16'h8007;
17'h78f:	data_out=16'h8003;
17'h790:	data_out=16'h8003;
17'h791:	data_out=16'h5;
17'h792:	data_out=16'h8;
17'h793:	data_out=16'h3;
17'h794:	data_out=16'h9;
17'h795:	data_out=16'h2;
17'h796:	data_out=16'hb;
17'h797:	data_out=16'h4;
17'h798:	data_out=16'h5;
17'h799:	data_out=16'h6;
17'h79a:	data_out=16'h8001;
17'h79b:	data_out=16'h8007;
17'h79c:	data_out=16'h8003;
17'h79d:	data_out=16'h2;
17'h79e:	data_out=16'h8003;
17'h79f:	data_out=16'h2;
17'h7a0:	data_out=16'h8003;
17'h7a1:	data_out=16'h8;
17'h7a2:	data_out=16'h8002;
17'h7a3:	data_out=16'h7;
17'h7a4:	data_out=16'h8008;
17'h7a5:	data_out=16'h8007;
17'h7a6:	data_out=16'h3;
17'h7a7:	data_out=16'h7;
17'h7a8:	data_out=16'h8007;
17'h7a9:	data_out=16'h4;
17'h7aa:	data_out=16'h8009;
17'h7ab:	data_out=16'h8001;
17'h7ac:	data_out=16'h2;
17'h7ad:	data_out=16'h8008;
17'h7ae:	data_out=16'h2;
17'h7af:	data_out=16'h9;
17'h7b0:	data_out=16'h6;
17'h7b1:	data_out=16'h3;
17'h7b2:	data_out=16'h8001;
17'h7b3:	data_out=16'h5;
17'h7b4:	data_out=16'h8008;
17'h7b5:	data_out=16'h8002;
17'h7b6:	data_out=16'h8001;
17'h7b7:	data_out=16'h5;
17'h7b8:	data_out=16'h8003;
17'h7b9:	data_out=16'h9;
17'h7ba:	data_out=16'h4;
17'h7bb:	data_out=16'h8003;
17'h7bc:	data_out=16'h8001;
17'h7bd:	data_out=16'h8007;
17'h7be:	data_out=16'h7;
17'h7bf:	data_out=16'h3;
17'h7c0:	data_out=16'h9;
17'h7c1:	data_out=16'h8003;
17'h7c2:	data_out=16'h8001;
17'h7c3:	data_out=16'h8009;
17'h7c4:	data_out=16'h8002;
17'h7c5:	data_out=16'h8005;
17'h7c6:	data_out=16'h7;
17'h7c7:	data_out=16'h8001;
17'h7c8:	data_out=16'h5;
17'h7c9:	data_out=16'h6;
17'h7ca:	data_out=16'h7;
17'h7cb:	data_out=16'h8003;
17'h7cc:	data_out=16'h8;
17'h7cd:	data_out=16'h8001;
17'h7ce:	data_out=16'h8003;
17'h7cf:	data_out=16'h4;
17'h7d0:	data_out=16'h9;
17'h7d1:	data_out=16'h6;
17'h7d2:	data_out=16'h8001;
17'h7d3:	data_out=16'h8006;
17'h7d4:	data_out=16'h8007;
17'h7d5:	data_out=16'h7;
17'h7d6:	data_out=16'h5;
17'h7d7:	data_out=16'h8006;
17'h7d8:	data_out=16'h5;
17'h7d9:	data_out=16'h0;
17'h7da:	data_out=16'h8001;
17'h7db:	data_out=16'h8006;
17'h7dc:	data_out=16'h1;
17'h7dd:	data_out=16'h8003;
17'h7de:	data_out=16'h5;
17'h7df:	data_out=16'h1;
17'h7e0:	data_out=16'h2;
17'h7e1:	data_out=16'h8004;
17'h7e2:	data_out=16'h1;
17'h7e3:	data_out=16'h8;
17'h7e4:	data_out=16'h8004;
17'h7e5:	data_out=16'h8003;
17'h7e6:	data_out=16'h8002;
17'h7e7:	data_out=16'h8009;
17'h7e8:	data_out=16'h8005;
17'h7e9:	data_out=16'h8003;
17'h7ea:	data_out=16'h8002;
17'h7eb:	data_out=16'h8005;
17'h7ec:	data_out=16'h5;
17'h7ed:	data_out=16'h4;
17'h7ee:	data_out=16'h6;
17'h7ef:	data_out=16'h6;
17'h7f0:	data_out=16'h8003;
17'h7f1:	data_out=16'h8004;
17'h7f2:	data_out=16'h6;
17'h7f3:	data_out=16'h8001;
17'h7f4:	data_out=16'h8006;
17'h7f5:	data_out=16'h2;
17'h7f6:	data_out=16'h1;
17'h7f7:	data_out=16'h6;
17'h7f8:	data_out=16'ha;
17'h7f9:	data_out=16'h9;
17'h7fa:	data_out=16'h9;
17'h7fb:	data_out=16'h1;
17'h7fc:	data_out=16'h8005;
17'h7fd:	data_out=16'h2;
17'h7fe:	data_out=16'ha;
17'h7ff:	data_out=16'h6;
17'h800:	data_out=16'h4;
17'h801:	data_out=16'h0;
17'h802:	data_out=16'h4;
17'h803:	data_out=16'h8;
17'h804:	data_out=16'h7;
17'h805:	data_out=16'h8008;
17'h806:	data_out=16'h9;
17'h807:	data_out=16'h8008;
17'h808:	data_out=16'h8003;
17'h809:	data_out=16'h8003;
17'h80a:	data_out=16'h8006;
17'h80b:	data_out=16'h8008;
17'h80c:	data_out=16'h8009;
17'h80d:	data_out=16'h8009;
17'h80e:	data_out=16'h5;
17'h80f:	data_out=16'h8003;
17'h810:	data_out=16'h8004;
17'h811:	data_out=16'h0;
17'h812:	data_out=16'h3;
17'h813:	data_out=16'h8001;
17'h814:	data_out=16'h8009;
17'h815:	data_out=16'h8005;
17'h816:	data_out=16'h8004;
17'h817:	data_out=16'h8009;
17'h818:	data_out=16'h8007;
17'h819:	data_out=16'h8005;
17'h81a:	data_out=16'h0;
17'h81b:	data_out=16'h8002;
17'h81c:	data_out=16'h6;
17'h81d:	data_out=16'h0;
17'h81e:	data_out=16'h8006;
17'h81f:	data_out=16'h1;
17'h820:	data_out=16'h8009;
17'h821:	data_out=16'h6;
17'h822:	data_out=16'h0;
17'h823:	data_out=16'h7;
17'h824:	data_out=16'h8;
17'h825:	data_out=16'h8000;
17'h826:	data_out=16'h8;
17'h827:	data_out=16'h8004;
17'h828:	data_out=16'h6;
17'h829:	data_out=16'h8007;
17'h82a:	data_out=16'h8003;
17'h82b:	data_out=16'h7;
17'h82c:	data_out=16'h8007;
17'h82d:	data_out=16'h8007;
17'h82e:	data_out=16'h8006;
17'h82f:	data_out=16'h8001;
17'h830:	data_out=16'h3;
17'h831:	data_out=16'h7;
17'h832:	data_out=16'h7;
17'h833:	data_out=16'h3;
17'h834:	data_out=16'h8008;
17'h835:	data_out=16'h8006;
17'h836:	data_out=16'h3;
17'h837:	data_out=16'h8005;
17'h838:	data_out=16'h8002;
17'h839:	data_out=16'h8006;
17'h83a:	data_out=16'h2;
17'h83b:	data_out=16'h8005;
17'h83c:	data_out=16'h4;
17'h83d:	data_out=16'h5;
17'h83e:	data_out=16'h5;
17'h83f:	data_out=16'h4;
17'h840:	data_out=16'h2;
17'h841:	data_out=16'h8004;
17'h842:	data_out=16'h2;
17'h843:	data_out=16'h1;
17'h844:	data_out=16'h5;
17'h845:	data_out=16'h1;
17'h846:	data_out=16'h6;
17'h847:	data_out=16'h2;
17'h848:	data_out=16'h3;
17'h849:	data_out=16'h8006;
17'h84a:	data_out=16'h8000;
17'h84b:	data_out=16'h5;
17'h84c:	data_out=16'h8004;
17'h84d:	data_out=16'h3;
17'h84e:	data_out=16'h8005;
17'h84f:	data_out=16'h8;
17'h850:	data_out=16'h1;
17'h851:	data_out=16'h8008;
17'h852:	data_out=16'h2;
17'h853:	data_out=16'h2;
17'h854:	data_out=16'h8005;
17'h855:	data_out=16'h8005;
17'h856:	data_out=16'h7;
17'h857:	data_out=16'h2;
17'h858:	data_out=16'h8001;
17'h859:	data_out=16'h8001;
17'h85a:	data_out=16'h6;
17'h85b:	data_out=16'h8007;
17'h85c:	data_out=16'h8005;
17'h85d:	data_out=16'h1;
17'h85e:	data_out=16'h7;
17'h85f:	data_out=16'h6;
17'h860:	data_out=16'h7;
17'h861:	data_out=16'h8000;
17'h862:	data_out=16'h8003;
17'h863:	data_out=16'h3;
17'h864:	data_out=16'h8009;
17'h865:	data_out=16'h8006;
17'h866:	data_out=16'h8004;
17'h867:	data_out=16'h4;
17'h868:	data_out=16'h8003;
17'h869:	data_out=16'h5;
17'h86a:	data_out=16'h8000;
17'h86b:	data_out=16'h2;
17'h86c:	data_out=16'h8001;
17'h86d:	data_out=16'h3;
17'h86e:	data_out=16'h1;
17'h86f:	data_out=16'h8009;
17'h870:	data_out=16'h4;
17'h871:	data_out=16'h8006;
17'h872:	data_out=16'h3;
17'h873:	data_out=16'h8;
17'h874:	data_out=16'h8001;
17'h875:	data_out=16'h0;
17'h876:	data_out=16'h1;
17'h877:	data_out=16'h7;
17'h878:	data_out=16'h9;
17'h879:	data_out=16'h8002;
17'h87a:	data_out=16'h9;
17'h87b:	data_out=16'h8006;
17'h87c:	data_out=16'h8;
17'h87d:	data_out=16'h6;
17'h87e:	data_out=16'h9;
17'h87f:	data_out=16'h6;
17'h880:	data_out=16'h8003;
17'h881:	data_out=16'h8003;
17'h882:	data_out=16'h8001;
17'h883:	data_out=16'h8003;
17'h884:	data_out=16'h8000;
17'h885:	data_out=16'h5;
17'h886:	data_out=16'h8008;
17'h887:	data_out=16'h6;
17'h888:	data_out=16'h1;
17'h889:	data_out=16'h0;
17'h88a:	data_out=16'h8001;
17'h88b:	data_out=16'h8009;
17'h88c:	data_out=16'h8005;
17'h88d:	data_out=16'h8009;
17'h88e:	data_out=16'h8009;
17'h88f:	data_out=16'h8;
17'h890:	data_out=16'h8006;
17'h891:	data_out=16'h3;
17'h892:	data_out=16'h7;
17'h893:	data_out=16'h2;
17'h894:	data_out=16'h8005;
17'h895:	data_out=16'h8001;
17'h896:	data_out=16'h8001;
17'h897:	data_out=16'h8006;
17'h898:	data_out=16'h6;
17'h899:	data_out=16'h8001;
17'h89a:	data_out=16'h8003;
17'h89b:	data_out=16'h5;
17'h89c:	data_out=16'h8004;
17'h89d:	data_out=16'h8003;
17'h89e:	data_out=16'h1;
17'h89f:	data_out=16'h2;
17'h8a0:	data_out=16'h3;
17'h8a1:	data_out=16'h8008;
17'h8a2:	data_out=16'h9;
17'h8a3:	data_out=16'h8006;
17'h8a4:	data_out=16'h6;
17'h8a5:	data_out=16'h8009;
17'h8a6:	data_out=16'h8;
17'h8a7:	data_out=16'h8003;
17'h8a8:	data_out=16'h1;
17'h8a9:	data_out=16'h8002;
17'h8aa:	data_out=16'h8003;
17'h8ab:	data_out=16'h5;
17'h8ac:	data_out=16'h8001;
17'h8ad:	data_out=16'h8002;
17'h8ae:	data_out=16'h4;
17'h8af:	data_out=16'h2;
17'h8b0:	data_out=16'h8008;
17'h8b1:	data_out=16'h2;
17'h8b2:	data_out=16'h8005;
17'h8b3:	data_out=16'h8004;
17'h8b4:	data_out=16'h8008;
17'h8b5:	data_out=16'h3;
17'h8b6:	data_out=16'h8001;
17'h8b7:	data_out=16'h7;
17'h8b8:	data_out=16'h8007;
17'h8b9:	data_out=16'h5;
17'h8ba:	data_out=16'h2;
17'h8bb:	data_out=16'h8001;
17'h8bc:	data_out=16'h8007;
17'h8bd:	data_out=16'h8006;
17'h8be:	data_out=16'h8008;
17'h8bf:	data_out=16'h5;
17'h8c0:	data_out=16'h8005;
17'h8c1:	data_out=16'h8009;
17'h8c2:	data_out=16'h8;
17'h8c3:	data_out=16'h8009;
17'h8c4:	data_out=16'h8008;
17'h8c5:	data_out=16'h7;
17'h8c6:	data_out=16'h8002;
17'h8c7:	data_out=16'h2;
17'h8c8:	data_out=16'h8004;
17'h8c9:	data_out=16'h4;
17'h8ca:	data_out=16'h8002;
17'h8cb:	data_out=16'h4;
17'h8cc:	data_out=16'h8007;
17'h8cd:	data_out=16'h8008;
17'h8ce:	data_out=16'h8003;
17'h8cf:	data_out=16'h8006;
17'h8d0:	data_out=16'h3;
17'h8d1:	data_out=16'h1;
17'h8d2:	data_out=16'h8001;
17'h8d3:	data_out=16'h4;
17'h8d4:	data_out=16'h8005;
17'h8d5:	data_out=16'h8;
17'h8d6:	data_out=16'h1;
17'h8d7:	data_out=16'h8003;
17'h8d8:	data_out=16'h4;
17'h8d9:	data_out=16'h8006;
17'h8da:	data_out=16'h5;
17'h8db:	data_out=16'h6;
17'h8dc:	data_out=16'h8003;
17'h8dd:	data_out=16'h6;
17'h8de:	data_out=16'h3;
17'h8df:	data_out=16'h2;
17'h8e0:	data_out=16'h7;
17'h8e1:	data_out=16'h2;
17'h8e2:	data_out=16'h2;
17'h8e3:	data_out=16'h8;
17'h8e4:	data_out=16'h8000;
17'h8e5:	data_out=16'h9;
17'h8e6:	data_out=16'h1;
17'h8e7:	data_out=16'h5;
17'h8e8:	data_out=16'h4;
17'h8e9:	data_out=16'h7;
17'h8ea:	data_out=16'h1;
17'h8eb:	data_out=16'h7;
17'h8ec:	data_out=16'h9;
17'h8ed:	data_out=16'h7;
17'h8ee:	data_out=16'h8008;
17'h8ef:	data_out=16'h2;
17'h8f0:	data_out=16'h8002;
17'h8f1:	data_out=16'h0;
17'h8f2:	data_out=16'h8003;
17'h8f3:	data_out=16'h3;
17'h8f4:	data_out=16'h8001;
17'h8f5:	data_out=16'h7;
17'h8f6:	data_out=16'h9;
17'h8f7:	data_out=16'h8006;
17'h8f8:	data_out=16'h8009;
17'h8f9:	data_out=16'h5;
17'h8fa:	data_out=16'h8009;
17'h8fb:	data_out=16'h8002;
17'h8fc:	data_out=16'h2;
17'h8fd:	data_out=16'h3;
17'h8fe:	data_out=16'h9;
17'h8ff:	data_out=16'h8001;
17'h900:	data_out=16'h8005;
17'h901:	data_out=16'h2;
17'h902:	data_out=16'h8002;
17'h903:	data_out=16'h4;
17'h904:	data_out=16'h2;
17'h905:	data_out=16'h8;
17'h906:	data_out=16'h1;
17'h907:	data_out=16'h8003;
17'h908:	data_out=16'h6;
17'h909:	data_out=16'h8008;
17'h90a:	data_out=16'h8006;
17'h90b:	data_out=16'h5;
17'h90c:	data_out=16'h8;
17'h90d:	data_out=16'h8005;
17'h90e:	data_out=16'h8002;
17'h90f:	data_out=16'h8003;
17'h910:	data_out=16'h5;
17'h911:	data_out=16'h4;
17'h912:	data_out=16'h9;
17'h913:	data_out=16'h8005;
17'h914:	data_out=16'h1;
17'h915:	data_out=16'h9;
17'h916:	data_out=16'h8003;
17'h917:	data_out=16'h2;
17'h918:	data_out=16'h5;
17'h919:	data_out=16'h8003;
17'h91a:	data_out=16'h9;
17'h91b:	data_out=16'h8002;
17'h91c:	data_out=16'h8009;
17'h91d:	data_out=16'h9;
17'h91e:	data_out=16'h6;
17'h91f:	data_out=16'h8004;
17'h920:	data_out=16'h1;
17'h921:	data_out=16'h8005;
17'h922:	data_out=16'h9;
17'h923:	data_out=16'h8006;
17'h924:	data_out=16'h8006;
17'h925:	data_out=16'h0;
17'h926:	data_out=16'h8000;
17'h927:	data_out=16'h9;
17'h928:	data_out=16'h1;
17'h929:	data_out=16'h3;
17'h92a:	data_out=16'h5;
17'h92b:	data_out=16'h0;
17'h92c:	data_out=16'h7;
17'h92d:	data_out=16'h8006;
17'h92e:	data_out=16'h6;
17'h92f:	data_out=16'h3;
17'h930:	data_out=16'h7;
17'h931:	data_out=16'h6;
17'h932:	data_out=16'h6;
17'h933:	data_out=16'h8001;
17'h934:	data_out=16'h6;
17'h935:	data_out=16'h8005;
17'h936:	data_out=16'h8008;
17'h937:	data_out=16'h1;
17'h938:	data_out=16'h1;
17'h939:	data_out=16'h8008;
17'h93a:	data_out=16'h8;
17'h93b:	data_out=16'h2;
17'h93c:	data_out=16'h8009;
17'h93d:	data_out=16'h5;
17'h93e:	data_out=16'h6;
17'h93f:	data_out=16'h2;
17'h940:	data_out=16'h8009;
17'h941:	data_out=16'h6;
17'h942:	data_out=16'h4;
17'h943:	data_out=16'h8006;
17'h944:	data_out=16'h8002;
17'h945:	data_out=16'h8005;
17'h946:	data_out=16'h8007;
17'h947:	data_out=16'h8;
17'h948:	data_out=16'h7;
17'h949:	data_out=16'h7;
17'h94a:	data_out=16'h8001;
17'h94b:	data_out=16'h5;
17'h94c:	data_out=16'h8008;
17'h94d:	data_out=16'h8004;
17'h94e:	data_out=16'h8002;
17'h94f:	data_out=16'h8;
17'h950:	data_out=16'h8007;
17'h951:	data_out=16'h8004;
17'h952:	data_out=16'h8002;
17'h953:	data_out=16'h8;
17'h954:	data_out=16'h8000;
17'h955:	data_out=16'h8001;
17'h956:	data_out=16'h0;
17'h957:	data_out=16'h8008;
17'h958:	data_out=16'h8000;
17'h959:	data_out=16'h8000;
17'h95a:	data_out=16'h2;
17'h95b:	data_out=16'h0;
17'h95c:	data_out=16'h8004;
17'h95d:	data_out=16'h8000;
17'h95e:	data_out=16'h8007;
17'h95f:	data_out=16'h8004;
17'h960:	data_out=16'h8003;
17'h961:	data_out=16'h6;
17'h962:	data_out=16'h8001;
17'h963:	data_out=16'h4;
17'h964:	data_out=16'h8008;
17'h965:	data_out=16'h2;
17'h966:	data_out=16'h3;
17'h967:	data_out=16'h8;
17'h968:	data_out=16'h8001;
17'h969:	data_out=16'h8008;
17'h96a:	data_out=16'h3;
17'h96b:	data_out=16'h0;
17'h96c:	data_out=16'h8002;
17'h96d:	data_out=16'h8007;
17'h96e:	data_out=16'h8001;
17'h96f:	data_out=16'h0;
17'h970:	data_out=16'h8003;
17'h971:	data_out=16'h6;
17'h972:	data_out=16'h8001;
17'h973:	data_out=16'h6;
17'h974:	data_out=16'h8004;
17'h975:	data_out=16'h9;
17'h976:	data_out=16'h7;
17'h977:	data_out=16'h5;
17'h978:	data_out=16'h8001;
17'h979:	data_out=16'h0;
17'h97a:	data_out=16'h8004;
17'h97b:	data_out=16'h4;
17'h97c:	data_out=16'h8009;
17'h97d:	data_out=16'h8002;
17'h97e:	data_out=16'h8009;
17'h97f:	data_out=16'h8003;
17'h980:	data_out=16'h8005;
17'h981:	data_out=16'h8000;
17'h982:	data_out=16'h8009;
17'h983:	data_out=16'h8004;
17'h984:	data_out=16'h8008;
17'h985:	data_out=16'h3;
17'h986:	data_out=16'h8006;
17'h987:	data_out=16'h0;
17'h988:	data_out=16'h5;
17'h989:	data_out=16'h6;
17'h98a:	data_out=16'h8008;
17'h98b:	data_out=16'h8007;
17'h98c:	data_out=16'h8;
17'h98d:	data_out=16'h8000;
17'h98e:	data_out=16'h3;
17'h98f:	data_out=16'h8004;
17'h990:	data_out=16'h8004;
17'h991:	data_out=16'h8007;
17'h992:	data_out=16'h8007;
17'h993:	data_out=16'h1;
17'h994:	data_out=16'h8008;
17'h995:	data_out=16'h8009;
17'h996:	data_out=16'h8004;
17'h997:	data_out=16'h1;
17'h998:	data_out=16'h1;
17'h999:	data_out=16'h1;
17'h99a:	data_out=16'h8004;
17'h99b:	data_out=16'h1;
17'h99c:	data_out=16'h8;
17'h99d:	data_out=16'h8004;
17'h99e:	data_out=16'h7;
17'h99f:	data_out=16'h8006;
17'h9a0:	data_out=16'h5;
17'h9a1:	data_out=16'h7;
17'h9a2:	data_out=16'h8002;
17'h9a3:	data_out=16'h6;
17'h9a4:	data_out=16'h1;
17'h9a5:	data_out=16'h1;
17'h9a6:	data_out=16'h8003;
17'h9a7:	data_out=16'h8004;
17'h9a8:	data_out=16'h8001;
17'h9a9:	data_out=16'h8002;
17'h9aa:	data_out=16'h8001;
17'h9ab:	data_out=16'h8002;
17'h9ac:	data_out=16'h7;
17'h9ad:	data_out=16'h8008;
17'h9ae:	data_out=16'h3;
17'h9af:	data_out=16'h8006;
17'h9b0:	data_out=16'h8006;
17'h9b1:	data_out=16'h6;
17'h9b2:	data_out=16'h4;
17'h9b3:	data_out=16'h8005;
17'h9b4:	data_out=16'h6;
17'h9b5:	data_out=16'h9;
17'h9b6:	data_out=16'h5;
17'h9b7:	data_out=16'h8003;
17'h9b8:	data_out=16'h1;
17'h9b9:	data_out=16'h8008;
17'h9ba:	data_out=16'h7;
17'h9bb:	data_out=16'h8000;
17'h9bc:	data_out=16'h8003;
17'h9bd:	data_out=16'h5;
17'h9be:	data_out=16'h3;
17'h9bf:	data_out=16'h8008;
17'h9c0:	data_out=16'h3;
17'h9c1:	data_out=16'h8008;
17'h9c2:	data_out=16'h7;
17'h9c3:	data_out=16'h8006;
17'h9c4:	data_out=16'h2;
17'h9c5:	data_out=16'h8005;
17'h9c6:	data_out=16'h8000;
17'h9c7:	data_out=16'h8008;
17'h9c8:	data_out=16'h2;
17'h9c9:	data_out=16'h8;
17'h9ca:	data_out=16'h8002;
17'h9cb:	data_out=16'h8000;
17'h9cc:	data_out=16'h8009;
17'h9cd:	data_out=16'h8008;
17'h9ce:	data_out=16'h2;
17'h9cf:	data_out=16'h8006;
17'h9d0:	data_out=16'h7;
17'h9d1:	data_out=16'h8003;
17'h9d2:	data_out=16'h8001;
17'h9d3:	data_out=16'h4;
17'h9d4:	data_out=16'h8003;
17'h9d5:	data_out=16'h8005;
17'h9d6:	data_out=16'h8008;
17'h9d7:	data_out=16'h7;
17'h9d8:	data_out=16'h8005;
17'h9d9:	data_out=16'h8;
17'h9da:	data_out=16'h8002;
17'h9db:	data_out=16'h1;
17'h9dc:	data_out=16'h4;
17'h9dd:	data_out=16'h8009;
17'h9de:	data_out=16'h3;
17'h9df:	data_out=16'h8002;
17'h9e0:	data_out=16'h8008;
17'h9e1:	data_out=16'h1;
17'h9e2:	data_out=16'h1;
17'h9e3:	data_out=16'h3;
17'h9e4:	data_out=16'h6;
17'h9e5:	data_out=16'h8008;
17'h9e6:	data_out=16'h4;
17'h9e7:	data_out=16'h8001;
17'h9e8:	data_out=16'h9;
17'h9e9:	data_out=16'h8007;
17'h9ea:	data_out=16'h8;
17'h9eb:	data_out=16'h9;
17'h9ec:	data_out=16'h8006;
17'h9ed:	data_out=16'h1;
17'h9ee:	data_out=16'h8006;
17'h9ef:	data_out=16'h8008;
17'h9f0:	data_out=16'h7;
17'h9f1:	data_out=16'h2;
17'h9f2:	data_out=16'h5;
17'h9f3:	data_out=16'h8006;
17'h9f4:	data_out=16'h5;
17'h9f5:	data_out=16'h6;
17'h9f6:	data_out=16'h8008;
17'h9f7:	data_out=16'h8008;
17'h9f8:	data_out=16'h6;
17'h9f9:	data_out=16'h8001;
17'h9fa:	data_out=16'h2;
17'h9fb:	data_out=16'h1;
17'h9fc:	data_out=16'h8001;
17'h9fd:	data_out=16'h8004;
17'h9fe:	data_out=16'h7;
17'h9ff:	data_out=16'h8000;
17'ha00:	data_out=16'h7;
17'ha01:	data_out=16'h8001;
17'ha02:	data_out=16'h8006;
17'ha03:	data_out=16'h3;
17'ha04:	data_out=16'h0;
17'ha05:	data_out=16'h6;
17'ha06:	data_out=16'h8007;
17'ha07:	data_out=16'h8000;
17'ha08:	data_out=16'h8;
17'ha09:	data_out=16'h8008;
17'ha0a:	data_out=16'h8000;
17'ha0b:	data_out=16'h8007;
17'ha0c:	data_out=16'h2;
17'ha0d:	data_out=16'h3;
17'ha0e:	data_out=16'h8005;
17'ha0f:	data_out=16'h8000;
17'ha10:	data_out=16'h8005;
17'ha11:	data_out=16'h9;
17'ha12:	data_out=16'h3;
17'ha13:	data_out=16'h8008;
17'ha14:	data_out=16'h6;
17'ha15:	data_out=16'h5;
17'ha16:	data_out=16'h8008;
17'ha17:	data_out=16'h3;
17'ha18:	data_out=16'h8006;
17'ha19:	data_out=16'h4;
17'ha1a:	data_out=16'h8006;
17'ha1b:	data_out=16'h2;
17'ha1c:	data_out=16'h9;
17'ha1d:	data_out=16'h8008;
17'ha1e:	data_out=16'h8007;
17'ha1f:	data_out=16'h6;
17'ha20:	data_out=16'h0;
17'ha21:	data_out=16'h8004;
17'ha22:	data_out=16'h1;
17'ha23:	data_out=16'h8009;
17'ha24:	data_out=16'h8007;
17'ha25:	data_out=16'h3;
17'ha26:	data_out=16'h1;
17'ha27:	data_out=16'h8008;
17'ha28:	data_out=16'h4;
17'ha29:	data_out=16'h8009;
17'ha2a:	data_out=16'h8005;
17'ha2b:	data_out=16'h8004;
17'ha2c:	data_out=16'h3;
17'ha2d:	data_out=16'h8002;
17'ha2e:	data_out=16'h5;
17'ha2f:	data_out=16'h8;
17'ha30:	data_out=16'h8002;
17'ha31:	data_out=16'h8001;
17'ha32:	data_out=16'h8;
17'ha33:	data_out=16'h8005;
17'ha34:	data_out=16'h8006;
17'ha35:	data_out=16'h8009;
17'ha36:	data_out=16'h7;
17'ha37:	data_out=16'h8002;
17'ha38:	data_out=16'h4;
17'ha39:	data_out=16'h8009;
17'ha3a:	data_out=16'h8009;
17'ha3b:	data_out=16'h4;
17'ha3c:	data_out=16'h8007;
17'ha3d:	data_out=16'h8007;
17'ha3e:	data_out=16'h1;
17'ha3f:	data_out=16'h2;
17'ha40:	data_out=16'h8002;
17'ha41:	data_out=16'h8007;
17'ha42:	data_out=16'h3;
17'ha43:	data_out=16'h0;
17'ha44:	data_out=16'h4;
17'ha45:	data_out=16'h8006;
17'ha46:	data_out=16'h2;
17'ha47:	data_out=16'h8001;
17'ha48:	data_out=16'h8005;
17'ha49:	data_out=16'h5;
17'ha4a:	data_out=16'h4;
17'ha4b:	data_out=16'h7;
17'ha4c:	data_out=16'h8005;
17'ha4d:	data_out=16'h0;
17'ha4e:	data_out=16'h5;
17'ha4f:	data_out=16'h2;
17'ha50:	data_out=16'h8;
17'ha51:	data_out=16'h5;
17'ha52:	data_out=16'h6;
17'ha53:	data_out=16'h8006;
17'ha54:	data_out=16'h5;
17'ha55:	data_out=16'h3;
17'ha56:	data_out=16'h1;
17'ha57:	data_out=16'h0;
17'ha58:	data_out=16'h4;
17'ha59:	data_out=16'h1;
17'ha5a:	data_out=16'h8005;
17'ha5b:	data_out=16'h6;
17'ha5c:	data_out=16'h3;
17'ha5d:	data_out=16'h5;
17'ha5e:	data_out=16'h8001;
17'ha5f:	data_out=16'h8008;
17'ha60:	data_out=16'h7;
17'ha61:	data_out=16'h8008;
17'ha62:	data_out=16'h2;
17'ha63:	data_out=16'h3;
17'ha64:	data_out=16'h8004;
17'ha65:	data_out=16'h8006;
17'ha66:	data_out=16'h8008;
17'ha67:	data_out=16'h8001;
17'ha68:	data_out=16'h9;
17'ha69:	data_out=16'h6;
17'ha6a:	data_out=16'h8003;
17'ha6b:	data_out=16'h8006;
17'ha6c:	data_out=16'h8003;
17'ha6d:	data_out=16'h8007;
17'ha6e:	data_out=16'h5;
17'ha6f:	data_out=16'h8004;
17'ha70:	data_out=16'h7;
17'ha71:	data_out=16'h2;
17'ha72:	data_out=16'h8001;
17'ha73:	data_out=16'h3;
17'ha74:	data_out=16'h8004;
17'ha75:	data_out=16'h9;
17'ha76:	data_out=16'h8006;
17'ha77:	data_out=16'h9;
17'ha78:	data_out=16'h0;
17'ha79:	data_out=16'h8002;
17'ha7a:	data_out=16'h5;
17'ha7b:	data_out=16'h8006;
17'ha7c:	data_out=16'h8005;
17'ha7d:	data_out=16'h8005;
17'ha7e:	data_out=16'h8004;
17'ha7f:	data_out=16'h8007;
17'ha80:	data_out=16'h8004;
17'ha81:	data_out=16'h7;
17'ha82:	data_out=16'h5;
17'ha83:	data_out=16'h1;
17'ha84:	data_out=16'h8008;
17'ha85:	data_out=16'h6;
17'ha86:	data_out=16'h9;
17'ha87:	data_out=16'h8009;
17'ha88:	data_out=16'h3;
17'ha89:	data_out=16'h8003;
17'ha8a:	data_out=16'h8005;
17'ha8b:	data_out=16'h9;
17'ha8c:	data_out=16'h8001;
17'ha8d:	data_out=16'h9;
17'ha8e:	data_out=16'h8004;
17'ha8f:	data_out=16'h8003;
17'ha90:	data_out=16'h1;
17'ha91:	data_out=16'h4;
17'ha92:	data_out=16'h8009;
17'ha93:	data_out=16'h6;
17'ha94:	data_out=16'h3;
17'ha95:	data_out=16'h8005;
17'ha96:	data_out=16'h6;
17'ha97:	data_out=16'h8006;
17'ha98:	data_out=16'h2;
17'ha99:	data_out=16'h2;
17'ha9a:	data_out=16'h8002;
17'ha9b:	data_out=16'h6;
17'ha9c:	data_out=16'h6;
17'ha9d:	data_out=16'h3;
17'ha9e:	data_out=16'h8;
17'ha9f:	data_out=16'h8008;
17'haa0:	data_out=16'h0;
17'haa1:	data_out=16'h4;
17'haa2:	data_out=16'h2;
17'haa3:	data_out=16'h1;
17'haa4:	data_out=16'h1;
17'haa5:	data_out=16'h2;
17'haa6:	data_out=16'h2;
17'haa7:	data_out=16'h8006;
17'haa8:	data_out=16'h8;
17'haa9:	data_out=16'h5;
17'haaa:	data_out=16'h8006;
17'haab:	data_out=16'h8002;
17'haac:	data_out=16'h5;
17'haad:	data_out=16'h8001;
17'haae:	data_out=16'h4;
17'haaf:	data_out=16'h8003;
17'hab0:	data_out=16'h8006;
17'hab1:	data_out=16'h5;
17'hab2:	data_out=16'h8006;
17'hab3:	data_out=16'h6;
17'hab4:	data_out=16'h8;
17'hab5:	data_out=16'h8009;
17'hab6:	data_out=16'h8008;
17'hab7:	data_out=16'h1;
17'hab8:	data_out=16'h2;
17'hab9:	data_out=16'h8001;
17'haba:	data_out=16'h8002;
17'habb:	data_out=16'h8001;
17'habc:	data_out=16'h8008;
17'habd:	data_out=16'h8003;
17'habe:	data_out=16'h0;
17'habf:	data_out=16'h1;
17'hac0:	data_out=16'h8008;
17'hac1:	data_out=16'h8007;
17'hac2:	data_out=16'h8007;
17'hac3:	data_out=16'h2;
17'hac4:	data_out=16'h4;
17'hac5:	data_out=16'h4;
17'hac6:	data_out=16'h5;
17'hac7:	data_out=16'h3;
17'hac8:	data_out=16'h8000;
17'hac9:	data_out=16'h9;
17'haca:	data_out=16'h8008;
17'hacb:	data_out=16'h8004;
17'hacc:	data_out=16'h8001;
17'hacd:	data_out=16'h6;
17'hace:	data_out=16'h2;
17'hacf:	data_out=16'h2;
17'had0:	data_out=16'h1;
17'had1:	data_out=16'h6;
17'had2:	data_out=16'h8001;
17'had3:	data_out=16'h0;
17'had4:	data_out=16'h6;
17'had5:	data_out=16'h0;
17'had6:	data_out=16'h8007;
17'had7:	data_out=16'h8001;
17'had8:	data_out=16'h8;
17'had9:	data_out=16'h0;
17'hada:	data_out=16'h6;
17'hadb:	data_out=16'h9;
17'hadc:	data_out=16'h7;
17'hadd:	data_out=16'h8003;
17'hade:	data_out=16'h1;
17'hadf:	data_out=16'h8;
17'hae0:	data_out=16'h8000;
17'hae1:	data_out=16'h3;
17'hae2:	data_out=16'h1;
17'hae3:	data_out=16'h8005;
17'hae4:	data_out=16'h8002;
17'hae5:	data_out=16'h8003;
17'hae6:	data_out=16'h7;
17'hae7:	data_out=16'h7;
17'hae8:	data_out=16'h8004;
17'hae9:	data_out=16'h8;
17'haea:	data_out=16'h8006;
17'haeb:	data_out=16'h4;
17'haec:	data_out=16'h4;
17'haed:	data_out=16'h5;
17'haee:	data_out=16'h8003;
17'haef:	data_out=16'h8004;
17'haf0:	data_out=16'h1;
17'haf1:	data_out=16'h5;
17'haf2:	data_out=16'h6;
17'haf3:	data_out=16'h8002;
17'haf4:	data_out=16'h8004;
17'haf5:	data_out=16'h8;
17'haf6:	data_out=16'h6;
17'haf7:	data_out=16'h8005;
17'haf8:	data_out=16'h8001;
17'haf9:	data_out=16'h3;
17'hafa:	data_out=16'h8005;
17'hafb:	data_out=16'h8003;
17'hafc:	data_out=16'h8009;
17'hafd:	data_out=16'h5;
17'hafe:	data_out=16'h8004;
17'haff:	data_out=16'h8000;
17'hb00:	data_out=16'h8001;
17'hb01:	data_out=16'h5;
17'hb02:	data_out=16'h4;
17'hb03:	data_out=16'h6;
17'hb04:	data_out=16'h8007;
17'hb05:	data_out=16'h1;
17'hb06:	data_out=16'h4;
17'hb07:	data_out=16'h8002;
17'hb08:	data_out=16'h8000;
17'hb09:	data_out=16'h7;
17'hb0a:	data_out=16'h8007;
17'hb0b:	data_out=16'h8005;
17'hb0c:	data_out=16'h3;
17'hb0d:	data_out=16'h8000;
17'hb0e:	data_out=16'h0;
17'hb0f:	data_out=16'h8005;
17'hb10:	data_out=16'h8004;
17'hb11:	data_out=16'h8003;
17'hb12:	data_out=16'h1;
17'hb13:	data_out=16'h2;
17'hb14:	data_out=16'h8004;
17'hb15:	data_out=16'h8002;
17'hb16:	data_out=16'h6;
17'hb17:	data_out=16'h4;
17'hb18:	data_out=16'h8008;
17'hb19:	data_out=16'h8008;
17'hb1a:	data_out=16'h8008;
17'hb1b:	data_out=16'h8008;
17'hb1c:	data_out=16'h6;
17'hb1d:	data_out=16'h8004;
17'hb1e:	data_out=16'h1;
17'hb1f:	data_out=16'h8004;
17'hb20:	data_out=16'h8007;
17'hb21:	data_out=16'h8005;
17'hb22:	data_out=16'h8006;
17'hb23:	data_out=16'h8005;
17'hb24:	data_out=16'h6;
17'hb25:	data_out=16'h7;
17'hb26:	data_out=16'h2;
17'hb27:	data_out=16'h8004;
17'hb28:	data_out=16'h5;
17'hb29:	data_out=16'h5;
17'hb2a:	data_out=16'h0;
17'hb2b:	data_out=16'h8002;
17'hb2c:	data_out=16'h8005;
17'hb2d:	data_out=16'h8008;
17'hb2e:	data_out=16'h2;
17'hb2f:	data_out=16'h1;
17'hb30:	data_out=16'h8002;
17'hb31:	data_out=16'h8006;
17'hb32:	data_out=16'h8007;
17'hb33:	data_out=16'h3;
17'hb34:	data_out=16'h1;
17'hb35:	data_out=16'h8;
17'hb36:	data_out=16'h8002;
17'hb37:	data_out=16'h2;
17'hb38:	data_out=16'h9;
17'hb39:	data_out=16'h8001;
17'hb3a:	data_out=16'h3;
17'hb3b:	data_out=16'h6;
17'hb3c:	data_out=16'h4;
17'hb3d:	data_out=16'h8006;
17'hb3e:	data_out=16'h8007;
17'hb3f:	data_out=16'h6;
17'hb40:	data_out=16'h8001;
17'hb41:	data_out=16'h8004;
17'hb42:	data_out=16'h8008;
17'hb43:	data_out=16'h8005;
17'hb44:	data_out=16'h8006;
17'hb45:	data_out=16'h3;
17'hb46:	data_out=16'h1;
17'hb47:	data_out=16'h8;
17'hb48:	data_out=16'h8001;
17'hb49:	data_out=16'h8008;
17'hb4a:	data_out=16'h8003;
17'hb4b:	data_out=16'h4;
17'hb4c:	data_out=16'h8007;
17'hb4d:	data_out=16'h8;
17'hb4e:	data_out=16'h8005;
17'hb4f:	data_out=16'h0;
17'hb50:	data_out=16'h8006;
17'hb51:	data_out=16'h8003;
17'hb52:	data_out=16'h8006;
17'hb53:	data_out=16'h4;
17'hb54:	data_out=16'h8004;
17'hb55:	data_out=16'h1;
17'hb56:	data_out=16'h8003;
17'hb57:	data_out=16'h8004;
17'hb58:	data_out=16'h8009;
17'hb59:	data_out=16'h9;
17'hb5a:	data_out=16'h8007;
17'hb5b:	data_out=16'h5;
17'hb5c:	data_out=16'h8006;
17'hb5d:	data_out=16'h8005;
17'hb5e:	data_out=16'h2;
17'hb5f:	data_out=16'h2;
17'hb60:	data_out=16'h1;
17'hb61:	data_out=16'h3;
17'hb62:	data_out=16'h6;
17'hb63:	data_out=16'h4;
17'hb64:	data_out=16'h8003;
17'hb65:	data_out=16'h8002;
17'hb66:	data_out=16'h3;
17'hb67:	data_out=16'h5;
17'hb68:	data_out=16'h8001;
17'hb69:	data_out=16'h8008;
17'hb6a:	data_out=16'h0;
17'hb6b:	data_out=16'h2;
17'hb6c:	data_out=16'h9;
17'hb6d:	data_out=16'h4;
17'hb6e:	data_out=16'h8007;
17'hb6f:	data_out=16'h8007;
17'hb70:	data_out=16'h8007;
17'hb71:	data_out=16'h8004;
17'hb72:	data_out=16'h6;
17'hb73:	data_out=16'h8002;
17'hb74:	data_out=16'h7;
17'hb75:	data_out=16'h8006;
17'hb76:	data_out=16'h3;
17'hb77:	data_out=16'h7;
17'hb78:	data_out=16'h8007;
17'hb79:	data_out=16'h5;
17'hb7a:	data_out=16'h2;
17'hb7b:	data_out=16'h8004;
17'hb7c:	data_out=16'h8009;
17'hb7d:	data_out=16'h8005;
17'hb7e:	data_out=16'h7;
17'hb7f:	data_out=16'h1;
17'hb80:	data_out=16'h6;
17'hb81:	data_out=16'h4;
17'hb82:	data_out=16'h8004;
17'hb83:	data_out=16'h8006;
17'hb84:	data_out=16'h8007;
17'hb85:	data_out=16'h8;
17'hb86:	data_out=16'h9;
17'hb87:	data_out=16'h2;
17'hb88:	data_out=16'h9;
17'hb89:	data_out=16'h8000;
17'hb8a:	data_out=16'h8006;
17'hb8b:	data_out=16'h9;
17'hb8c:	data_out=16'h8005;
17'hb8d:	data_out=16'h8004;
17'hb8e:	data_out=16'h8007;
17'hb8f:	data_out=16'h8003;
17'hb90:	data_out=16'h1;
17'hb91:	data_out=16'h9;
17'hb92:	data_out=16'h4;
17'hb93:	data_out=16'h8001;
17'hb94:	data_out=16'h8006;
17'hb95:	data_out=16'h8002;
17'hb96:	data_out=16'h8004;
17'hb97:	data_out=16'h8004;
17'hb98:	data_out=16'h8006;
17'hb99:	data_out=16'h7;
17'hb9a:	data_out=16'h2;
17'hb9b:	data_out=16'h8006;
17'hb9c:	data_out=16'h8007;
17'hb9d:	data_out=16'h8000;
17'hb9e:	data_out=16'h4;
17'hb9f:	data_out=16'h8;
17'hba0:	data_out=16'h8005;
17'hba1:	data_out=16'h8009;
17'hba2:	data_out=16'h8007;
17'hba3:	data_out=16'h8002;
17'hba4:	data_out=16'h8;
17'hba5:	data_out=16'h8007;
17'hba6:	data_out=16'h9;
17'hba7:	data_out=16'h8;
17'hba8:	data_out=16'h1;
17'hba9:	data_out=16'h8006;
17'hbaa:	data_out=16'h8;
17'hbab:	data_out=16'h5;
17'hbac:	data_out=16'h8001;
17'hbad:	data_out=16'h8008;
17'hbae:	data_out=16'h8007;
17'hbaf:	data_out=16'h8009;
17'hbb0:	data_out=16'h8008;
17'hbb1:	data_out=16'h6;
17'hbb2:	data_out=16'h8001;
17'hbb3:	data_out=16'h8005;
17'hbb4:	data_out=16'h8006;
17'hbb5:	data_out=16'h4;
17'hbb6:	data_out=16'h1;
17'hbb7:	data_out=16'h8003;
17'hbb8:	data_out=16'h2;
17'hbb9:	data_out=16'h8007;
17'hbba:	data_out=16'h0;
17'hbbb:	data_out=16'h4;
17'hbbc:	data_out=16'h2;
17'hbbd:	data_out=16'h8005;
17'hbbe:	data_out=16'h3;
17'hbbf:	data_out=16'h7;
17'hbc0:	data_out=16'h8004;
17'hbc1:	data_out=16'h5;
17'hbc2:	data_out=16'h8004;
17'hbc3:	data_out=16'h8005;
17'hbc4:	data_out=16'h7;
17'hbc5:	data_out=16'h8005;
17'hbc6:	data_out=16'h8006;
17'hbc7:	data_out=16'h8001;
17'hbc8:	data_out=16'h8002;
17'hbc9:	data_out=16'h8007;
17'hbca:	data_out=16'h8005;
17'hbcb:	data_out=16'h6;
17'hbcc:	data_out=16'h8005;
17'hbcd:	data_out=16'h8003;
17'hbce:	data_out=16'h7;
17'hbcf:	data_out=16'h8004;
17'hbd0:	data_out=16'h8006;
17'hbd1:	data_out=16'h8004;
17'hbd2:	data_out=16'h0;
17'hbd3:	data_out=16'h8002;
17'hbd4:	data_out=16'h8009;
17'hbd5:	data_out=16'h8008;
17'hbd6:	data_out=16'h4;
17'hbd7:	data_out=16'h2;
17'hbd8:	data_out=16'h8006;
17'hbd9:	data_out=16'h8005;
17'hbda:	data_out=16'h8003;
17'hbdb:	data_out=16'h6;
17'hbdc:	data_out=16'h8000;
17'hbdd:	data_out=16'h9;
17'hbde:	data_out=16'h4;
17'hbdf:	data_out=16'h5;
17'hbe0:	data_out=16'h5;
17'hbe1:	data_out=16'h8;
17'hbe2:	data_out=16'h9;
17'hbe3:	data_out=16'h2;
17'hbe4:	data_out=16'h8006;
17'hbe5:	data_out=16'h8006;
17'hbe6:	data_out=16'h8008;
17'hbe7:	data_out=16'h2;
17'hbe8:	data_out=16'h8004;
17'hbe9:	data_out=16'h8003;
17'hbea:	data_out=16'h8001;
17'hbeb:	data_out=16'h8000;
17'hbec:	data_out=16'h3;
17'hbed:	data_out=16'h8004;
17'hbee:	data_out=16'h5;
17'hbef:	data_out=16'h6;
17'hbf0:	data_out=16'h2;
17'hbf1:	data_out=16'h8004;
17'hbf2:	data_out=16'h8005;
17'hbf3:	data_out=16'h2;
17'hbf4:	data_out=16'h8003;
17'hbf5:	data_out=16'h8;
17'hbf6:	data_out=16'h8005;
17'hbf7:	data_out=16'h0;
17'hbf8:	data_out=16'h8006;
17'hbf9:	data_out=16'h1;
17'hbfa:	data_out=16'h8003;
17'hbfb:	data_out=16'h3;
17'hbfc:	data_out=16'h0;
17'hbfd:	data_out=16'h8009;
17'hbfe:	data_out=16'h8001;
17'hbff:	data_out=16'h8004;
17'hc00:	data_out=16'h9;
17'hc01:	data_out=16'h8002;
17'hc02:	data_out=16'h7;
17'hc03:	data_out=16'h8006;
17'hc04:	data_out=16'h1;
17'hc05:	data_out=16'h8;
17'hc06:	data_out=16'h5;
17'hc07:	data_out=16'h6;
17'hc08:	data_out=16'h8004;
17'hc09:	data_out=16'h8006;
17'hc0a:	data_out=16'h8004;
17'hc0b:	data_out=16'h8;
17'hc0c:	data_out=16'h8000;
17'hc0d:	data_out=16'h8008;
17'hc0e:	data_out=16'h5;
17'hc0f:	data_out=16'h8008;
17'hc10:	data_out=16'h8003;
17'hc11:	data_out=16'h8009;
17'hc12:	data_out=16'h3;
17'hc13:	data_out=16'h3;
17'hc14:	data_out=16'h8;
17'hc15:	data_out=16'h7;
17'hc16:	data_out=16'h8006;
17'hc17:	data_out=16'h8007;
17'hc18:	data_out=16'h8001;
17'hc19:	data_out=16'h0;
17'hc1a:	data_out=16'h6;
17'hc1b:	data_out=16'h8;
17'hc1c:	data_out=16'h1;
17'hc1d:	data_out=16'h8004;
17'hc1e:	data_out=16'h8006;
17'hc1f:	data_out=16'h0;
17'hc20:	data_out=16'h3;
17'hc21:	data_out=16'h8008;
17'hc22:	data_out=16'h3;
17'hc23:	data_out=16'h8005;
17'hc24:	data_out=16'h8008;
17'hc25:	data_out=16'h8001;
17'hc26:	data_out=16'h8008;
17'hc27:	data_out=16'h8003;
17'hc28:	data_out=16'h3;
17'hc29:	data_out=16'h8003;
17'hc2a:	data_out=16'h8004;
17'hc2b:	data_out=16'h8007;
17'hc2c:	data_out=16'h8002;
17'hc2d:	data_out=16'h8008;
17'hc2e:	data_out=16'h8005;
17'hc2f:	data_out=16'h4;
17'hc30:	data_out=16'h8008;
17'hc31:	data_out=16'h7;
17'hc32:	data_out=16'h8002;
17'hc33:	data_out=16'h8009;
17'hc34:	data_out=16'h5;
17'hc35:	data_out=16'h2;
17'hc36:	data_out=16'h8006;
17'hc37:	data_out=16'h8006;
17'hc38:	data_out=16'h8007;
17'hc39:	data_out=16'h8009;
17'hc3a:	data_out=16'h8007;
17'hc3b:	data_out=16'h3;
17'hc3c:	data_out=16'h8004;
17'hc3d:	data_out=16'h8003;
17'hc3e:	data_out=16'h8006;
17'hc3f:	data_out=16'h8;
17'hc40:	data_out=16'h8002;
17'hc41:	data_out=16'h7;
17'hc42:	data_out=16'h8006;
17'hc43:	data_out=16'h8001;
17'hc44:	data_out=16'h8003;
17'hc45:	data_out=16'h8005;
17'hc46:	data_out=16'h5;
17'hc47:	data_out=16'h8;
17'hc48:	data_out=16'h1;
17'hc49:	data_out=16'h8008;
17'hc4a:	data_out=16'h8007;
17'hc4b:	data_out=16'h9;
17'hc4c:	data_out=16'h8007;
17'hc4d:	data_out=16'h8004;
17'hc4e:	data_out=16'h4;
17'hc4f:	data_out=16'h8005;
17'hc50:	data_out=16'h8006;
17'hc51:	data_out=16'h8007;
17'hc52:	data_out=16'h8005;
17'hc53:	data_out=16'h9;
17'hc54:	data_out=16'h4;
17'hc55:	data_out=16'h8002;
17'hc56:	data_out=16'h8006;
17'hc57:	data_out=16'h6;
17'hc58:	data_out=16'h8002;
17'hc59:	data_out=16'h8004;
17'hc5a:	data_out=16'h8001;
17'hc5b:	data_out=16'h3;
17'hc5c:	data_out=16'h2;
17'hc5d:	data_out=16'h3;
17'hc5e:	data_out=16'h2;
17'hc5f:	data_out=16'h8008;
17'hc60:	data_out=16'h0;
17'hc61:	data_out=16'h6;
17'hc62:	data_out=16'h0;
17'hc63:	data_out=16'h6;
17'hc64:	data_out=16'h8009;
17'hc65:	data_out=16'h8004;
17'hc66:	data_out=16'h5;
17'hc67:	data_out=16'h2;
17'hc68:	data_out=16'h8003;
17'hc69:	data_out=16'h7;
17'hc6a:	data_out=16'h1;
17'hc6b:	data_out=16'h8000;
17'hc6c:	data_out=16'h8006;
17'hc6d:	data_out=16'h8004;
17'hc6e:	data_out=16'h4;
17'hc6f:	data_out=16'h8002;
17'hc70:	data_out=16'h8002;
17'hc71:	data_out=16'h8;
17'hc72:	data_out=16'h8003;
17'hc73:	data_out=16'h8008;
17'hc74:	data_out=16'h8003;
17'hc75:	data_out=16'h0;
17'hc76:	data_out=16'h7;
17'hc77:	data_out=16'h5;
17'hc78:	data_out=16'h6;
17'hc79:	data_out=16'h8003;
17'hc7a:	data_out=16'h8001;
17'hc7b:	data_out=16'h8001;
17'hc7c:	data_out=16'h9;
17'hc7d:	data_out=16'h8008;
17'hc7e:	data_out=16'h0;
17'hc7f:	data_out=16'h0;
17'hc80:	data_out=16'h7;
17'hc81:	data_out=16'h8009;
17'hc82:	data_out=16'h8003;
17'hc83:	data_out=16'h7;
17'hc84:	data_out=16'h8003;
17'hc85:	data_out=16'h8006;
17'hc86:	data_out=16'h8000;
17'hc87:	data_out=16'h3;
17'hc88:	data_out=16'h8008;
17'hc89:	data_out=16'h8008;
17'hc8a:	data_out=16'h8006;
17'hc8b:	data_out=16'h8005;
17'hc8c:	data_out=16'h8004;
17'hc8d:	data_out=16'h7;
17'hc8e:	data_out=16'h2;
17'hc8f:	data_out=16'h3;
17'hc90:	data_out=16'h5;
17'hc91:	data_out=16'h9;
17'hc92:	data_out=16'h4;
17'hc93:	data_out=16'h8007;
17'hc94:	data_out=16'h0;
17'hc95:	data_out=16'h2;
17'hc96:	data_out=16'h7;
17'hc97:	data_out=16'h8003;
17'hc98:	data_out=16'h8;
17'hc99:	data_out=16'h8003;
17'hc9a:	data_out=16'h5;
17'hc9b:	data_out=16'h8;
17'hc9c:	data_out=16'h8002;
17'hc9d:	data_out=16'h8004;
17'hc9e:	data_out=16'h8001;
17'hc9f:	data_out=16'h8004;
17'hca0:	data_out=16'h8003;
17'hca1:	data_out=16'h5;
17'hca2:	data_out=16'h8006;
17'hca3:	data_out=16'h3;
17'hca4:	data_out=16'h8;
17'hca5:	data_out=16'h3;
17'hca6:	data_out=16'h8003;
17'hca7:	data_out=16'h9;
17'hca8:	data_out=16'h4;
17'hca9:	data_out=16'h0;
17'hcaa:	data_out=16'h8005;
17'hcab:	data_out=16'h9;
17'hcac:	data_out=16'h8002;
17'hcad:	data_out=16'h6;
17'hcae:	data_out=16'h3;
17'hcaf:	data_out=16'h8006;
17'hcb0:	data_out=16'h6;
17'hcb1:	data_out=16'h8002;
17'hcb2:	data_out=16'h8003;
17'hcb3:	data_out=16'h8003;
17'hcb4:	data_out=16'h9;
17'hcb5:	data_out=16'h8005;
17'hcb6:	data_out=16'h3;
17'hcb7:	data_out=16'h8;
17'hcb8:	data_out=16'h1;
17'hcb9:	data_out=16'h8000;
17'hcba:	data_out=16'h7;
17'hcbb:	data_out=16'h9;
17'hcbc:	data_out=16'h5;
17'hcbd:	data_out=16'h8003;
17'hcbe:	data_out=16'h8004;
17'hcbf:	data_out=16'h8007;
17'hcc0:	data_out=16'h8007;
17'hcc1:	data_out=16'h8001;
17'hcc2:	data_out=16'h5;
17'hcc3:	data_out=16'h8008;
17'hcc4:	data_out=16'h8007;
17'hcc5:	data_out=16'h8007;
17'hcc6:	data_out=16'h8008;
17'hcc7:	data_out=16'h6;
17'hcc8:	data_out=16'h2;
17'hcc9:	data_out=16'h8004;
17'hcca:	data_out=16'h6;
17'hccb:	data_out=16'h8009;
17'hccc:	data_out=16'h8007;
17'hccd:	data_out=16'h8001;
17'hcce:	data_out=16'h8005;
17'hccf:	data_out=16'h8;
17'hcd0:	data_out=16'h6;
17'hcd1:	data_out=16'h1;
17'hcd2:	data_out=16'h8004;
17'hcd3:	data_out=16'h6;
17'hcd4:	data_out=16'h5;
17'hcd5:	data_out=16'h8;
17'hcd6:	data_out=16'h5;
17'hcd7:	data_out=16'h8003;
17'hcd8:	data_out=16'h8001;
17'hcd9:	data_out=16'h3;
17'hcda:	data_out=16'h8003;
17'hcdb:	data_out=16'h8005;
17'hcdc:	data_out=16'h8009;
17'hcdd:	data_out=16'h1;
17'hcde:	data_out=16'h8003;
17'hcdf:	data_out=16'h8006;
17'hce0:	data_out=16'h8009;
17'hce1:	data_out=16'h8007;
17'hce2:	data_out=16'h8005;
17'hce3:	data_out=16'h8007;
17'hce4:	data_out=16'h8005;
17'hce5:	data_out=16'h8003;
17'hce6:	data_out=16'h8;
17'hce7:	data_out=16'h6;
17'hce8:	data_out=16'h2;
17'hce9:	data_out=16'h4;
17'hcea:	data_out=16'h7;
17'hceb:	data_out=16'h4;
17'hcec:	data_out=16'h8006;
17'hced:	data_out=16'h8008;
17'hcee:	data_out=16'h3;
17'hcef:	data_out=16'h8008;
17'hcf0:	data_out=16'h2;
17'hcf1:	data_out=16'h8;
17'hcf2:	data_out=16'h7;
17'hcf3:	data_out=16'h8002;
17'hcf4:	data_out=16'h7;
17'hcf5:	data_out=16'h3;
17'hcf6:	data_out=16'h4;
17'hcf7:	data_out=16'h8003;
17'hcf8:	data_out=16'h8002;
17'hcf9:	data_out=16'h8008;
17'hcfa:	data_out=16'h1;
17'hcfb:	data_out=16'h8002;
17'hcfc:	data_out=16'h2;
17'hcfd:	data_out=16'h7;
17'hcfe:	data_out=16'h1;
17'hcff:	data_out=16'h2;
17'hd00:	data_out=16'h9;
17'hd01:	data_out=16'h6;
17'hd02:	data_out=16'h4;
17'hd03:	data_out=16'h8006;
17'hd04:	data_out=16'h8007;
17'hd05:	data_out=16'h3;
17'hd06:	data_out=16'h8009;
17'hd07:	data_out=16'h4;
17'hd08:	data_out=16'h8002;
17'hd09:	data_out=16'h7;
17'hd0a:	data_out=16'h8001;
17'hd0b:	data_out=16'h2;
17'hd0c:	data_out=16'h8;
17'hd0d:	data_out=16'h8007;
17'hd0e:	data_out=16'h2;
17'hd0f:	data_out=16'h1;
17'hd10:	data_out=16'h8008;
17'hd11:	data_out=16'h0;
17'hd12:	data_out=16'h9;
17'hd13:	data_out=16'h8;
17'hd14:	data_out=16'h8005;
17'hd15:	data_out=16'h4;
17'hd16:	data_out=16'h8004;
17'hd17:	data_out=16'h2;
17'hd18:	data_out=16'h4;
17'hd19:	data_out=16'h6;
17'hd1a:	data_out=16'h9;
17'hd1b:	data_out=16'h8003;
17'hd1c:	data_out=16'h4;
17'hd1d:	data_out=16'h1;
17'hd1e:	data_out=16'h8;
17'hd1f:	data_out=16'h4;
17'hd20:	data_out=16'h8003;
17'hd21:	data_out=16'h3;
17'hd22:	data_out=16'h7;
17'hd23:	data_out=16'h8000;
17'hd24:	data_out=16'h8003;
17'hd25:	data_out=16'h7;
17'hd26:	data_out=16'h8006;
17'hd27:	data_out=16'h4;
17'hd28:	data_out=16'h5;
17'hd29:	data_out=16'h2;
17'hd2a:	data_out=16'h8003;
17'hd2b:	data_out=16'h4;
17'hd2c:	data_out=16'h4;
17'hd2d:	data_out=16'h8;
17'hd2e:	data_out=16'h8003;
17'hd2f:	data_out=16'h5;
17'hd30:	data_out=16'h8000;
17'hd31:	data_out=16'h8004;
17'hd32:	data_out=16'h4;
17'hd33:	data_out=16'h4;
17'hd34:	data_out=16'h9;
17'hd35:	data_out=16'h8009;
17'hd36:	data_out=16'h8004;
17'hd37:	data_out=16'h4;
17'hd38:	data_out=16'h6;
17'hd39:	data_out=16'h8004;
17'hd3a:	data_out=16'h8008;
17'hd3b:	data_out=16'h1;
17'hd3c:	data_out=16'h6;
17'hd3d:	data_out=16'h8009;
17'hd3e:	data_out=16'h8004;
17'hd3f:	data_out=16'h8006;
17'hd40:	data_out=16'h4;
17'hd41:	data_out=16'h8006;
17'hd42:	data_out=16'h2;
17'hd43:	data_out=16'h8008;
17'hd44:	data_out=16'h8008;
17'hd45:	data_out=16'h6;
17'hd46:	data_out=16'h5;
17'hd47:	data_out=16'h6;
17'hd48:	data_out=16'h8001;
17'hd49:	data_out=16'h8007;
17'hd4a:	data_out=16'h2;
17'hd4b:	data_out=16'h8006;
17'hd4c:	data_out=16'h8008;
17'hd4d:	data_out=16'h7;
17'hd4e:	data_out=16'h8;
17'hd4f:	data_out=16'h1;
17'hd50:	data_out=16'h8006;
17'hd51:	data_out=16'h3;
17'hd52:	data_out=16'h8004;
17'hd53:	data_out=16'h8006;
17'hd54:	data_out=16'h3;
17'hd55:	data_out=16'h1;
17'hd56:	data_out=16'h7;
17'hd57:	data_out=16'h1;
17'hd58:	data_out=16'h6;
17'hd59:	data_out=16'h8;
17'hd5a:	data_out=16'h8007;
17'hd5b:	data_out=16'h2;
17'hd5c:	data_out=16'h8;
17'hd5d:	data_out=16'h8002;
17'hd5e:	data_out=16'h5;
17'hd5f:	data_out=16'h2;
17'hd60:	data_out=16'h1;
17'hd61:	data_out=16'h8002;
17'hd62:	data_out=16'h3;
17'hd63:	data_out=16'h2;
17'hd64:	data_out=16'h8005;
17'hd65:	data_out=16'h8001;
17'hd66:	data_out=16'h8000;
17'hd67:	data_out=16'h4;
17'hd68:	data_out=16'h1;
17'hd69:	data_out=16'h8008;
17'hd6a:	data_out=16'h7;
17'hd6b:	data_out=16'h2;
17'hd6c:	data_out=16'h8;
17'hd6d:	data_out=16'h6;
17'hd6e:	data_out=16'h8006;
17'hd6f:	data_out=16'h8007;
17'hd70:	data_out=16'h0;
17'hd71:	data_out=16'h8001;
17'hd72:	data_out=16'h8004;
17'hd73:	data_out=16'h8005;
17'hd74:	data_out=16'h9;
17'hd75:	data_out=16'h8006;
17'hd76:	data_out=16'h4;
17'hd77:	data_out=16'h5;
17'hd78:	data_out=16'h8008;
17'hd79:	data_out=16'h7;
17'hd7a:	data_out=16'h8002;
17'hd7b:	data_out=16'h9;
17'hd7c:	data_out=16'h8004;
17'hd7d:	data_out=16'h8006;
17'hd7e:	data_out=16'h2;
17'hd7f:	data_out=16'h6;
17'hd80:	data_out=16'h2;
17'hd81:	data_out=16'h8004;
17'hd82:	data_out=16'h8001;
17'hd83:	data_out=16'h6;
17'hd84:	data_out=16'h4;
17'hd85:	data_out=16'h8;
17'hd86:	data_out=16'h0;
17'hd87:	data_out=16'h8005;
17'hd88:	data_out=16'h9;
17'hd89:	data_out=16'h8002;
17'hd8a:	data_out=16'h7;
17'hd8b:	data_out=16'h8;
17'hd8c:	data_out=16'h8005;
17'hd8d:	data_out=16'h8008;
17'hd8e:	data_out=16'h8008;
17'hd8f:	data_out=16'h5;
17'hd90:	data_out=16'h8000;
17'hd91:	data_out=16'h8002;
17'hd92:	data_out=16'h8;
17'hd93:	data_out=16'h8001;
17'hd94:	data_out=16'h0;
17'hd95:	data_out=16'h4;
17'hd96:	data_out=16'h8005;
17'hd97:	data_out=16'h2;
17'hd98:	data_out=16'h1;
17'hd99:	data_out=16'h3;
17'hd9a:	data_out=16'h1;
17'hd9b:	data_out=16'h6;
17'hd9c:	data_out=16'h6;
17'hd9d:	data_out=16'h8006;
17'hd9e:	data_out=16'h3;
17'hd9f:	data_out=16'h8001;
17'hda0:	data_out=16'h8001;
17'hda1:	data_out=16'h8007;
17'hda2:	data_out=16'h8004;
17'hda3:	data_out=16'h8007;
17'hda4:	data_out=16'h8009;
17'hda5:	data_out=16'h5;
17'hda6:	data_out=16'h8003;
17'hda7:	data_out=16'h8009;
17'hda8:	data_out=16'h8006;
17'hda9:	data_out=16'h8005;
17'hdaa:	data_out=16'h8;
17'hdab:	data_out=16'h8001;
17'hdac:	data_out=16'h8004;
17'hdad:	data_out=16'h8008;
17'hdae:	data_out=16'h8006;
17'hdaf:	data_out=16'h4;
17'hdb0:	data_out=16'h8002;
17'hdb1:	data_out=16'h8007;
17'hdb2:	data_out=16'h8006;
17'hdb3:	data_out=16'h8;
17'hdb4:	data_out=16'h6;
17'hdb5:	data_out=16'h8001;
17'hdb6:	data_out=16'h0;
17'hdb7:	data_out=16'h8002;
17'hdb8:	data_out=16'h8007;
17'hdb9:	data_out=16'h8008;
17'hdba:	data_out=16'h8005;
17'hdbb:	data_out=16'h8;
17'hdbc:	data_out=16'h8005;
17'hdbd:	data_out=16'h7;
17'hdbe:	data_out=16'h8002;
17'hdbf:	data_out=16'h3;
17'hdc0:	data_out=16'h8;
17'hdc1:	data_out=16'h2;
17'hdc2:	data_out=16'h5;
17'hdc3:	data_out=16'h9;
17'hdc4:	data_out=16'h8002;
17'hdc5:	data_out=16'h8007;
17'hdc6:	data_out=16'h9;
17'hdc7:	data_out=16'h2;
17'hdc8:	data_out=16'h8003;
17'hdc9:	data_out=16'h8;
17'hdca:	data_out=16'h8009;
17'hdcb:	data_out=16'h2;
17'hdcc:	data_out=16'h9;
17'hdcd:	data_out=16'h8006;
17'hdce:	data_out=16'h8003;
17'hdcf:	data_out=16'h8002;
17'hdd0:	data_out=16'h8003;
17'hdd1:	data_out=16'h1;
17'hdd2:	data_out=16'h8003;
17'hdd3:	data_out=16'h8007;
17'hdd4:	data_out=16'h9;
17'hdd5:	data_out=16'h7;
17'hdd6:	data_out=16'h1;
17'hdd7:	data_out=16'h8008;
17'hdd8:	data_out=16'h8;
17'hdd9:	data_out=16'h5;
17'hdda:	data_out=16'h8009;
17'hddb:	data_out=16'h8006;
17'hddc:	data_out=16'h2;
17'hddd:	data_out=16'h8002;
17'hdde:	data_out=16'h7;
17'hddf:	data_out=16'h1;
17'hde0:	data_out=16'h8009;
17'hde1:	data_out=16'h3;
17'hde2:	data_out=16'h1;
17'hde3:	data_out=16'h8001;
17'hde4:	data_out=16'h5;
17'hde5:	data_out=16'h1;
17'hde6:	data_out=16'h8009;
17'hde7:	data_out=16'h8007;
17'hde8:	data_out=16'h8000;
17'hde9:	data_out=16'h8009;
17'hdea:	data_out=16'h5;
17'hdeb:	data_out=16'h8000;
17'hdec:	data_out=16'h8005;
17'hded:	data_out=16'h8007;
17'hdee:	data_out=16'h7;
17'hdef:	data_out=16'h0;
17'hdf0:	data_out=16'h3;
17'hdf1:	data_out=16'h8005;
17'hdf2:	data_out=16'h3;
17'hdf3:	data_out=16'h2;
17'hdf4:	data_out=16'h8008;
17'hdf5:	data_out=16'h8006;
17'hdf6:	data_out=16'h4;
17'hdf7:	data_out=16'h8009;
17'hdf8:	data_out=16'h8;
17'hdf9:	data_out=16'h4;
17'hdfa:	data_out=16'h8005;
17'hdfb:	data_out=16'h1;
17'hdfc:	data_out=16'h8007;
17'hdfd:	data_out=16'h8007;
17'hdfe:	data_out=16'h8007;
17'hdff:	data_out=16'h8007;
17'he00:	data_out=16'h4;
17'he01:	data_out=16'h4;
17'he02:	data_out=16'h1;
17'he03:	data_out=16'h0;
17'he04:	data_out=16'h8005;
17'he05:	data_out=16'h1;
17'he06:	data_out=16'h3;
17'he07:	data_out=16'h4;
17'he08:	data_out=16'h2;
17'he09:	data_out=16'h8001;
17'he0a:	data_out=16'h8005;
17'he0b:	data_out=16'h5;
17'he0c:	data_out=16'h0;
17'he0d:	data_out=16'h8007;
17'he0e:	data_out=16'h8003;
17'he0f:	data_out=16'h8006;
17'he10:	data_out=16'h8003;
17'he11:	data_out=16'h9;
17'he12:	data_out=16'h5;
17'he13:	data_out=16'h8002;
17'he14:	data_out=16'h8006;
17'he15:	data_out=16'h8000;
17'he16:	data_out=16'h8001;
17'he17:	data_out=16'h8007;
17'he18:	data_out=16'h8005;
17'he19:	data_out=16'h3;
17'he1a:	data_out=16'h3;
17'he1b:	data_out=16'h8004;
17'he1c:	data_out=16'h4;
17'he1d:	data_out=16'h6;
17'he1e:	data_out=16'h8001;
17'he1f:	data_out=16'h8000;
17'he20:	data_out=16'h0;
17'he21:	data_out=16'h9;
17'he22:	data_out=16'h8009;
17'he23:	data_out=16'h5;
17'he24:	data_out=16'h1;
17'he25:	data_out=16'h3;
17'he26:	data_out=16'h8000;
17'he27:	data_out=16'h8007;
17'he28:	data_out=16'h8007;
17'he29:	data_out=16'h4;
17'he2a:	data_out=16'h8;
17'he2b:	data_out=16'h2;
17'he2c:	data_out=16'h5;
17'he2d:	data_out=16'h8005;
17'he2e:	data_out=16'h5;
17'he2f:	data_out=16'h8007;
17'he30:	data_out=16'h8005;
17'he31:	data_out=16'h1;
17'he32:	data_out=16'h0;
17'he33:	data_out=16'h8002;
17'he34:	data_out=16'h8008;
17'he35:	data_out=16'h8;
17'he36:	data_out=16'h0;
17'he37:	data_out=16'h8004;
17'he38:	data_out=16'h2;
17'he39:	data_out=16'h8006;
17'he3a:	data_out=16'h1;
17'he3b:	data_out=16'h8003;
17'he3c:	data_out=16'h8009;
17'he3d:	data_out=16'h9;
17'he3e:	data_out=16'h6;
17'he3f:	data_out=16'h1;
17'he40:	data_out=16'h8;
17'he41:	data_out=16'h6;
17'he42:	data_out=16'h8004;
17'he43:	data_out=16'h0;
17'he44:	data_out=16'h0;
17'he45:	data_out=16'h5;
17'he46:	data_out=16'h3;
17'he47:	data_out=16'h2;
17'he48:	data_out=16'h8000;
17'he49:	data_out=16'h1;
17'he4a:	data_out=16'h8005;
17'he4b:	data_out=16'h8004;
17'he4c:	data_out=16'h6;
17'he4d:	data_out=16'h8009;
17'he4e:	data_out=16'h8002;
17'he4f:	data_out=16'h8008;
17'he50:	data_out=16'h2;
17'he51:	data_out=16'h8;
17'he52:	data_out=16'h8001;
17'he53:	data_out=16'h3;
17'he54:	data_out=16'h7;
17'he55:	data_out=16'h8;
17'he56:	data_out=16'h7;
17'he57:	data_out=16'h8000;
17'he58:	data_out=16'h8007;
17'he59:	data_out=16'h8001;
17'he5a:	data_out=16'h6;
17'he5b:	data_out=16'h8006;
17'he5c:	data_out=16'h8001;
17'he5d:	data_out=16'h3;
17'he5e:	data_out=16'h3;
17'he5f:	data_out=16'h8002;
17'he60:	data_out=16'h0;
17'he61:	data_out=16'h9;
17'he62:	data_out=16'h8;
17'he63:	data_out=16'h8008;
17'he64:	data_out=16'h5;
17'he65:	data_out=16'h1;
17'he66:	data_out=16'h3;
17'he67:	data_out=16'h8004;
17'he68:	data_out=16'h8007;
17'he69:	data_out=16'h7;
17'he6a:	data_out=16'h1;
17'he6b:	data_out=16'h9;
17'he6c:	data_out=16'h8;
17'he6d:	data_out=16'h9;
17'he6e:	data_out=16'h8009;
17'he6f:	data_out=16'h0;
17'he70:	data_out=16'h8;
17'he71:	data_out=16'h8001;
17'he72:	data_out=16'h8006;
17'he73:	data_out=16'h6;
17'he74:	data_out=16'h8002;
17'he75:	data_out=16'h8008;
17'he76:	data_out=16'h8003;
17'he77:	data_out=16'h1;
17'he78:	data_out=16'h0;
17'he79:	data_out=16'h8006;
17'he7a:	data_out=16'h4;
17'he7b:	data_out=16'h8;
17'he7c:	data_out=16'h6;
17'he7d:	data_out=16'h8002;
17'he7e:	data_out=16'h8003;
17'he7f:	data_out=16'h8003;
17'he80:	data_out=16'h8002;
17'he81:	data_out=16'h8004;
17'he82:	data_out=16'h8002;
17'he83:	data_out=16'h8006;
17'he84:	data_out=16'h6;
17'he85:	data_out=16'h8008;
17'he86:	data_out=16'h8001;
17'he87:	data_out=16'h9;
17'he88:	data_out=16'h8;
17'he89:	data_out=16'h9;
17'he8a:	data_out=16'h8;
17'he8b:	data_out=16'h7;
17'he8c:	data_out=16'h9;
17'he8d:	data_out=16'h9;
17'he8e:	data_out=16'h8002;
17'he8f:	data_out=16'h7;
17'he90:	data_out=16'h8001;
17'he91:	data_out=16'h0;
17'he92:	data_out=16'h4;
17'he93:	data_out=16'h6;
17'he94:	data_out=16'h1;
17'he95:	data_out=16'h8009;
17'he96:	data_out=16'h8002;
17'he97:	data_out=16'h8008;
17'he98:	data_out=16'h8006;
17'he99:	data_out=16'h8008;
17'he9a:	data_out=16'h8009;
17'he9b:	data_out=16'h8009;
17'he9c:	data_out=16'h8000;
17'he9d:	data_out=16'h8002;
17'he9e:	data_out=16'h8002;
17'he9f:	data_out=16'h6;
17'hea0:	data_out=16'h3;
17'hea1:	data_out=16'h5;
17'hea2:	data_out=16'h9;
17'hea3:	data_out=16'h0;
17'hea4:	data_out=16'h6;
17'hea5:	data_out=16'h8002;
17'hea6:	data_out=16'h8000;
17'hea7:	data_out=16'h5;
17'hea8:	data_out=16'h8002;
17'hea9:	data_out=16'h8001;
17'heaa:	data_out=16'h2;
17'heab:	data_out=16'h8002;
17'heac:	data_out=16'h8002;
17'head:	data_out=16'h9;
17'heae:	data_out=16'h8004;
17'heaf:	data_out=16'h6;
17'heb0:	data_out=16'h0;
17'heb1:	data_out=16'h8;
17'heb2:	data_out=16'h3;
17'heb3:	data_out=16'h8008;
17'heb4:	data_out=16'h9;
17'heb5:	data_out=16'h8008;
17'heb6:	data_out=16'h8007;
17'heb7:	data_out=16'h8006;
17'heb8:	data_out=16'h8006;
17'heb9:	data_out=16'h8006;
17'heba:	data_out=16'h8006;
17'hebb:	data_out=16'h2;
17'hebc:	data_out=16'h1;
17'hebd:	data_out=16'h0;
17'hebe:	data_out=16'h8001;
17'hebf:	data_out=16'h8005;
17'hec0:	data_out=16'h8004;
17'hec1:	data_out=16'h8001;
17'hec2:	data_out=16'h4;
17'hec3:	data_out=16'h8007;
17'hec4:	data_out=16'h7;
17'hec5:	data_out=16'h8006;
17'hec6:	data_out=16'h7;
17'hec7:	data_out=16'h8004;
17'hec8:	data_out=16'h2;
17'hec9:	data_out=16'h8000;
17'heca:	data_out=16'h2;
17'hecb:	data_out=16'h8009;
17'hecc:	data_out=16'h8001;
17'hecd:	data_out=16'h7;
17'hece:	data_out=16'h6;
17'hecf:	data_out=16'h9;
17'hed0:	data_out=16'h6;
17'hed1:	data_out=16'h0;
17'hed2:	data_out=16'h8008;
17'hed3:	data_out=16'h6;
17'hed4:	data_out=16'h2;
17'hed5:	data_out=16'h8006;
17'hed6:	data_out=16'h9;
17'hed7:	data_out=16'h4;
17'hed8:	data_out=16'h8003;
17'hed9:	data_out=16'h8007;
17'heda:	data_out=16'h8003;
17'hedb:	data_out=16'h7;
17'hedc:	data_out=16'h3;
17'hedd:	data_out=16'h6;
17'hede:	data_out=16'h8008;
17'hedf:	data_out=16'h8;
17'hee0:	data_out=16'h8004;
17'hee1:	data_out=16'h5;
17'hee2:	data_out=16'h8009;
17'hee3:	data_out=16'h8006;
17'hee4:	data_out=16'h9;
17'hee5:	data_out=16'h7;
17'hee6:	data_out=16'h8002;
17'hee7:	data_out=16'h2;
17'hee8:	data_out=16'h8002;
17'hee9:	data_out=16'h8008;
17'heea:	data_out=16'h2;
17'heeb:	data_out=16'h6;
17'heec:	data_out=16'h8;
17'heed:	data_out=16'h8000;
17'heee:	data_out=16'h6;
17'heef:	data_out=16'h5;
17'hef0:	data_out=16'h9;
17'hef1:	data_out=16'h7;
17'hef2:	data_out=16'h2;
17'hef3:	data_out=16'h1;
17'hef4:	data_out=16'h8008;
17'hef5:	data_out=16'h1;
17'hef6:	data_out=16'h8003;
17'hef7:	data_out=16'h8002;
17'hef8:	data_out=16'h3;
17'hef9:	data_out=16'h3;
17'hefa:	data_out=16'h8005;
17'hefb:	data_out=16'h8003;
17'hefc:	data_out=16'h8000;
17'hefd:	data_out=16'h8003;
17'hefe:	data_out=16'h8005;
17'heff:	data_out=16'h5;
17'hf00:	data_out=16'h8007;
17'hf01:	data_out=16'h8004;
17'hf02:	data_out=16'h8;
17'hf03:	data_out=16'h8007;
17'hf04:	data_out=16'h8006;
17'hf05:	data_out=16'h8003;
17'hf06:	data_out=16'h4;
17'hf07:	data_out=16'h1;
17'hf08:	data_out=16'h8002;
17'hf09:	data_out=16'h8003;
17'hf0a:	data_out=16'h8002;
17'hf0b:	data_out=16'h8004;
17'hf0c:	data_out=16'h5;
17'hf0d:	data_out=16'h8005;
17'hf0e:	data_out=16'h8008;
17'hf0f:	data_out=16'h5;
17'hf10:	data_out=16'h8008;
17'hf11:	data_out=16'h3;
17'hf12:	data_out=16'h8002;
17'hf13:	data_out=16'h8007;
17'hf14:	data_out=16'h8005;
17'hf15:	data_out=16'h3;
17'hf16:	data_out=16'h8000;
17'hf17:	data_out=16'h7;
17'hf18:	data_out=16'h8003;
17'hf19:	data_out=16'h4;
17'hf1a:	data_out=16'h8005;
17'hf1b:	data_out=16'h6;
17'hf1c:	data_out=16'h8008;
17'hf1d:	data_out=16'h8001;
17'hf1e:	data_out=16'h3;
17'hf1f:	data_out=16'h8006;
17'hf20:	data_out=16'h4;
17'hf21:	data_out=16'h1;
17'hf22:	data_out=16'h8005;
17'hf23:	data_out=16'h7;
17'hf24:	data_out=16'h7;
17'hf25:	data_out=16'h8;
17'hf26:	data_out=16'h8001;
17'hf27:	data_out=16'h8004;
17'hf28:	data_out=16'h8004;
17'hf29:	data_out=16'h6;
17'hf2a:	data_out=16'h2;
17'hf2b:	data_out=16'h8008;
17'hf2c:	data_out=16'h8008;
17'hf2d:	data_out=16'h3;
17'hf2e:	data_out=16'h6;
17'hf2f:	data_out=16'h8007;
17'hf30:	data_out=16'h8004;
17'hf31:	data_out=16'h8005;
17'hf32:	data_out=16'h8005;
17'hf33:	data_out=16'h0;
17'hf34:	data_out=16'h7;
17'hf35:	data_out=16'h3;
17'hf36:	data_out=16'h8002;
17'hf37:	data_out=16'h8005;
17'hf38:	data_out=16'h8002;
17'hf39:	data_out=16'h1;
17'hf3a:	data_out=16'h8007;
17'hf3b:	data_out=16'h8001;
17'hf3c:	data_out=16'h8009;
17'hf3d:	data_out=16'h4;
17'hf3e:	data_out=16'h2;
17'hf3f:	data_out=16'h5;
17'hf40:	data_out=16'h8004;
17'hf41:	data_out=16'h7;
17'hf42:	data_out=16'h3;
17'hf43:	data_out=16'h8005;
17'hf44:	data_out=16'h6;
17'hf45:	data_out=16'h8007;
17'hf46:	data_out=16'h0;
17'hf47:	data_out=16'h8008;
17'hf48:	data_out=16'h8;
17'hf49:	data_out=16'h8007;
17'hf4a:	data_out=16'h8007;
17'hf4b:	data_out=16'h9;
17'hf4c:	data_out=16'h4;
17'hf4d:	data_out=16'h9;
17'hf4e:	data_out=16'h8008;
17'hf4f:	data_out=16'h8008;
17'hf50:	data_out=16'h8006;
17'hf51:	data_out=16'h8004;
17'hf52:	data_out=16'h1;
17'hf53:	data_out=16'h8008;
17'hf54:	data_out=16'h9;
17'hf55:	data_out=16'h8;
17'hf56:	data_out=16'h8003;
17'hf57:	data_out=16'h8002;
17'hf58:	data_out=16'h8000;
17'hf59:	data_out=16'h8001;
17'hf5a:	data_out=16'h6;
17'hf5b:	data_out=16'h1;
17'hf5c:	data_out=16'h8006;
17'hf5d:	data_out=16'h8001;
17'hf5e:	data_out=16'h8004;
17'hf5f:	data_out=16'h8000;
17'hf60:	data_out=16'h8003;
17'hf61:	data_out=16'h8;
17'hf62:	data_out=16'h4;
17'hf63:	data_out=16'h8007;
17'hf64:	data_out=16'h8008;
17'hf65:	data_out=16'h8005;
17'hf66:	data_out=16'h8005;
17'hf67:	data_out=16'h9;
17'hf68:	data_out=16'h8004;
17'hf69:	data_out=16'h8003;
17'hf6a:	data_out=16'h8;
17'hf6b:	data_out=16'h8009;
17'hf6c:	data_out=16'h8003;
17'hf6d:	data_out=16'h8008;
17'hf6e:	data_out=16'h8008;
17'hf6f:	data_out=16'h0;
17'hf70:	data_out=16'h8003;
17'hf71:	data_out=16'h2;
17'hf72:	data_out=16'h2;
17'hf73:	data_out=16'h8003;
17'hf74:	data_out=16'h0;
17'hf75:	data_out=16'h8;
17'hf76:	data_out=16'h4;
17'hf77:	data_out=16'h8009;
17'hf78:	data_out=16'h8003;
17'hf79:	data_out=16'h1;
17'hf7a:	data_out=16'h1;
17'hf7b:	data_out=16'h1;
17'hf7c:	data_out=16'h8009;
17'hf7d:	data_out=16'h6;
17'hf7e:	data_out=16'h8009;
17'hf7f:	data_out=16'h8003;
17'hf80:	data_out=16'h5;
17'hf81:	data_out=16'h4;
17'hf82:	data_out=16'h8001;
17'hf83:	data_out=16'h6;
17'hf84:	data_out=16'h8;
17'hf85:	data_out=16'h3;
17'hf86:	data_out=16'h6;
17'hf87:	data_out=16'h8005;
17'hf88:	data_out=16'h8009;
17'hf89:	data_out=16'h6;
17'hf8a:	data_out=16'h8005;
17'hf8b:	data_out=16'h8003;
17'hf8c:	data_out=16'h6;
17'hf8d:	data_out=16'h8003;
17'hf8e:	data_out=16'h6;
17'hf8f:	data_out=16'h8006;
17'hf90:	data_out=16'h8;
17'hf91:	data_out=16'h8001;
17'hf92:	data_out=16'h8000;
17'hf93:	data_out=16'h8001;
17'hf94:	data_out=16'h8003;
17'hf95:	data_out=16'h8006;
17'hf96:	data_out=16'h8001;
17'hf97:	data_out=16'h4;
17'hf98:	data_out=16'h4;
17'hf99:	data_out=16'h8009;
17'hf9a:	data_out=16'h8005;
17'hf9b:	data_out=16'h4;
17'hf9c:	data_out=16'h7;
17'hf9d:	data_out=16'h8004;
17'hf9e:	data_out=16'h8008;
17'hf9f:	data_out=16'h3;
17'hfa0:	data_out=16'h9;
17'hfa1:	data_out=16'h0;
17'hfa2:	data_out=16'h0;
17'hfa3:	data_out=16'h7;
17'hfa4:	data_out=16'h8006;
17'hfa5:	data_out=16'h8003;
17'hfa6:	data_out=16'h8007;
17'hfa7:	data_out=16'h8006;
17'hfa8:	data_out=16'h8006;
17'hfa9:	data_out=16'h8003;
17'hfaa:	data_out=16'h0;
17'hfab:	data_out=16'h9;
17'hfac:	data_out=16'h3;
17'hfad:	data_out=16'h8003;
17'hfae:	data_out=16'h8006;
17'hfaf:	data_out=16'h2;
17'hfb0:	data_out=16'h5;
17'hfb1:	data_out=16'h3;
17'hfb2:	data_out=16'h8008;
17'hfb3:	data_out=16'h8007;
17'hfb4:	data_out=16'h6;
17'hfb5:	data_out=16'h1;
17'hfb6:	data_out=16'h6;
17'hfb7:	data_out=16'h1;
17'hfb8:	data_out=16'h1;
17'hfb9:	data_out=16'h8008;
17'hfba:	data_out=16'h8004;
17'hfbb:	data_out=16'h8001;
17'hfbc:	data_out=16'h8003;
17'hfbd:	data_out=16'h8003;
17'hfbe:	data_out=16'h8008;
17'hfbf:	data_out=16'h8004;
17'hfc0:	data_out=16'h7;
17'hfc1:	data_out=16'h1;
17'hfc2:	data_out=16'h8006;
17'hfc3:	data_out=16'h8008;
17'hfc4:	data_out=16'h8;
17'hfc5:	data_out=16'h8004;
17'hfc6:	data_out=16'h8005;
17'hfc7:	data_out=16'h8008;
17'hfc8:	data_out=16'h3;
17'hfc9:	data_out=16'h5;
17'hfca:	data_out=16'h8008;
17'hfcb:	data_out=16'h8003;
17'hfcc:	data_out=16'h8007;
17'hfcd:	data_out=16'h8005;
17'hfce:	data_out=16'h8;
17'hfcf:	data_out=16'h7;
17'hfd0:	data_out=16'h7;
17'hfd1:	data_out=16'h8009;
17'hfd2:	data_out=16'h9;
17'hfd3:	data_out=16'h4;
17'hfd4:	data_out=16'h1;
17'hfd5:	data_out=16'h6;
17'hfd6:	data_out=16'h8004;
17'hfd7:	data_out=16'h8007;
17'hfd8:	data_out=16'h7;
17'hfd9:	data_out=16'h1;
17'hfda:	data_out=16'h0;
17'hfdb:	data_out=16'h8006;
17'hfdc:	data_out=16'h8;
17'hfdd:	data_out=16'h2;
17'hfde:	data_out=16'h8000;
17'hfdf:	data_out=16'h6;
17'hfe0:	data_out=16'h8006;
17'hfe1:	data_out=16'h3;
17'hfe2:	data_out=16'h7;
17'hfe3:	data_out=16'h8007;
17'hfe4:	data_out=16'h9;
17'hfe5:	data_out=16'h8007;
17'hfe6:	data_out=16'h8006;
17'hfe7:	data_out=16'h2;
17'hfe8:	data_out=16'h7;
17'hfe9:	data_out=16'h8005;
17'hfea:	data_out=16'h9;
17'hfeb:	data_out=16'h9;
17'hfec:	data_out=16'h8001;
17'hfed:	data_out=16'h8;
17'hfee:	data_out=16'h7;
17'hfef:	data_out=16'h8003;
17'hff0:	data_out=16'h8;
17'hff1:	data_out=16'h7;
17'hff2:	data_out=16'h8008;
17'hff3:	data_out=16'h8000;
17'hff4:	data_out=16'h3;
17'hff5:	data_out=16'h8003;
17'hff6:	data_out=16'h2;
17'hff7:	data_out=16'h1;
17'hff8:	data_out=16'h7;
17'hff9:	data_out=16'h8007;
17'hffa:	data_out=16'h4;
17'hffb:	data_out=16'h6;
17'hffc:	data_out=16'h4;
17'hffd:	data_out=16'h8005;
17'hffe:	data_out=16'h3;
17'hfff:	data_out=16'h7;
17'h1000:	data_out=16'h8;
17'h1001:	data_out=16'h2;
17'h1002:	data_out=16'ha;
17'h1003:	data_out=16'ha;
17'h1004:	data_out=16'h5;
17'h1005:	data_out=16'h8003;
17'h1006:	data_out=16'h1;
17'h1007:	data_out=16'h1;
17'h1008:	data_out=16'h8001;
17'h1009:	data_out=16'h8000;
17'h100a:	data_out=16'h3;
17'h100b:	data_out=16'ha;
17'h100c:	data_out=16'h2;
17'h100d:	data_out=16'h0;
17'h100e:	data_out=16'h8005;
17'h100f:	data_out=16'h8001;
17'h1010:	data_out=16'h8003;
17'h1011:	data_out=16'h8001;
17'h1012:	data_out=16'h7;
17'h1013:	data_out=16'hb;
17'h1014:	data_out=16'h2;
17'h1015:	data_out=16'h0;
17'h1016:	data_out=16'h1;
17'h1017:	data_out=16'h1;
17'h1018:	data_out=16'h1;
17'h1019:	data_out=16'h8003;
17'h101a:	data_out=16'h8001;
17'h101b:	data_out=16'h8002;
17'h101c:	data_out=16'h2;
17'h101d:	data_out=16'ha;
17'h101e:	data_out=16'h8004;
17'h101f:	data_out=16'h8002;
17'h1020:	data_out=16'h1;
17'h1021:	data_out=16'h8005;
17'h1022:	data_out=16'h8004;
17'h1023:	data_out=16'h8007;
17'h1024:	data_out=16'h8002;
17'h1025:	data_out=16'h7;
17'h1026:	data_out=16'h4;
17'h1027:	data_out=16'h8;
17'h1028:	data_out=16'h8003;
17'h1029:	data_out=16'h8004;
17'h102a:	data_out=16'h4;
17'h102b:	data_out=16'h5;
17'h102c:	data_out=16'h5;
17'h102d:	data_out=16'h9;
17'h102e:	data_out=16'h8006;
17'h102f:	data_out=16'h9;
17'h1030:	data_out=16'h8002;
17'h1031:	data_out=16'h8006;
17'h1032:	data_out=16'hc;
17'h1033:	data_out=16'h4;
17'h1034:	data_out=16'h1;
17'h1035:	data_out=16'h2;
17'h1036:	data_out=16'h8005;
17'h1037:	data_out=16'h8006;
17'h1038:	data_out=16'h3;
17'h1039:	data_out=16'h8001;
17'h103a:	data_out=16'h8002;
17'h103b:	data_out=16'h8005;
17'h103c:	data_out=16'h8000;
17'h103d:	data_out=16'h4;
17'h103e:	data_out=16'h8000;
17'h103f:	data_out=16'ha;
17'h1040:	data_out=16'h6;
17'h1041:	data_out=16'h7;
17'h1042:	data_out=16'ha;
17'h1043:	data_out=16'h8004;
17'h1044:	data_out=16'h4;
17'h1045:	data_out=16'h2;
17'h1046:	data_out=16'h8007;
17'h1047:	data_out=16'h6;
17'h1048:	data_out=16'h5;
17'h1049:	data_out=16'h4;
17'h104a:	data_out=16'h4;
17'h104b:	data_out=16'h0;
17'h104c:	data_out=16'h2;
17'h104d:	data_out=16'h5;
17'h104e:	data_out=16'h8001;
17'h104f:	data_out=16'h4;
17'h1050:	data_out=16'h4;
17'h1051:	data_out=16'h8004;
17'h1052:	data_out=16'h8003;
17'h1053:	data_out=16'h8001;
17'h1054:	data_out=16'h2;
17'h1055:	data_out=16'h1;
17'h1056:	data_out=16'h8002;
17'h1057:	data_out=16'h8007;
17'h1058:	data_out=16'h9;
17'h1059:	data_out=16'h5;
17'h105a:	data_out=16'h8004;
17'h105b:	data_out=16'h8002;
17'h105c:	data_out=16'h0;
17'h105d:	data_out=16'h4;
17'h105e:	data_out=16'h8006;
17'h105f:	data_out=16'h8005;
17'h1060:	data_out=16'h8001;
17'h1061:	data_out=16'hc;
17'h1062:	data_out=16'h1;
17'h1063:	data_out=16'h9;
17'h1064:	data_out=16'h2;
17'h1065:	data_out=16'h2;
17'h1066:	data_out=16'h7;
17'h1067:	data_out=16'h8003;
17'h1068:	data_out=16'h8005;
17'h1069:	data_out=16'h1;
17'h106a:	data_out=16'h5;
17'h106b:	data_out=16'h5;
17'h106c:	data_out=16'h8003;
17'h106d:	data_out=16'h8007;
17'h106e:	data_out=16'h8002;
17'h106f:	data_out=16'hb;
17'h1070:	data_out=16'h8005;
17'h1071:	data_out=16'h3;
17'h1072:	data_out=16'h8002;
17'h1073:	data_out=16'h7;
17'h1074:	data_out=16'h8002;
17'h1075:	data_out=16'h6;
17'h1076:	data_out=16'h6;
17'h1077:	data_out=16'h8007;
17'h1078:	data_out=16'h8003;
17'h1079:	data_out=16'h8008;
17'h107a:	data_out=16'h8004;
17'h107b:	data_out=16'h4;
17'h107c:	data_out=16'h3;
17'h107d:	data_out=16'h8004;
17'h107e:	data_out=16'h8;
17'h107f:	data_out=16'h8007;
17'h1080:	data_out=16'h800d;
17'h1081:	data_out=16'h8007;
17'h1082:	data_out=16'h8010;
17'h1083:	data_out=16'h6;
17'h1084:	data_out=16'h16;
17'h1085:	data_out=16'he;
17'h1086:	data_out=16'h8007;
17'h1087:	data_out=16'h8009;
17'h1088:	data_out=16'h800b;
17'h1089:	data_out=16'h4;
17'h108a:	data_out=16'h4;
17'h108b:	data_out=16'h8;
17'h108c:	data_out=16'h17;
17'h108d:	data_out=16'h8005;
17'h108e:	data_out=16'h8001;
17'h108f:	data_out=16'h800e;
17'h1090:	data_out=16'h5;
17'h1091:	data_out=16'he;
17'h1092:	data_out=16'h1;
17'h1093:	data_out=16'h8006;
17'h1094:	data_out=16'h800e;
17'h1095:	data_out=16'h2;
17'h1096:	data_out=16'h8009;
17'h1097:	data_out=16'h8007;
17'h1098:	data_out=16'h8001;
17'h1099:	data_out=16'h2;
17'h109a:	data_out=16'he;
17'h109b:	data_out=16'h8006;
17'h109c:	data_out=16'h8003;
17'h109d:	data_out=16'h800a;
17'h109e:	data_out=16'h800b;
17'h109f:	data_out=16'h8001;
17'h10a0:	data_out=16'h8002;
17'h10a1:	data_out=16'h8001;
17'h10a2:	data_out=16'h0;
17'h10a3:	data_out=16'h8004;
17'h10a4:	data_out=16'h8008;
17'h10a5:	data_out=16'h7;
17'h10a6:	data_out=16'h8007;
17'h10a7:	data_out=16'h8003;
17'h10a8:	data_out=16'h0;
17'h10a9:	data_out=16'h8007;
17'h10aa:	data_out=16'h8010;
17'h10ab:	data_out=16'h8002;
17'h10ac:	data_out=16'h4;
17'h10ad:	data_out=16'h8;
17'h10ae:	data_out=16'h8004;
17'h10af:	data_out=16'h8001;
17'h10b0:	data_out=16'h17;
17'h10b1:	data_out=16'h8001;
17'h10b2:	data_out=16'h1b;
17'h10b3:	data_out=16'h800c;
17'h10b4:	data_out=16'h800a;
17'h10b5:	data_out=16'hf;
17'h10b6:	data_out=16'h4;
17'h10b7:	data_out=16'h2;
17'h10b8:	data_out=16'h8006;
17'h10b9:	data_out=16'h8011;
17'h10ba:	data_out=16'h8009;
17'h10bb:	data_out=16'h8000;
17'h10bc:	data_out=16'h8006;
17'h10bd:	data_out=16'h2;
17'h10be:	data_out=16'h8;
17'h10bf:	data_out=16'h19;
17'h10c0:	data_out=16'h1;
17'h10c1:	data_out=16'h8002;
17'h10c2:	data_out=16'hb;
17'h10c3:	data_out=16'h5;
17'h10c4:	data_out=16'h8002;
17'h10c5:	data_out=16'h800d;
17'h10c6:	data_out=16'h800a;
17'h10c7:	data_out=16'h8002;
17'h10c8:	data_out=16'h8005;
17'h10c9:	data_out=16'h8002;
17'h10ca:	data_out=16'h8001;
17'h10cb:	data_out=16'h12;
17'h10cc:	data_out=16'hb;
17'h10cd:	data_out=16'h2;
17'h10ce:	data_out=16'h8003;
17'h10cf:	data_out=16'he;
17'h10d0:	data_out=16'h8006;
17'h10d1:	data_out=16'h8001;
17'h10d2:	data_out=16'h8006;
17'h10d3:	data_out=16'h8005;
17'h10d4:	data_out=16'h800a;
17'h10d5:	data_out=16'h800a;
17'h10d6:	data_out=16'h800a;
17'h10d7:	data_out=16'h8003;
17'h10d8:	data_out=16'h8006;
17'h10d9:	data_out=16'h4;
17'h10da:	data_out=16'h2;
17'h10db:	data_out=16'h4;
17'h10dc:	data_out=16'h8002;
17'h10dd:	data_out=16'h8;
17'h10de:	data_out=16'hc;
17'h10df:	data_out=16'h8001;
17'h10e0:	data_out=16'h8008;
17'h10e1:	data_out=16'h4;
17'h10e2:	data_out=16'h800c;
17'h10e3:	data_out=16'h800a;
17'h10e4:	data_out=16'h8007;
17'h10e5:	data_out=16'h9;
17'h10e6:	data_out=16'h8001;
17'h10e7:	data_out=16'h1;
17'h10e8:	data_out=16'h3;
17'h10e9:	data_out=16'h800a;
17'h10ea:	data_out=16'h2;
17'h10eb:	data_out=16'h5;
17'h10ec:	data_out=16'h2;
17'h10ed:	data_out=16'h8002;
17'h10ee:	data_out=16'h8003;
17'h10ef:	data_out=16'h16;
17'h10f0:	data_out=16'h2;
17'h10f1:	data_out=16'h8007;
17'h10f2:	data_out=16'h3;
17'h10f3:	data_out=16'h9;
17'h10f4:	data_out=16'h14;
17'h10f5:	data_out=16'h8;
17'h10f6:	data_out=16'h8004;
17'h10f7:	data_out=16'ha;
17'h10f8:	data_out=16'h8007;
17'h10f9:	data_out=16'h8009;
17'h10fa:	data_out=16'h8009;
17'h10fb:	data_out=16'h8001;
17'h10fc:	data_out=16'h8008;
17'h10fd:	data_out=16'h8004;
17'h10fe:	data_out=16'h800a;
17'h10ff:	data_out=16'h9;
17'h1100:	data_out=16'h825e;
17'h1101:	data_out=16'h82bd;
17'h1102:	data_out=16'h82a3;
17'h1103:	data_out=16'h8186;
17'h1104:	data_out=16'h234;
17'h1105:	data_out=16'h10;
17'h1106:	data_out=16'h80bf;
17'h1107:	data_out=16'h80ac;
17'h1108:	data_out=16'h8302;
17'h1109:	data_out=16'h80b2;
17'h110a:	data_out=16'h8212;
17'h110b:	data_out=16'h80ef;
17'h110c:	data_out=16'h275;
17'h110d:	data_out=16'h81a3;
17'h110e:	data_out=16'h8088;
17'h110f:	data_out=16'h82d6;
17'h1110:	data_out=16'h80e4;
17'h1111:	data_out=16'h9d;
17'h1112:	data_out=16'h8229;
17'h1113:	data_out=16'h812c;
17'h1114:	data_out=16'h8396;
17'h1115:	data_out=16'h813e;
17'h1116:	data_out=16'h8165;
17'h1117:	data_out=16'h8372;
17'h1118:	data_out=16'h8103;
17'h1119:	data_out=16'h105;
17'h111a:	data_out=16'h30f;
17'h111b:	data_out=16'h8250;
17'h111c:	data_out=16'h82a7;
17'h111d:	data_out=16'h82e1;
17'h111e:	data_out=16'h8395;
17'h111f:	data_out=16'h81d9;
17'h1120:	data_out=16'h81d9;
17'h1121:	data_out=16'h8077;
17'h1122:	data_out=16'h809e;
17'h1123:	data_out=16'h8160;
17'h1124:	data_out=16'h8160;
17'h1125:	data_out=16'h4b;
17'h1126:	data_out=16'h82b2;
17'h1127:	data_out=16'h82ea;
17'h1128:	data_out=16'h807f;
17'h1129:	data_out=16'h8206;
17'h112a:	data_out=16'h82c5;
17'h112b:	data_out=16'h810f;
17'h112c:	data_out=16'h810d;
17'h112d:	data_out=16'hec;
17'h112e:	data_out=16'h8227;
17'h112f:	data_out=16'h813c;
17'h1130:	data_out=16'h368;
17'h1131:	data_out=16'h8230;
17'h1132:	data_out=16'h36d;
17'h1133:	data_out=16'h83a3;
17'h1134:	data_out=16'h81e4;
17'h1135:	data_out=16'h194;
17'h1136:	data_out=16'h8242;
17'h1137:	data_out=16'h82a6;
17'h1138:	data_out=16'h832c;
17'h1139:	data_out=16'h837a;
17'h113a:	data_out=16'h8149;
17'h113b:	data_out=16'h8013;
17'h113c:	data_out=16'h82ca;
17'h113d:	data_out=16'h816c;
17'h113e:	data_out=16'h8080;
17'h113f:	data_out=16'h13c;
17'h1140:	data_out=16'h162;
17'h1141:	data_out=16'h81de;
17'h1142:	data_out=16'h23b;
17'h1143:	data_out=16'h806c;
17'h1144:	data_out=16'h8062;
17'h1145:	data_out=16'h8170;
17'h1146:	data_out=16'h81e5;
17'h1147:	data_out=16'h80d8;
17'h1148:	data_out=16'h80d4;
17'h1149:	data_out=16'h26;
17'h114a:	data_out=16'ha3;
17'h114b:	data_out=16'h1ba;
17'h114c:	data_out=16'hb2;
17'h114d:	data_out=16'h80c9;
17'h114e:	data_out=16'h816b;
17'h114f:	data_out=16'hbd;
17'h1150:	data_out=16'h3e;
17'h1151:	data_out=16'h82d8;
17'h1152:	data_out=16'h814d;
17'h1153:	data_out=16'h82b6;
17'h1154:	data_out=16'h81e8;
17'h1155:	data_out=16'h834c;
17'h1156:	data_out=16'h8234;
17'h1157:	data_out=16'h820a;
17'h1158:	data_out=16'h82f4;
17'h1159:	data_out=16'h2d;
17'h115a:	data_out=16'h8340;
17'h115b:	data_out=16'h82f3;
17'h115c:	data_out=16'h812c;
17'h115d:	data_out=16'h810b;
17'h115e:	data_out=16'h8021;
17'h115f:	data_out=16'h80f3;
17'h1160:	data_out=16'h8251;
17'h1161:	data_out=16'h8156;
17'h1162:	data_out=16'h836f;
17'h1163:	data_out=16'h836c;
17'h1164:	data_out=16'h8231;
17'h1165:	data_out=16'h1a9;
17'h1166:	data_out=16'h109;
17'h1167:	data_out=16'h8151;
17'h1168:	data_out=16'h8085;
17'h1169:	data_out=16'h82b1;
17'h116a:	data_out=16'h8089;
17'h116b:	data_out=16'h165;
17'h116c:	data_out=16'h8261;
17'h116d:	data_out=16'h839b;
17'h116e:	data_out=16'h8084;
17'h116f:	data_out=16'h19d;
17'h1170:	data_out=16'h8087;
17'h1171:	data_out=16'h8315;
17'h1172:	data_out=16'h802a;
17'h1173:	data_out=16'h8065;
17'h1174:	data_out=16'h36e;
17'h1175:	data_out=16'h8154;
17'h1176:	data_out=16'h815d;
17'h1177:	data_out=16'h119;
17'h1178:	data_out=16'h8051;
17'h1179:	data_out=16'h82f8;
17'h117a:	data_out=16'h839a;
17'h117b:	data_out=16'h807d;
17'h117c:	data_out=16'h8185;
17'h117d:	data_out=16'h8149;
17'h117e:	data_out=16'h80d2;
17'h117f:	data_out=16'h1e;
17'h1180:	data_out=16'h8381;
17'h1181:	data_out=16'h83f2;
17'h1182:	data_out=16'h83b7;
17'h1183:	data_out=16'h81f1;
17'h1184:	data_out=16'h4c8;
17'h1185:	data_out=16'h11d;
17'h1186:	data_out=16'h8089;
17'h1187:	data_out=16'h8069;
17'h1188:	data_out=16'h849a;
17'h1189:	data_out=16'h8181;
17'h118a:	data_out=16'h83ae;
17'h118b:	data_out=16'h8181;
17'h118c:	data_out=16'h4a8;
17'h118d:	data_out=16'h8301;
17'h118e:	data_out=16'h80ee;
17'h118f:	data_out=16'h8434;
17'h1190:	data_out=16'h80d8;
17'h1191:	data_out=16'h1be;
17'h1192:	data_out=16'h8321;
17'h1193:	data_out=16'h81f1;
17'h1194:	data_out=16'h85fd;
17'h1195:	data_out=16'h81c5;
17'h1196:	data_out=16'h8214;
17'h1197:	data_out=16'h8589;
17'h1198:	data_out=16'h8205;
17'h1199:	data_out=16'h243;
17'h119a:	data_out=16'h646;
17'h119b:	data_out=16'h8405;
17'h119c:	data_out=16'h8401;
17'h119d:	data_out=16'h845c;
17'h119e:	data_out=16'h85ec;
17'h119f:	data_out=16'h82ba;
17'h11a0:	data_out=16'h82df;
17'h11a1:	data_out=16'h80e2;
17'h11a2:	data_out=16'h80af;
17'h11a3:	data_out=16'h81cf;
17'h11a4:	data_out=16'h81cf;
17'h11a5:	data_out=16'hb4;
17'h11a6:	data_out=16'h84e7;
17'h11a7:	data_out=16'h846a;
17'h11a8:	data_out=16'h80e2;
17'h11a9:	data_out=16'h83cf;
17'h11aa:	data_out=16'h8499;
17'h11ab:	data_out=16'h8202;
17'h11ac:	data_out=16'h819b;
17'h11ad:	data_out=16'h1c1;
17'h11ae:	data_out=16'h83d1;
17'h11af:	data_out=16'h8111;
17'h11b0:	data_out=16'h618;
17'h11b1:	data_out=16'h83fe;
17'h11b2:	data_out=16'h62b;
17'h11b3:	data_out=16'h8641;
17'h11b4:	data_out=16'h836c;
17'h11b5:	data_out=16'h324;
17'h11b6:	data_out=16'h8322;
17'h11b7:	data_out=16'h83bf;
17'h11b8:	data_out=16'h8501;
17'h11b9:	data_out=16'h863e;
17'h11ba:	data_out=16'h81a7;
17'h11bb:	data_out=16'h67;
17'h11bc:	data_out=16'h83d9;
17'h11bd:	data_out=16'h8275;
17'h11be:	data_out=16'h80e3;
17'h11bf:	data_out=16'h29a;
17'h11c0:	data_out=16'h2a9;
17'h11c1:	data_out=16'h825c;
17'h11c2:	data_out=16'h41c;
17'h11c3:	data_out=16'h80c3;
17'h11c4:	data_out=16'h806f;
17'h11c5:	data_out=16'h81ca;
17'h11c6:	data_out=16'h824f;
17'h11c7:	data_out=16'h8145;
17'h11c8:	data_out=16'h819e;
17'h11c9:	data_out=16'h83;
17'h11ca:	data_out=16'h17d;
17'h11cb:	data_out=16'h335;
17'h11cc:	data_out=16'h171;
17'h11cd:	data_out=16'h80a7;
17'h11ce:	data_out=16'h8261;
17'h11cf:	data_out=16'h190;
17'h11d0:	data_out=16'h7e;
17'h11d1:	data_out=16'h842e;
17'h11d2:	data_out=16'h81a8;
17'h11d3:	data_out=16'h843a;
17'h11d4:	data_out=16'h82cc;
17'h11d5:	data_out=16'h8504;
17'h11d6:	data_out=16'h8333;
17'h11d7:	data_out=16'h82fe;
17'h11d8:	data_out=16'h843f;
17'h11d9:	data_out=16'h161;
17'h11da:	data_out=16'h8540;
17'h11db:	data_out=16'h846d;
17'h11dc:	data_out=16'h812e;
17'h11dd:	data_out=16'h8151;
17'h11de:	data_out=16'h2;
17'h11df:	data_out=16'h81d2;
17'h11e0:	data_out=16'h8430;
17'h11e1:	data_out=16'h8243;
17'h11e2:	data_out=16'h8567;
17'h11e3:	data_out=16'h8625;
17'h11e4:	data_out=16'h8422;
17'h11e5:	data_out=16'h395;
17'h11e6:	data_out=16'h23a;
17'h11e7:	data_out=16'h8203;
17'h11e8:	data_out=16'h80ec;
17'h11e9:	data_out=16'h847a;
17'h11ea:	data_out=16'h80f4;
17'h11eb:	data_out=16'h330;
17'h11ec:	data_out=16'h830e;
17'h11ed:	data_out=16'h8626;
17'h11ee:	data_out=16'h80ee;
17'h11ef:	data_out=16'h3d4;
17'h11f0:	data_out=16'h80f9;
17'h11f1:	data_out=16'h85f3;
17'h11f2:	data_out=16'h45;
17'h11f3:	data_out=16'h3d;
17'h11f4:	data_out=16'h623;
17'h11f5:	data_out=16'h8237;
17'h11f6:	data_out=16'h8260;
17'h11f7:	data_out=16'h1c1;
17'h11f8:	data_out=16'h8079;
17'h11f9:	data_out=16'h8581;
17'h11fa:	data_out=16'h85ff;
17'h11fb:	data_out=16'h80dd;
17'h11fc:	data_out=16'h8211;
17'h11fd:	data_out=16'h81a1;
17'h11fe:	data_out=16'h8173;
17'h11ff:	data_out=16'h6a;
17'h1200:	data_out=16'h84dc;
17'h1201:	data_out=16'h848d;
17'h1202:	data_out=16'h82ea;
17'h1203:	data_out=16'h81aa;
17'h1204:	data_out=16'h5cc;
17'h1205:	data_out=16'h193;
17'h1206:	data_out=16'h8017;
17'h1207:	data_out=16'h8035;
17'h1208:	data_out=16'h83b8;
17'h1209:	data_out=16'h81a5;
17'h120a:	data_out=16'h8386;
17'h120b:	data_out=16'h8071;
17'h120c:	data_out=16'h5d0;
17'h120d:	data_out=16'h81c4;
17'h120e:	data_out=16'h8092;
17'h120f:	data_out=16'h8333;
17'h1210:	data_out=16'h809f;
17'h1211:	data_out=16'h1cd;
17'h1212:	data_out=16'h829a;
17'h1213:	data_out=16'h80a8;
17'h1214:	data_out=16'h861c;
17'h1215:	data_out=16'h81e1;
17'h1216:	data_out=16'h819e;
17'h1217:	data_out=16'h8536;
17'h1218:	data_out=16'h818f;
17'h1219:	data_out=16'h22b;
17'h121a:	data_out=16'h75f;
17'h121b:	data_out=16'h8325;
17'h121c:	data_out=16'h84e3;
17'h121d:	data_out=16'h852c;
17'h121e:	data_out=16'h8603;
17'h121f:	data_out=16'h8216;
17'h1220:	data_out=16'h8415;
17'h1221:	data_out=16'h808d;
17'h1222:	data_out=16'h806d;
17'h1223:	data_out=16'h8192;
17'h1224:	data_out=16'h8192;
17'h1225:	data_out=16'h123;
17'h1226:	data_out=16'h83e7;
17'h1227:	data_out=16'h856e;
17'h1228:	data_out=16'h8088;
17'h1229:	data_out=16'h83a8;
17'h122a:	data_out=16'h82fa;
17'h122b:	data_out=16'h8213;
17'h122c:	data_out=16'h8099;
17'h122d:	data_out=16'h1cc;
17'h122e:	data_out=16'h824c;
17'h122f:	data_out=16'h8113;
17'h1230:	data_out=16'h711;
17'h1231:	data_out=16'h853a;
17'h1232:	data_out=16'h73c;
17'h1233:	data_out=16'h86c2;
17'h1234:	data_out=16'h84db;
17'h1235:	data_out=16'h3a5;
17'h1236:	data_out=16'h8299;
17'h1237:	data_out=16'h82ef;
17'h1238:	data_out=16'h8696;
17'h1239:	data_out=16'h86bd;
17'h123a:	data_out=16'h8184;
17'h123b:	data_out=16'h9e;
17'h123c:	data_out=16'h830a;
17'h123d:	data_out=16'h83e8;
17'h123e:	data_out=16'h8088;
17'h123f:	data_out=16'h2a2;
17'h1240:	data_out=16'h288;
17'h1241:	data_out=16'h8197;
17'h1242:	data_out=16'h547;
17'h1243:	data_out=16'h67;
17'h1244:	data_out=16'h812a;
17'h1245:	data_out=16'h81e1;
17'h1246:	data_out=16'h81ac;
17'h1247:	data_out=16'h8115;
17'h1248:	data_out=16'h8051;
17'h1249:	data_out=16'hed;
17'h124a:	data_out=16'h23e;
17'h124b:	data_out=16'h4cf;
17'h124c:	data_out=16'h1bf;
17'h124d:	data_out=16'h80ba;
17'h124e:	data_out=16'h8099;
17'h124f:	data_out=16'h1ba;
17'h1250:	data_out=16'hf9;
17'h1251:	data_out=16'h8335;
17'h1252:	data_out=16'h8171;
17'h1253:	data_out=16'h8428;
17'h1254:	data_out=16'h835f;
17'h1255:	data_out=16'h83ff;
17'h1256:	data_out=16'h8316;
17'h1257:	data_out=16'h82d6;
17'h1258:	data_out=16'h8355;
17'h1259:	data_out=16'h139;
17'h125a:	data_out=16'h84a9;
17'h125b:	data_out=16'h853d;
17'h125c:	data_out=16'h8191;
17'h125d:	data_out=16'h806f;
17'h125e:	data_out=16'haf;
17'h125f:	data_out=16'h816d;
17'h1260:	data_out=16'h83aa;
17'h1261:	data_out=16'h8270;
17'h1262:	data_out=16'h8472;
17'h1263:	data_out=16'h863d;
17'h1264:	data_out=16'h85d3;
17'h1265:	data_out=16'h416;
17'h1266:	data_out=16'h248;
17'h1267:	data_out=16'h815d;
17'h1268:	data_out=16'h8086;
17'h1269:	data_out=16'h8385;
17'h126a:	data_out=16'h809c;
17'h126b:	data_out=16'h438;
17'h126c:	data_out=16'h8329;
17'h126d:	data_out=16'h86a1;
17'h126e:	data_out=16'h809b;
17'h126f:	data_out=16'h557;
17'h1270:	data_out=16'h80a1;
17'h1271:	data_out=16'h8489;
17'h1272:	data_out=16'h67;
17'h1273:	data_out=16'h8011;
17'h1274:	data_out=16'h720;
17'h1275:	data_out=16'h8149;
17'h1276:	data_out=16'h822b;
17'h1277:	data_out=16'h276;
17'h1278:	data_out=16'h9e;
17'h1279:	data_out=16'h8369;
17'h127a:	data_out=16'h8626;
17'h127b:	data_out=16'h8079;
17'h127c:	data_out=16'h822c;
17'h127d:	data_out=16'h8169;
17'h127e:	data_out=16'h8161;
17'h127f:	data_out=16'hd6;
17'h1280:	data_out=16'h819d;
17'h1281:	data_out=16'h806f;
17'h1282:	data_out=16'h5c;
17'h1283:	data_out=16'h188;
17'h1284:	data_out=16'h49f;
17'h1285:	data_out=16'h3ab;
17'h1286:	data_out=16'h805d;
17'h1287:	data_out=16'h808f;
17'h1288:	data_out=16'hcf;
17'h1289:	data_out=16'h8193;
17'h128a:	data_out=16'hc3;
17'h128b:	data_out=16'h2a3;
17'h128c:	data_out=16'h4f8;
17'h128d:	data_out=16'h106;
17'h128e:	data_out=16'h21;
17'h128f:	data_out=16'h8051;
17'h1290:	data_out=16'hf;
17'h1291:	data_out=16'h264;
17'h1292:	data_out=16'h8051;
17'h1293:	data_out=16'h2a4;
17'h1294:	data_out=16'h8164;
17'h1295:	data_out=16'h80ca;
17'h1296:	data_out=16'hc6;
17'h1297:	data_out=16'h801f;
17'h1298:	data_out=16'h80df;
17'h1299:	data_out=16'h17a;
17'h129a:	data_out=16'h567;
17'h129b:	data_out=16'h155;
17'h129c:	data_out=16'h807b;
17'h129d:	data_out=16'h8074;
17'h129e:	data_out=16'h8182;
17'h129f:	data_out=16'h810c;
17'h12a0:	data_out=16'h8125;
17'h12a1:	data_out=16'h31;
17'h12a2:	data_out=16'h804d;
17'h12a3:	data_out=16'h8109;
17'h12a4:	data_out=16'h8109;
17'h12a5:	data_out=16'h189;
17'h12a6:	data_out=16'h61;
17'h12a7:	data_out=16'h80d3;
17'h12a8:	data_out=16'h30;
17'h12a9:	data_out=16'h95;
17'h12aa:	data_out=16'h83;
17'h12ab:	data_out=16'h815e;
17'h12ac:	data_out=16'h1c8;
17'h12ad:	data_out=16'h33e;
17'h12ae:	data_out=16'h127;
17'h12af:	data_out=16'h10d;
17'h12b0:	data_out=16'h682;
17'h12b1:	data_out=16'h8075;
17'h12b2:	data_out=16'h687;
17'h12b3:	data_out=16'h8255;
17'h12b4:	data_out=16'h8142;
17'h12b5:	data_out=16'h532;
17'h12b6:	data_out=16'h2e;
17'h12b7:	data_out=16'h84;
17'h12b8:	data_out=16'h81f2;
17'h12b9:	data_out=16'h82c3;
17'h12ba:	data_out=16'h8179;
17'h12bb:	data_out=16'h27d;
17'h12bc:	data_out=16'h240;
17'h12bd:	data_out=16'h815c;
17'h12be:	data_out=16'h3a;
17'h12bf:	data_out=16'h407;
17'h12c0:	data_out=16'h1ce;
17'h12c1:	data_out=16'h1ca;
17'h12c2:	data_out=16'h422;
17'h12c3:	data_out=16'h13e;
17'h12c4:	data_out=16'h1c5;
17'h12c5:	data_out=16'h80bc;
17'h12c6:	data_out=16'h14a;
17'h12c7:	data_out=16'h811d;
17'h12c8:	data_out=16'h8b;
17'h12c9:	data_out=16'h120;
17'h12ca:	data_out=16'h282;
17'h12cb:	data_out=16'h470;
17'h12cc:	data_out=16'h1ab;
17'h12cd:	data_out=16'h80d7;
17'h12ce:	data_out=16'h283;
17'h12cf:	data_out=16'h15f;
17'h12d0:	data_out=16'hcb;
17'h12d1:	data_out=16'h124;
17'h12d2:	data_out=16'h80fa;
17'h12d3:	data_out=16'hd9;
17'h12d4:	data_out=16'h41;
17'h12d5:	data_out=16'hbb;
17'h12d6:	data_out=16'h80c6;
17'h12d7:	data_out=16'h8176;
17'h12d8:	data_out=16'h10c;
17'h12d9:	data_out=16'hc6;
17'h12da:	data_out=16'h101;
17'h12db:	data_out=16'h8057;
17'h12dc:	data_out=16'hf8;
17'h12dd:	data_out=16'h245;
17'h12de:	data_out=16'h2b9;
17'h12df:	data_out=16'h80f1;
17'h12e0:	data_out=16'hea;
17'h12e1:	data_out=16'h1bb;
17'h12e2:	data_out=16'h8028;
17'h12e3:	data_out=16'h818d;
17'h12e4:	data_out=16'h825e;
17'h12e5:	data_out=16'h2d0;
17'h12e6:	data_out=16'h15d;
17'h12e7:	data_out=16'h8012;
17'h12e8:	data_out=16'h35;
17'h12e9:	data_out=16'hda;
17'h12ea:	data_out=16'h1f;
17'h12eb:	data_out=16'h33e;
17'h12ec:	data_out=16'ha0;
17'h12ed:	data_out=16'h823e;
17'h12ee:	data_out=16'h26;
17'h12ef:	data_out=16'h4f1;
17'h12f0:	data_out=16'h2e;
17'h12f1:	data_out=16'h8175;
17'h12f2:	data_out=16'h341;
17'h12f3:	data_out=16'h21b;
17'h12f4:	data_out=16'h68f;
17'h12f5:	data_out=16'h40e;
17'h12f6:	data_out=16'h816d;
17'h12f7:	data_out=16'h2c1;
17'h12f8:	data_out=16'h123;
17'h12f9:	data_out=16'hed;
17'h12fa:	data_out=16'h8183;
17'h12fb:	data_out=16'h2f;
17'h12fc:	data_out=16'h81ae;
17'h12fd:	data_out=16'h80a4;
17'h12fe:	data_out=16'h80d8;
17'h12ff:	data_out=16'h155;
17'h1300:	data_out=16'h81cf;
17'h1301:	data_out=16'h8094;
17'h1302:	data_out=16'h80f1;
17'h1303:	data_out=16'h32e;
17'h1304:	data_out=16'h8f0;
17'h1305:	data_out=16'h6de;
17'h1306:	data_out=16'h8015;
17'h1307:	data_out=16'h5;
17'h1308:	data_out=16'h4e;
17'h1309:	data_out=16'h822e;
17'h130a:	data_out=16'hed;
17'h130b:	data_out=16'h1e3;
17'h130c:	data_out=16'h94e;
17'h130d:	data_out=16'hb1;
17'h130e:	data_out=16'h21;
17'h130f:	data_out=16'h8255;
17'h1310:	data_out=16'h101;
17'h1311:	data_out=16'h542;
17'h1312:	data_out=16'h820b;
17'h1313:	data_out=16'h348;
17'h1314:	data_out=16'h83e9;
17'h1315:	data_out=16'h80aa;
17'h1316:	data_out=16'h167;
17'h1317:	data_out=16'h8222;
17'h1318:	data_out=16'h826a;
17'h1319:	data_out=16'h2bf;
17'h131a:	data_out=16'ha00;
17'h131b:	data_out=16'h15;
17'h131c:	data_out=16'h8003;
17'h131d:	data_out=16'h80a6;
17'h131e:	data_out=16'h8429;
17'h131f:	data_out=16'h8299;
17'h1320:	data_out=16'h8102;
17'h1321:	data_out=16'h2a;
17'h1322:	data_out=16'h8052;
17'h1323:	data_out=16'h8116;
17'h1324:	data_out=16'h8115;
17'h1325:	data_out=16'h236;
17'h1326:	data_out=16'h8088;
17'h1327:	data_out=16'h80ee;
17'h1328:	data_out=16'h2d;
17'h1329:	data_out=16'h8125;
17'h132a:	data_out=16'h8213;
17'h132b:	data_out=16'h81c4;
17'h132c:	data_out=16'h286;
17'h132d:	data_out=16'h504;
17'h132e:	data_out=16'h8097;
17'h132f:	data_out=16'h299;
17'h1330:	data_out=16'ha00;
17'h1331:	data_out=16'h8066;
17'h1332:	data_out=16'ha00;
17'h1333:	data_out=16'h8561;
17'h1334:	data_out=16'h81ff;
17'h1335:	data_out=16'h973;
17'h1336:	data_out=16'h8138;
17'h1337:	data_out=16'h80f8;
17'h1338:	data_out=16'h8252;
17'h1339:	data_out=16'h85cb;
17'h133a:	data_out=16'h822b;
17'h133b:	data_out=16'h533;
17'h133c:	data_out=16'h2cb;
17'h133d:	data_out=16'h81b5;
17'h133e:	data_out=16'h31;
17'h133f:	data_out=16'h701;
17'h1340:	data_out=16'h4c3;
17'h1341:	data_out=16'h191;
17'h1342:	data_out=16'h675;
17'h1343:	data_out=16'h171;
17'h1344:	data_out=16'h1f2;
17'h1345:	data_out=16'h8096;
17'h1346:	data_out=16'h15b;
17'h1347:	data_out=16'h818b;
17'h1348:	data_out=16'h8050;
17'h1349:	data_out=16'h240;
17'h134a:	data_out=16'h3ae;
17'h134b:	data_out=16'h67e;
17'h134c:	data_out=16'h246;
17'h134d:	data_out=16'h8057;
17'h134e:	data_out=16'h106;
17'h134f:	data_out=16'h1b9;
17'h1350:	data_out=16'h2b5;
17'h1351:	data_out=16'he5;
17'h1352:	data_out=16'h80eb;
17'h1353:	data_out=16'hd6;
17'h1354:	data_out=16'he5;
17'h1355:	data_out=16'h8036;
17'h1356:	data_out=16'h81f8;
17'h1357:	data_out=16'h823f;
17'h1358:	data_out=16'h4e;
17'h1359:	data_out=16'h2a9;
17'h135a:	data_out=16'h4e;
17'h135b:	data_out=16'h802f;
17'h135c:	data_out=16'h221;
17'h135d:	data_out=16'h381;
17'h135e:	data_out=16'h415;
17'h135f:	data_out=16'h81cc;
17'h1360:	data_out=16'h8020;
17'h1361:	data_out=16'h2a7;
17'h1362:	data_out=16'h8243;
17'h1363:	data_out=16'h8405;
17'h1364:	data_out=16'h8386;
17'h1365:	data_out=16'h577;
17'h1366:	data_out=16'h273;
17'h1367:	data_out=16'h80ff;
17'h1368:	data_out=16'h33;
17'h1369:	data_out=16'hf;
17'h136a:	data_out=16'h800f;
17'h136b:	data_out=16'h6ea;
17'h136c:	data_out=16'h108;
17'h136d:	data_out=16'h8538;
17'h136e:	data_out=16'hf;
17'h136f:	data_out=16'ha00;
17'h1370:	data_out=16'h16;
17'h1371:	data_out=16'h85ce;
17'h1372:	data_out=16'h649;
17'h1373:	data_out=16'h4e4;
17'h1374:	data_out=16'ha00;
17'h1375:	data_out=16'h4c2;
17'h1376:	data_out=16'h8237;
17'h1377:	data_out=16'h3ec;
17'h1378:	data_out=16'h21a;
17'h1379:	data_out=16'h81cf;
17'h137a:	data_out=16'h8426;
17'h137b:	data_out=16'h30;
17'h137c:	data_out=16'h8287;
17'h137d:	data_out=16'h80b8;
17'h137e:	data_out=16'h80df;
17'h137f:	data_out=16'h2d2;
17'h1380:	data_out=16'h7b;
17'h1381:	data_out=16'h26f;
17'h1382:	data_out=16'h8d;
17'h1383:	data_out=16'h531;
17'h1384:	data_out=16'ha00;
17'h1385:	data_out=16'h9f7;
17'h1386:	data_out=16'h809d;
17'h1387:	data_out=16'h88;
17'h1388:	data_out=16'h2df;
17'h1389:	data_out=16'h8321;
17'h138a:	data_out=16'h4d0;
17'h138b:	data_out=16'h2cc;
17'h138c:	data_out=16'ha00;
17'h138d:	data_out=16'hf2;
17'h138e:	data_out=16'h4a;
17'h138f:	data_out=16'h8166;
17'h1390:	data_out=16'h180;
17'h1391:	data_out=16'h8b1;
17'h1392:	data_out=16'h831f;
17'h1393:	data_out=16'h4a7;
17'h1394:	data_out=16'h8405;
17'h1395:	data_out=16'h8006;
17'h1396:	data_out=16'h32e;
17'h1397:	data_out=16'h81af;
17'h1398:	data_out=16'h8338;
17'h1399:	data_out=16'h31c;
17'h139a:	data_out=16'ha00;
17'h139b:	data_out=16'h18d;
17'h139c:	data_out=16'h2e7;
17'h139d:	data_out=16'h292;
17'h139e:	data_out=16'h8397;
17'h139f:	data_out=16'h8359;
17'h13a0:	data_out=16'h2e;
17'h13a1:	data_out=16'h45;
17'h13a2:	data_out=16'h806a;
17'h13a3:	data_out=16'h80c6;
17'h13a4:	data_out=16'h80c4;
17'h13a5:	data_out=16'h27d;
17'h13a6:	data_out=16'h38;
17'h13a7:	data_out=16'h227;
17'h13a8:	data_out=16'h66;
17'h13a9:	data_out=16'h8015;
17'h13aa:	data_out=16'h816b;
17'h13ab:	data_out=16'h8053;
17'h13ac:	data_out=16'h3f5;
17'h13ad:	data_out=16'h706;
17'h13ae:	data_out=16'h80d3;
17'h13af:	data_out=16'h4e6;
17'h13b0:	data_out=16'ha00;
17'h13b1:	data_out=16'h2ce;
17'h13b2:	data_out=16'ha00;
17'h13b3:	data_out=16'h85b2;
17'h13b4:	data_out=16'h8d;
17'h13b5:	data_out=16'ha00;
17'h13b6:	data_out=16'h7a;
17'h13b7:	data_out=16'h81;
17'h13b8:	data_out=16'h803d;
17'h13b9:	data_out=16'h85d2;
17'h13ba:	data_out=16'h8361;
17'h13bb:	data_out=16'h898;
17'h13bc:	data_out=16'h64c;
17'h13bd:	data_out=16'h25;
17'h13be:	data_out=16'h6d;
17'h13bf:	data_out=16'h9f4;
17'h13c0:	data_out=16'h569;
17'h13c1:	data_out=16'h35d;
17'h13c2:	data_out=16'h857;
17'h13c3:	data_out=16'h75;
17'h13c4:	data_out=16'h4d1;
17'h13c5:	data_out=16'h1a;
17'h13c6:	data_out=16'h2d5;
17'h13c7:	data_out=16'h822b;
17'h13c8:	data_out=16'h819d;
17'h13c9:	data_out=16'h28e;
17'h13ca:	data_out=16'h519;
17'h13cb:	data_out=16'h917;
17'h13cc:	data_out=16'h282;
17'h13cd:	data_out=16'h806d;
17'h13ce:	data_out=16'h25a;
17'h13cf:	data_out=16'h1d7;
17'h13d0:	data_out=16'h2c2;
17'h13d1:	data_out=16'h319;
17'h13d2:	data_out=16'h8083;
17'h13d3:	data_out=16'h3cf;
17'h13d4:	data_out=16'h28b;
17'h13d5:	data_out=16'h1f6;
17'h13d6:	data_out=16'h8240;
17'h13d7:	data_out=16'h82cf;
17'h13d8:	data_out=16'h2c1;
17'h13d9:	data_out=16'h37d;
17'h13da:	data_out=16'h277;
17'h13db:	data_out=16'h31c;
17'h13dc:	data_out=16'h532;
17'h13dd:	data_out=16'h4d6;
17'h13de:	data_out=16'h638;
17'h13df:	data_out=16'h81f7;
17'h13e0:	data_out=16'h192;
17'h13e1:	data_out=16'h5de;
17'h13e2:	data_out=16'h8166;
17'h13e3:	data_out=16'h844a;
17'h13e4:	data_out=16'h825e;
17'h13e5:	data_out=16'h7d3;
17'h13e6:	data_out=16'h2b8;
17'h13e7:	data_out=16'h815d;
17'h13e8:	data_out=16'h5d;
17'h13e9:	data_out=16'h233;
17'h13ea:	data_out=16'h31;
17'h13eb:	data_out=16'h942;
17'h13ec:	data_out=16'h47f;
17'h13ed:	data_out=16'h8553;
17'h13ee:	data_out=16'h37;
17'h13ef:	data_out=16'ha00;
17'h13f0:	data_out=16'h3d;
17'h13f1:	data_out=16'h8760;
17'h13f2:	data_out=16'h957;
17'h13f3:	data_out=16'h841;
17'h13f4:	data_out=16'ha00;
17'h13f5:	data_out=16'h897;
17'h13f6:	data_out=16'h8218;
17'h13f7:	data_out=16'h43c;
17'h13f8:	data_out=16'h154;
17'h13f9:	data_out=16'h81ae;
17'h13fa:	data_out=16'h843e;
17'h13fb:	data_out=16'h69;
17'h13fc:	data_out=16'h82e3;
17'h13fd:	data_out=16'h819e;
17'h13fe:	data_out=16'h8142;
17'h13ff:	data_out=16'h335;
17'h1400:	data_out=16'h81a6;
17'h1401:	data_out=16'h8045;
17'h1402:	data_out=16'h83f6;
17'h1403:	data_out=16'h469;
17'h1404:	data_out=16'ha00;
17'h1405:	data_out=16'ha00;
17'h1406:	data_out=16'h80c6;
17'h1407:	data_out=16'h1f8;
17'h1408:	data_out=16'h816a;
17'h1409:	data_out=16'h83f8;
17'h140a:	data_out=16'h14a;
17'h140b:	data_out=16'h836e;
17'h140c:	data_out=16'ha00;
17'h140d:	data_out=16'h8321;
17'h140e:	data_out=16'h80f8;
17'h140f:	data_out=16'h86bd;
17'h1410:	data_out=16'h5a;
17'h1411:	data_out=16'h96a;
17'h1412:	data_out=16'h86f6;
17'h1413:	data_out=16'h2a8;
17'h1414:	data_out=16'h8a00;
17'h1415:	data_out=16'h80a4;
17'h1416:	data_out=16'h21a;
17'h1417:	data_out=16'h8847;
17'h1418:	data_out=16'h8503;
17'h1419:	data_out=16'h556;
17'h141a:	data_out=16'ha00;
17'h141b:	data_out=16'h8375;
17'h141c:	data_out=16'h65;
17'h141d:	data_out=16'h1a;
17'h141e:	data_out=16'h89d0;
17'h141f:	data_out=16'h856d;
17'h1420:	data_out=16'h816b;
17'h1421:	data_out=16'h80df;
17'h1422:	data_out=16'h19;
17'h1423:	data_out=16'h80c1;
17'h1424:	data_out=16'h80be;
17'h1425:	data_out=16'h364;
17'h1426:	data_out=16'h8577;
17'h1427:	data_out=16'h8046;
17'h1428:	data_out=16'h80bd;
17'h1429:	data_out=16'h855d;
17'h142a:	data_out=16'h881a;
17'h142b:	data_out=16'h803e;
17'h142c:	data_out=16'h21b;
17'h142d:	data_out=16'h6f5;
17'h142e:	data_out=16'h85e3;
17'h142f:	data_out=16'h50d;
17'h1430:	data_out=16'ha00;
17'h1431:	data_out=16'h3d;
17'h1432:	data_out=16'ha00;
17'h1433:	data_out=16'h8a00;
17'h1434:	data_out=16'h8279;
17'h1435:	data_out=16'h9f9;
17'h1436:	data_out=16'h83f6;
17'h1437:	data_out=16'h8407;
17'h1438:	data_out=16'h8287;
17'h1439:	data_out=16'h8a00;
17'h143a:	data_out=16'h8575;
17'h143b:	data_out=16'h946;
17'h143c:	data_out=16'h2eb;
17'h143d:	data_out=16'h814b;
17'h143e:	data_out=16'h80ba;
17'h143f:	data_out=16'ha00;
17'h1440:	data_out=16'h829;
17'h1441:	data_out=16'h104;
17'h1442:	data_out=16'ha00;
17'h1443:	data_out=16'h80a2;
17'h1444:	data_out=16'h35c;
17'h1445:	data_out=16'h8089;
17'h1446:	data_out=16'h119;
17'h1447:	data_out=16'h82f3;
17'h1448:	data_out=16'h82ed;
17'h1449:	data_out=16'h384;
17'h144a:	data_out=16'h765;
17'h144b:	data_out=16'ha00;
17'h144c:	data_out=16'h36c;
17'h144d:	data_out=16'h25;
17'h144e:	data_out=16'h834c;
17'h144f:	data_out=16'h25d;
17'h1450:	data_out=16'h3e2;
17'h1451:	data_out=16'h8021;
17'h1452:	data_out=16'h805f;
17'h1453:	data_out=16'h10c;
17'h1454:	data_out=16'heb;
17'h1455:	data_out=16'h82b8;
17'h1456:	data_out=16'h8542;
17'h1457:	data_out=16'h84b4;
17'h1458:	data_out=16'h81a5;
17'h1459:	data_out=16'h540;
17'h145a:	data_out=16'h81e6;
17'h145b:	data_out=16'h9e;
17'h145c:	data_out=16'h5a1;
17'h145d:	data_out=16'h420;
17'h145e:	data_out=16'h5ac;
17'h145f:	data_out=16'h8302;
17'h1460:	data_out=16'h8427;
17'h1461:	data_out=16'h3a7;
17'h1462:	data_out=16'h8753;
17'h1463:	data_out=16'h8a00;
17'h1464:	data_out=16'h863d;
17'h1465:	data_out=16'ha00;
17'h1466:	data_out=16'h4c0;
17'h1467:	data_out=16'h82e5;
17'h1468:	data_out=16'h80d6;
17'h1469:	data_out=16'h823c;
17'h146a:	data_out=16'h811e;
17'h146b:	data_out=16'ha00;
17'h146c:	data_out=16'h218;
17'h146d:	data_out=16'h8a00;
17'h146e:	data_out=16'h8108;
17'h146f:	data_out=16'ha00;
17'h1470:	data_out=16'h80f5;
17'h1471:	data_out=16'h8a00;
17'h1472:	data_out=16'ha00;
17'h1473:	data_out=16'ha00;
17'h1474:	data_out=16'ha00;
17'h1475:	data_out=16'h50d;
17'h1476:	data_out=16'h842b;
17'h1477:	data_out=16'h46d;
17'h1478:	data_out=16'h220;
17'h1479:	data_out=16'h88df;
17'h147a:	data_out=16'h8a00;
17'h147b:	data_out=16'h80b9;
17'h147c:	data_out=16'h8439;
17'h147d:	data_out=16'h8296;
17'h147e:	data_out=16'h8246;
17'h147f:	data_out=16'h42e;
17'h1480:	data_out=16'h69;
17'h1481:	data_out=16'h2f6;
17'h1482:	data_out=16'h163;
17'h1483:	data_out=16'h560;
17'h1484:	data_out=16'ha00;
17'h1485:	data_out=16'h95f;
17'h1486:	data_out=16'hbd;
17'h1487:	data_out=16'h74;
17'h1488:	data_out=16'h35e;
17'h1489:	data_out=16'h81eb;
17'h148a:	data_out=16'h4cf;
17'h148b:	data_out=16'h33f;
17'h148c:	data_out=16'ha00;
17'h148d:	data_out=16'h1c9;
17'h148e:	data_out=16'he9;
17'h148f:	data_out=16'h815a;
17'h1490:	data_out=16'h1a8;
17'h1491:	data_out=16'h958;
17'h1492:	data_out=16'h825d;
17'h1493:	data_out=16'h5fe;
17'h1494:	data_out=16'h824c;
17'h1495:	data_out=16'hfe;
17'h1496:	data_out=16'h42a;
17'h1497:	data_out=16'h803d;
17'h1498:	data_out=16'h823a;
17'h1499:	data_out=16'h30f;
17'h149a:	data_out=16'ha00;
17'h149b:	data_out=16'h35c;
17'h149c:	data_out=16'h451;
17'h149d:	data_out=16'h4a6;
17'h149e:	data_out=16'h821e;
17'h149f:	data_out=16'h818e;
17'h14a0:	data_out=16'h2bb;
17'h14a1:	data_out=16'he8;
17'h14a2:	data_out=16'h15d;
17'h14a3:	data_out=16'h2d;
17'h14a4:	data_out=16'h1d;
17'h14a5:	data_out=16'h253;
17'h14a6:	data_out=16'h7f;
17'h14a7:	data_out=16'h41b;
17'h14a8:	data_out=16'h117;
17'h14a9:	data_out=16'h55;
17'h14aa:	data_out=16'h817f;
17'h14ab:	data_out=16'h101;
17'h14ac:	data_out=16'h453;
17'h14ad:	data_out=16'h63a;
17'h14ae:	data_out=16'ha0;
17'h14af:	data_out=16'h663;
17'h14b0:	data_out=16'ha00;
17'h14b1:	data_out=16'h368;
17'h14b2:	data_out=16'ha00;
17'h14b3:	data_out=16'h835b;
17'h14b4:	data_out=16'hc1;
17'h14b5:	data_out=16'ha00;
17'h14b6:	data_out=16'h19c;
17'h14b7:	data_out=16'h1e2;
17'h14b8:	data_out=16'hd4;
17'h14b9:	data_out=16'h848b;
17'h14ba:	data_out=16'h839f;
17'h14bb:	data_out=16'h783;
17'h14bc:	data_out=16'h72b;
17'h14bd:	data_out=16'h166;
17'h14be:	data_out=16'h11c;
17'h14bf:	data_out=16'h95b;
17'h14c0:	data_out=16'h419;
17'h14c1:	data_out=16'h54e;
17'h14c2:	data_out=16'h8b0;
17'h14c3:	data_out=16'h1b1;
17'h14c4:	data_out=16'h46f;
17'h14c5:	data_out=16'h4e;
17'h14c6:	data_out=16'h47b;
17'h14c7:	data_out=16'h81d1;
17'h14c8:	data_out=16'h80df;
17'h14c9:	data_out=16'h262;
17'h14ca:	data_out=16'h484;
17'h14cb:	data_out=16'h9ed;
17'h14cc:	data_out=16'h243;
17'h14cd:	data_out=16'h157;
17'h14ce:	data_out=16'h23b;
17'h14cf:	data_out=16'h190;
17'h14d0:	data_out=16'h1ec;
17'h14d1:	data_out=16'h305;
17'h14d2:	data_out=16'h17;
17'h14d3:	data_out=16'h628;
17'h14d4:	data_out=16'h497;
17'h14d5:	data_out=16'h2e4;
17'h14d6:	data_out=16'h809b;
17'h14d7:	data_out=16'h81cd;
17'h14d8:	data_out=16'h389;
17'h14d9:	data_out=16'h357;
17'h14da:	data_out=16'h2bf;
17'h14db:	data_out=16'h455;
17'h14dc:	data_out=16'h493;
17'h14dd:	data_out=16'h5a5;
17'h14de:	data_out=16'h7d5;
17'h14df:	data_out=16'h8077;
17'h14e0:	data_out=16'h19c;
17'h14e1:	data_out=16'h65f;
17'h14e2:	data_out=16'hf;
17'h14e3:	data_out=16'h8306;
17'h14e4:	data_out=16'h817d;
17'h14e5:	data_out=16'h8c2;
17'h14e6:	data_out=16'h2be;
17'h14e7:	data_out=16'h80b1;
17'h14e8:	data_out=16'hf7;
17'h14e9:	data_out=16'h3d2;
17'h14ea:	data_out=16'hd1;
17'h14eb:	data_out=16'ha00;
17'h14ec:	data_out=16'h567;
17'h14ed:	data_out=16'h8309;
17'h14ee:	data_out=16'hd2;
17'h14ef:	data_out=16'ha00;
17'h14f0:	data_out=16'hda;
17'h14f1:	data_out=16'h8639;
17'h14f2:	data_out=16'h968;
17'h14f3:	data_out=16'h7e1;
17'h14f4:	data_out=16'ha00;
17'h14f5:	data_out=16'h84f;
17'h14f6:	data_out=16'h802f;
17'h14f7:	data_out=16'h375;
17'h14f8:	data_out=16'h27e;
17'h14f9:	data_out=16'h804b;
17'h14fa:	data_out=16'h8274;
17'h14fb:	data_out=16'h11a;
17'h14fc:	data_out=16'h82a9;
17'h14fd:	data_out=16'h8013;
17'h14fe:	data_out=16'h11;
17'h14ff:	data_out=16'h2b1;
17'h1500:	data_out=16'h364;
17'h1501:	data_out=16'h2cc;
17'h1502:	data_out=16'h4;
17'h1503:	data_out=16'h691;
17'h1504:	data_out=16'h4bc;
17'h1505:	data_out=16'h771;
17'h1506:	data_out=16'h1cd;
17'h1507:	data_out=16'h8300;
17'h1508:	data_out=16'h803d;
17'h1509:	data_out=16'h84fb;
17'h150a:	data_out=16'h34a;
17'h150b:	data_out=16'h320;
17'h150c:	data_out=16'h34f;
17'h150d:	data_out=16'h68e;
17'h150e:	data_out=16'h96;
17'h150f:	data_out=16'h160;
17'h1510:	data_out=16'h81d7;
17'h1511:	data_out=16'h3ae;
17'h1512:	data_out=16'h818f;
17'h1513:	data_out=16'h7d9;
17'h1514:	data_out=16'h442;
17'h1515:	data_out=16'h327;
17'h1516:	data_out=16'h838;
17'h1517:	data_out=16'h662;
17'h1518:	data_out=16'h8122;
17'h1519:	data_out=16'h800d;
17'h151a:	data_out=16'h63f;
17'h151b:	data_out=16'h491;
17'h151c:	data_out=16'h7bc;
17'h151d:	data_out=16'h163;
17'h151e:	data_out=16'h48f;
17'h151f:	data_out=16'h8025;
17'h1520:	data_out=16'h259;
17'h1521:	data_out=16'h8f;
17'h1522:	data_out=16'h83b3;
17'h1523:	data_out=16'h8594;
17'h1524:	data_out=16'h8595;
17'h1525:	data_out=16'h82bb;
17'h1526:	data_out=16'h8178;
17'h1527:	data_out=16'h155;
17'h1528:	data_out=16'hb6;
17'h1529:	data_out=16'h638;
17'h152a:	data_out=16'h8063;
17'h152b:	data_out=16'h833a;
17'h152c:	data_out=16'h747;
17'h152d:	data_out=16'h7e;
17'h152e:	data_out=16'h1;
17'h152f:	data_out=16'h53d;
17'h1530:	data_out=16'h760;
17'h1531:	data_out=16'h36a;
17'h1532:	data_out=16'h765;
17'h1533:	data_out=16'h344;
17'h1534:	data_out=16'h8076;
17'h1535:	data_out=16'h4ce;
17'h1536:	data_out=16'h80c6;
17'h1537:	data_out=16'h95;
17'h1538:	data_out=16'h8057;
17'h1539:	data_out=16'h313;
17'h153a:	data_out=16'h8581;
17'h153b:	data_out=16'h55a;
17'h153c:	data_out=16'h496;
17'h153d:	data_out=16'h288;
17'h153e:	data_out=16'hbb;
17'h153f:	data_out=16'h774;
17'h1540:	data_out=16'h80a8;
17'h1541:	data_out=16'h39e;
17'h1542:	data_out=16'h800c;
17'h1543:	data_out=16'h29c;
17'h1544:	data_out=16'h4d0;
17'h1545:	data_out=16'h351;
17'h1546:	data_out=16'h80fe;
17'h1547:	data_out=16'h845d;
17'h1548:	data_out=16'h82a8;
17'h1549:	data_out=16'h8315;
17'h154a:	data_out=16'h819f;
17'h154b:	data_out=16'h8170;
17'h154c:	data_out=16'h8348;
17'h154d:	data_out=16'h82ec;
17'h154e:	data_out=16'h19a;
17'h154f:	data_out=16'h8387;
17'h1550:	data_out=16'h80fe;
17'h1551:	data_out=16'h78c;
17'h1552:	data_out=16'h8579;
17'h1553:	data_out=16'h2a0;
17'h1554:	data_out=16'h2f7;
17'h1555:	data_out=16'h4d3;
17'h1556:	data_out=16'h8253;
17'h1557:	data_out=16'h8451;
17'h1558:	data_out=16'h2ff;
17'h1559:	data_out=16'h8166;
17'h155a:	data_out=16'h1f6;
17'h155b:	data_out=16'h5d9;
17'h155c:	data_out=16'h33a;
17'h155d:	data_out=16'h3a2;
17'h155e:	data_out=16'h528;
17'h155f:	data_out=16'h803b;
17'h1560:	data_out=16'h8;
17'h1561:	data_out=16'h6f8;
17'h1562:	data_out=16'h5b9;
17'h1563:	data_out=16'h35c;
17'h1564:	data_out=16'h81ca;
17'h1565:	data_out=16'h2a3;
17'h1566:	data_out=16'h8130;
17'h1567:	data_out=16'h836f;
17'h1568:	data_out=16'ha0;
17'h1569:	data_out=16'h80d8;
17'h156a:	data_out=16'h7e;
17'h156b:	data_out=16'h61c;
17'h156c:	data_out=16'h5d9;
17'h156d:	data_out=16'h359;
17'h156e:	data_out=16'h85;
17'h156f:	data_out=16'h6f9;
17'h1570:	data_out=16'h9a;
17'h1571:	data_out=16'h809f;
17'h1572:	data_out=16'h8b6;
17'h1573:	data_out=16'h6f7;
17'h1574:	data_out=16'h76d;
17'h1575:	data_out=16'h9ff;
17'h1576:	data_out=16'h836a;
17'h1577:	data_out=16'h80f6;
17'h1578:	data_out=16'h3b8;
17'h1579:	data_out=16'h4a;
17'h157a:	data_out=16'h3c8;
17'h157b:	data_out=16'hb9;
17'h157c:	data_out=16'h8156;
17'h157d:	data_out=16'h2f3;
17'h157e:	data_out=16'h82d8;
17'h157f:	data_out=16'h8050;
17'h1580:	data_out=16'h898;
17'h1581:	data_out=16'h4ba;
17'h1582:	data_out=16'h84c2;
17'h1583:	data_out=16'h6f1;
17'h1584:	data_out=16'h500;
17'h1585:	data_out=16'h746;
17'h1586:	data_out=16'h35;
17'h1587:	data_out=16'h85c4;
17'h1588:	data_out=16'h8242;
17'h1589:	data_out=16'h8657;
17'h158a:	data_out=16'h6a9;
17'h158b:	data_out=16'h1c5;
17'h158c:	data_out=16'h1d4;
17'h158d:	data_out=16'h525;
17'h158e:	data_out=16'h80e9;
17'h158f:	data_out=16'h840e;
17'h1590:	data_out=16'h8415;
17'h1591:	data_out=16'h615;
17'h1592:	data_out=16'h873b;
17'h1593:	data_out=16'h740;
17'h1594:	data_out=16'h27d;
17'h1595:	data_out=16'h3ca;
17'h1596:	data_out=16'h958;
17'h1597:	data_out=16'h4d3;
17'h1598:	data_out=16'h8341;
17'h1599:	data_out=16'h25d;
17'h159a:	data_out=16'h6c4;
17'h159b:	data_out=16'h228;
17'h159c:	data_out=16'h941;
17'h159d:	data_out=16'h38e;
17'h159e:	data_out=16'h21d;
17'h159f:	data_out=16'h84a2;
17'h15a0:	data_out=16'h40a;
17'h15a1:	data_out=16'h80ed;
17'h15a2:	data_out=16'h868c;
17'h15a3:	data_out=16'h8601;
17'h15a4:	data_out=16'h85ff;
17'h15a5:	data_out=16'h85fc;
17'h15a6:	data_out=16'h82bc;
17'h15a7:	data_out=16'h34a;
17'h15a8:	data_out=16'h80cf;
17'h15a9:	data_out=16'h453;
17'h15aa:	data_out=16'h86b6;
17'h15ab:	data_out=16'h8211;
17'h15ac:	data_out=16'h884;
17'h15ad:	data_out=16'h821e;
17'h15ae:	data_out=16'h874d;
17'h15af:	data_out=16'h537;
17'h15b0:	data_out=16'h842;
17'h15b1:	data_out=16'h9cc;
17'h15b2:	data_out=16'h88d;
17'h15b3:	data_out=16'h176;
17'h15b4:	data_out=16'h326;
17'h15b5:	data_out=16'h33b;
17'h15b6:	data_out=16'h848a;
17'h15b7:	data_out=16'h84c2;
17'h15b8:	data_out=16'h1eb;
17'h15b9:	data_out=16'h13b;
17'h15ba:	data_out=16'h87fa;
17'h15bb:	data_out=16'h761;
17'h15bc:	data_out=16'h2b5;
17'h15bd:	data_out=16'h5cb;
17'h15be:	data_out=16'h80da;
17'h15bf:	data_out=16'h837;
17'h15c0:	data_out=16'h81e4;
17'h15c1:	data_out=16'h126;
17'h15c2:	data_out=16'h8314;
17'h15c3:	data_out=16'h55;
17'h15c4:	data_out=16'h69e;
17'h15c5:	data_out=16'h3f5;
17'h15c6:	data_out=16'h82d7;
17'h15c7:	data_out=16'h8748;
17'h15c8:	data_out=16'h88b8;
17'h15c9:	data_out=16'h85f0;
17'h15ca:	data_out=16'h8552;
17'h15cb:	data_out=16'h84c8;
17'h15cc:	data_out=16'h87eb;
17'h15cd:	data_out=16'h85a3;
17'h15ce:	data_out=16'h849c;
17'h15cf:	data_out=16'h8805;
17'h15d0:	data_out=16'h82c6;
17'h15d1:	data_out=16'h5d2;
17'h15d2:	data_out=16'h85d9;
17'h15d3:	data_out=16'h16a;
17'h15d4:	data_out=16'h331;
17'h15d5:	data_out=16'h2d4;
17'h15d6:	data_out=16'h8656;
17'h15d7:	data_out=16'h8844;
17'h15d8:	data_out=16'h4c;
17'h15d9:	data_out=16'h82bf;
17'h15da:	data_out=16'h800c;
17'h15db:	data_out=16'h7d8;
17'h15dc:	data_out=16'h54c;
17'h15dd:	data_out=16'h169;
17'h15de:	data_out=16'h4f3;
17'h15df:	data_out=16'h8218;
17'h15e0:	data_out=16'h81a1;
17'h15e1:	data_out=16'h993;
17'h15e2:	data_out=16'h480;
17'h15e3:	data_out=16'h189;
17'h15e4:	data_out=16'h68;
17'h15e5:	data_out=16'h2a4;
17'h15e6:	data_out=16'h57;
17'h15e7:	data_out=16'h88f8;
17'h15e8:	data_out=16'h80e2;
17'h15e9:	data_out=16'h847d;
17'h15ea:	data_out=16'h8102;
17'h15eb:	data_out=16'h779;
17'h15ec:	data_out=16'ha00;
17'h15ed:	data_out=16'h18b;
17'h15ee:	data_out=16'h80fc;
17'h15ef:	data_out=16'h6fc;
17'h15f0:	data_out=16'h80e6;
17'h15f1:	data_out=16'h86fb;
17'h15f2:	data_out=16'h8b8;
17'h15f3:	data_out=16'h7d5;
17'h15f4:	data_out=16'h846;
17'h15f5:	data_out=16'h9b9;
17'h15f6:	data_out=16'h8317;
17'h15f7:	data_out=16'h8613;
17'h15f8:	data_out=16'h339;
17'h15f9:	data_out=16'h876f;
17'h15fa:	data_out=16'h1e3;
17'h15fb:	data_out=16'h80d6;
17'h15fc:	data_out=16'h82d1;
17'h15fd:	data_out=16'h802c;
17'h15fe:	data_out=16'h846f;
17'h15ff:	data_out=16'h8367;
17'h1600:	data_out=16'h942;
17'h1601:	data_out=16'h70c;
17'h1602:	data_out=16'h846e;
17'h1603:	data_out=16'h2d7;
17'h1604:	data_out=16'h5ee;
17'h1605:	data_out=16'h49f;
17'h1606:	data_out=16'h8284;
17'h1607:	data_out=16'h802f;
17'h1608:	data_out=16'h2ac;
17'h1609:	data_out=16'h8025;
17'h160a:	data_out=16'h9c9;
17'h160b:	data_out=16'h32a;
17'h160c:	data_out=16'h71a;
17'h160d:	data_out=16'h8093;
17'h160e:	data_out=16'h8115;
17'h160f:	data_out=16'h8593;
17'h1610:	data_out=16'h1a7;
17'h1611:	data_out=16'ha00;
17'h1612:	data_out=16'h84c5;
17'h1613:	data_out=16'h309;
17'h1614:	data_out=16'h842b;
17'h1615:	data_out=16'h294;
17'h1616:	data_out=16'h3f1;
17'h1617:	data_out=16'h8349;
17'h1618:	data_out=16'h82f8;
17'h1619:	data_out=16'h909;
17'h161a:	data_out=16'h66e;
17'h161b:	data_out=16'hde;
17'h161c:	data_out=16'h541;
17'h161d:	data_out=16'h8c4;
17'h161e:	data_out=16'h822b;
17'h161f:	data_out=16'h8532;
17'h1620:	data_out=16'h544;
17'h1621:	data_out=16'h810d;
17'h1622:	data_out=16'h8064;
17'h1623:	data_out=16'h262;
17'h1624:	data_out=16'h267;
17'h1625:	data_out=16'ha;
17'h1626:	data_out=16'h42e;
17'h1627:	data_out=16'h84f;
17'h1628:	data_out=16'h8102;
17'h1629:	data_out=16'h81f9;
17'h162a:	data_out=16'h8493;
17'h162b:	data_out=16'ha00;
17'h162c:	data_out=16'h3ca;
17'h162d:	data_out=16'h462;
17'h162e:	data_out=16'h8599;
17'h162f:	data_out=16'h363;
17'h1630:	data_out=16'h876;
17'h1631:	data_out=16'ha00;
17'h1632:	data_out=16'h8c2;
17'h1633:	data_out=16'h843b;
17'h1634:	data_out=16'h8f6;
17'h1635:	data_out=16'h7fc;
17'h1636:	data_out=16'h80fa;
17'h1637:	data_out=16'h846c;
17'h1638:	data_out=16'h704;
17'h1639:	data_out=16'h834e;
17'h163a:	data_out=16'h8374;
17'h163b:	data_out=16'h980;
17'h163c:	data_out=16'h11d;
17'h163d:	data_out=16'h651;
17'h163e:	data_out=16'h8104;
17'h163f:	data_out=16'h587;
17'h1640:	data_out=16'h8010;
17'h1641:	data_out=16'h814a;
17'h1642:	data_out=16'h1a1;
17'h1643:	data_out=16'h8392;
17'h1644:	data_out=16'h7fb;
17'h1645:	data_out=16'h2a8;
17'h1646:	data_out=16'h78;
17'h1647:	data_out=16'h8272;
17'h1648:	data_out=16'h85de;
17'h1649:	data_out=16'h13;
17'h164a:	data_out=16'h80c6;
17'h164b:	data_out=16'h2b6;
17'h164c:	data_out=16'h83cf;
17'h164d:	data_out=16'h8075;
17'h164e:	data_out=16'h8273;
17'h164f:	data_out=16'h832b;
17'h1650:	data_out=16'h825f;
17'h1651:	data_out=16'h48;
17'h1652:	data_out=16'h2fe;
17'h1653:	data_out=16'h51f;
17'h1654:	data_out=16'h3f6;
17'h1655:	data_out=16'h825f;
17'h1656:	data_out=16'h83f9;
17'h1657:	data_out=16'h83b9;
17'h1658:	data_out=16'h8268;
17'h1659:	data_out=16'h80aa;
17'h165a:	data_out=16'hc5;
17'h165b:	data_out=16'h5c4;
17'h165c:	data_out=16'h5f7;
17'h165d:	data_out=16'h178;
17'h165e:	data_out=16'h360;
17'h165f:	data_out=16'h81a1;
17'h1660:	data_out=16'h627;
17'h1661:	data_out=16'h7eb;
17'h1662:	data_out=16'h82cb;
17'h1663:	data_out=16'h8421;
17'h1664:	data_out=16'h850;
17'h1665:	data_out=16'h6c8;
17'h1666:	data_out=16'h7ad;
17'h1667:	data_out=16'h8480;
17'h1668:	data_out=16'h8115;
17'h1669:	data_out=16'h86;
17'h166a:	data_out=16'h8133;
17'h166b:	data_out=16'h686;
17'h166c:	data_out=16'h859;
17'h166d:	data_out=16'h83fc;
17'h166e:	data_out=16'h812a;
17'h166f:	data_out=16'h436;
17'h1670:	data_out=16'h8114;
17'h1671:	data_out=16'h881f;
17'h1672:	data_out=16'h543;
17'h1673:	data_out=16'h534;
17'h1674:	data_out=16'h86c;
17'h1675:	data_out=16'h3df;
17'h1676:	data_out=16'h7ea;
17'h1677:	data_out=16'h8305;
17'h1678:	data_out=16'h80f1;
17'h1679:	data_out=16'h866b;
17'h167a:	data_out=16'h8427;
17'h167b:	data_out=16'h80fe;
17'h167c:	data_out=16'h825d;
17'h167d:	data_out=16'h841b;
17'h167e:	data_out=16'hd7;
17'h167f:	data_out=16'h81fd;
17'h1680:	data_out=16'h691;
17'h1681:	data_out=16'h6c3;
17'h1682:	data_out=16'hd4;
17'h1683:	data_out=16'h48f;
17'h1684:	data_out=16'h6ff;
17'h1685:	data_out=16'h671;
17'h1686:	data_out=16'h818f;
17'h1687:	data_out=16'h7b;
17'h1688:	data_out=16'h795;
17'h1689:	data_out=16'h8071;
17'h168a:	data_out=16'h93b;
17'h168b:	data_out=16'h646;
17'h168c:	data_out=16'h995;
17'h168d:	data_out=16'h20e;
17'h168e:	data_out=16'h33;
17'h168f:	data_out=16'h80a2;
17'h1690:	data_out=16'h270;
17'h1691:	data_out=16'h8ca;
17'h1692:	data_out=16'h821b;
17'h1693:	data_out=16'h561;
17'h1694:	data_out=16'h80f3;
17'h1695:	data_out=16'h1b1;
17'h1696:	data_out=16'h50a;
17'h1697:	data_out=16'h98;
17'h1698:	data_out=16'h8170;
17'h1699:	data_out=16'h484;
17'h169a:	data_out=16'h75d;
17'h169b:	data_out=16'h4e0;
17'h169c:	data_out=16'h615;
17'h169d:	data_out=16'h7e9;
17'h169e:	data_out=16'h4b;
17'h169f:	data_out=16'h8337;
17'h16a0:	data_out=16'h34b;
17'h16a1:	data_out=16'h49;
17'h16a2:	data_out=16'h8052;
17'h16a3:	data_out=16'h17a;
17'h16a4:	data_out=16'h17c;
17'h16a5:	data_out=16'h16b;
17'h16a6:	data_out=16'h641;
17'h16a7:	data_out=16'h76a;
17'h16a8:	data_out=16'h65;
17'h16a9:	data_out=16'h245;
17'h16aa:	data_out=16'h10d;
17'h16ab:	data_out=16'h6e4;
17'h16ac:	data_out=16'h4c4;
17'h16ad:	data_out=16'h6e5;
17'h16ae:	data_out=16'h48;
17'h16af:	data_out=16'h512;
17'h16b0:	data_out=16'h9fe;
17'h16b1:	data_out=16'h9c0;
17'h16b2:	data_out=16'ha00;
17'h16b3:	data_out=16'h817b;
17'h16b4:	data_out=16'h6b4;
17'h16b5:	data_out=16'ha00;
17'h16b6:	data_out=16'h2c3;
17'h16b7:	data_out=16'hd3;
17'h16b8:	data_out=16'h3df;
17'h16b9:	data_out=16'h8133;
17'h16ba:	data_out=16'h833c;
17'h16bb:	data_out=16'h8fa;
17'h16bc:	data_out=16'h6f1;
17'h16bd:	data_out=16'h3f1;
17'h16be:	data_out=16'h5c;
17'h16bf:	data_out=16'h713;
17'h16c0:	data_out=16'h13b;
17'h16c1:	data_out=16'h370;
17'h16c2:	data_out=16'h3dd;
17'h16c3:	data_out=16'h8176;
17'h16c4:	data_out=16'h723;
17'h16c5:	data_out=16'h117;
17'h16c6:	data_out=16'h505;
17'h16c7:	data_out=16'h8183;
17'h16c8:	data_out=16'h830a;
17'h16c9:	data_out=16'h179;
17'h16ca:	data_out=16'h38a;
17'h16cb:	data_out=16'h67a;
17'h16cc:	data_out=16'he8;
17'h16cd:	data_out=16'h8028;
17'h16ce:	data_out=16'h376;
17'h16cf:	data_out=16'hb9;
17'h16d0:	data_out=16'h8066;
17'h16d1:	data_out=16'h381;
17'h16d2:	data_out=16'h1b3;
17'h16d3:	data_out=16'h7ab;
17'h16d4:	data_out=16'h46c;
17'h16d5:	data_out=16'h30c;
17'h16d6:	data_out=16'h8185;
17'h16d7:	data_out=16'h81e0;
17'h16d8:	data_out=16'h33a;
17'h16d9:	data_out=16'h8a;
17'h16da:	data_out=16'h52d;
17'h16db:	data_out=16'h629;
17'h16dc:	data_out=16'h692;
17'h16dd:	data_out=16'h441;
17'h16de:	data_out=16'h5ac;
17'h16df:	data_out=16'h8113;
17'h16e0:	data_out=16'h75d;
17'h16e1:	data_out=16'h84b;
17'h16e2:	data_out=16'h87;
17'h16e3:	data_out=16'h80d2;
17'h16e4:	data_out=16'h462;
17'h16e5:	data_out=16'h575;
17'h16e6:	data_out=16'h40e;
17'h16e7:	data_out=16'h81a9;
17'h16e8:	data_out=16'h4b;
17'h16e9:	data_out=16'h575;
17'h16ea:	data_out=16'h2a;
17'h16eb:	data_out=16'h6aa;
17'h16ec:	data_out=16'h83f;
17'h16ed:	data_out=16'h8124;
17'h16ee:	data_out=16'h22;
17'h16ef:	data_out=16'h71b;
17'h16f0:	data_out=16'h37;
17'h16f1:	data_out=16'h8470;
17'h16f2:	data_out=16'h706;
17'h16f3:	data_out=16'h593;
17'h16f4:	data_out=16'h9fd;
17'h16f5:	data_out=16'h950;
17'h16f6:	data_out=16'h460;
17'h16f7:	data_out=16'h139;
17'h16f8:	data_out=16'hce;
17'h16f9:	data_out=16'h6a;
17'h16fa:	data_out=16'h811c;
17'h16fb:	data_out=16'h67;
17'h16fc:	data_out=16'h81f6;
17'h16fd:	data_out=16'h82a7;
17'h16fe:	data_out=16'h157;
17'h16ff:	data_out=16'hf2;
17'h1700:	data_out=16'h54;
17'h1701:	data_out=16'h2e0;
17'h1702:	data_out=16'h19d;
17'h1703:	data_out=16'h41c;
17'h1704:	data_out=16'h616;
17'h1705:	data_out=16'h637;
17'h1706:	data_out=16'h60;
17'h1707:	data_out=16'h10a;
17'h1708:	data_out=16'h2fb;
17'h1709:	data_out=16'h81a4;
17'h170a:	data_out=16'h42b;
17'h170b:	data_out=16'h3ef;
17'h170c:	data_out=16'h7f3;
17'h170d:	data_out=16'h29b;
17'h170e:	data_out=16'h9c;
17'h170f:	data_out=16'h14;
17'h1710:	data_out=16'h121;
17'h1711:	data_out=16'h50e;
17'h1712:	data_out=16'h8085;
17'h1713:	data_out=16'h47e;
17'h1714:	data_out=16'h5a;
17'h1715:	data_out=16'h98;
17'h1716:	data_out=16'h317;
17'h1717:	data_out=16'h1da;
17'h1718:	data_out=16'h80a9;
17'h1719:	data_out=16'h224;
17'h171a:	data_out=16'h73a;
17'h171b:	data_out=16'h3c7;
17'h171c:	data_out=16'h385;
17'h171d:	data_out=16'h3a9;
17'h171e:	data_out=16'hd;
17'h171f:	data_out=16'h811f;
17'h1720:	data_out=16'h1de;
17'h1721:	data_out=16'hb1;
17'h1722:	data_out=16'ha1;
17'h1723:	data_out=16'h8089;
17'h1724:	data_out=16'h8083;
17'h1725:	data_out=16'h1af;
17'h1726:	data_out=16'hfd;
17'h1727:	data_out=16'h33b;
17'h1728:	data_out=16'hc3;
17'h1729:	data_out=16'h1fc;
17'h172a:	data_out=16'hb1;
17'h172b:	data_out=16'h8086;
17'h172c:	data_out=16'h399;
17'h172d:	data_out=16'h3b7;
17'h172e:	data_out=16'h169;
17'h172f:	data_out=16'h456;
17'h1730:	data_out=16'h9cf;
17'h1731:	data_out=16'h31b;
17'h1732:	data_out=16'h9bf;
17'h1733:	data_out=16'h8084;
17'h1734:	data_out=16'h21b;
17'h1735:	data_out=16'h81c;
17'h1736:	data_out=16'h1e5;
17'h1737:	data_out=16'h219;
17'h1738:	data_out=16'h7e;
17'h1739:	data_out=16'h81c9;
17'h173a:	data_out=16'h81df;
17'h173b:	data_out=16'h560;
17'h173c:	data_out=16'h5eb;
17'h173d:	data_out=16'h53;
17'h173e:	data_out=16'hcd;
17'h173f:	data_out=16'h634;
17'h1740:	data_out=16'h23f;
17'h1741:	data_out=16'h41f;
17'h1742:	data_out=16'h357;
17'h1743:	data_out=16'h194;
17'h1744:	data_out=16'h358;
17'h1745:	data_out=16'h8009;
17'h1746:	data_out=16'h445;
17'h1747:	data_out=16'h81b0;
17'h1748:	data_out=16'h8085;
17'h1749:	data_out=16'h1ba;
17'h174a:	data_out=16'h3b5;
17'h174b:	data_out=16'h60a;
17'h174c:	data_out=16'h1e6;
17'h174d:	data_out=16'hb1;
17'h174e:	data_out=16'h375;
17'h174f:	data_out=16'h174;
17'h1750:	data_out=16'h10a;
17'h1751:	data_out=16'h2cb;
17'h1752:	data_out=16'h8059;
17'h1753:	data_out=16'h50f;
17'h1754:	data_out=16'h361;
17'h1755:	data_out=16'h30a;
17'h1756:	data_out=16'h74;
17'h1757:	data_out=16'h80c9;
17'h1758:	data_out=16'h348;
17'h1759:	data_out=16'h22a;
17'h175a:	data_out=16'h331;
17'h175b:	data_out=16'h38c;
17'h175c:	data_out=16'h3b0;
17'h175d:	data_out=16'h438;
17'h175e:	data_out=16'h590;
17'h175f:	data_out=16'h8027;
17'h1760:	data_out=16'h271;
17'h1761:	data_out=16'h504;
17'h1762:	data_out=16'h197;
17'h1763:	data_out=16'h803a;
17'h1764:	data_out=16'h48;
17'h1765:	data_out=16'h462;
17'h1766:	data_out=16'h1c6;
17'h1767:	data_out=16'h8042;
17'h1768:	data_out=16'hba;
17'h1769:	data_out=16'h3bf;
17'h176a:	data_out=16'h90;
17'h176b:	data_out=16'h547;
17'h176c:	data_out=16'h43d;
17'h176d:	data_out=16'h804e;
17'h176e:	data_out=16'h91;
17'h176f:	data_out=16'h82d;
17'h1770:	data_out=16'h9b;
17'h1771:	data_out=16'h823c;
17'h1772:	data_out=16'h605;
17'h1773:	data_out=16'h4b8;
17'h1774:	data_out=16'h9ea;
17'h1775:	data_out=16'h757;
17'h1776:	data_out=16'h8150;
17'h1777:	data_out=16'h277;
17'h1778:	data_out=16'h251;
17'h1779:	data_out=16'h1e0;
17'h177a:	data_out=16'h3d;
17'h177b:	data_out=16'hcc;
17'h177c:	data_out=16'h8126;
17'h177d:	data_out=16'h8014;
17'h177e:	data_out=16'h80b7;
17'h177f:	data_out=16'h21c;
17'h1780:	data_out=16'h43;
17'h1781:	data_out=16'h24f;
17'h1782:	data_out=16'hea;
17'h1783:	data_out=16'h35e;
17'h1784:	data_out=16'h5d6;
17'h1785:	data_out=16'h51a;
17'h1786:	data_out=16'ha1;
17'h1787:	data_out=16'h190;
17'h1788:	data_out=16'h13c;
17'h1789:	data_out=16'h8166;
17'h178a:	data_out=16'h300;
17'h178b:	data_out=16'h223;
17'h178c:	data_out=16'h664;
17'h178d:	data_out=16'h1b8;
17'h178e:	data_out=16'h70;
17'h178f:	data_out=16'h8059;
17'h1790:	data_out=16'he8;
17'h1791:	data_out=16'h46a;
17'h1792:	data_out=16'h80f1;
17'h1793:	data_out=16'h346;
17'h1794:	data_out=16'h8042;
17'h1795:	data_out=16'he1;
17'h1796:	data_out=16'h23e;
17'h1797:	data_out=16'hc6;
17'h1798:	data_out=16'h808a;
17'h1799:	data_out=16'h2d7;
17'h179a:	data_out=16'h697;
17'h179b:	data_out=16'h2a7;
17'h179c:	data_out=16'h2f0;
17'h179d:	data_out=16'h321;
17'h179e:	data_out=16'h806f;
17'h179f:	data_out=16'h8078;
17'h17a0:	data_out=16'h210;
17'h17a1:	data_out=16'h7f;
17'h17a2:	data_out=16'h12d;
17'h17a3:	data_out=16'h6;
17'h17a4:	data_out=16'h2;
17'h17a5:	data_out=16'h1a2;
17'h17a6:	data_out=16'h80b5;
17'h17a7:	data_out=16'h2d1;
17'h17a8:	data_out=16'h8e;
17'h17a9:	data_out=16'hb8;
17'h17aa:	data_out=16'h809b;
17'h17ab:	data_out=16'h8026;
17'h17ac:	data_out=16'h2b1;
17'h17ad:	data_out=16'h33d;
17'h17ae:	data_out=16'ha;
17'h17af:	data_out=16'h40c;
17'h17b0:	data_out=16'h815;
17'h17b1:	data_out=16'h291;
17'h17b2:	data_out=16'h80c;
17'h17b3:	data_out=16'h80d4;
17'h17b4:	data_out=16'h1ef;
17'h17b5:	data_out=16'h684;
17'h17b6:	data_out=16'h114;
17'h17b7:	data_out=16'h13a;
17'h17b8:	data_out=16'h90;
17'h17b9:	data_out=16'h81b6;
17'h17ba:	data_out=16'h8101;
17'h17bb:	data_out=16'h3f1;
17'h17bc:	data_out=16'h422;
17'h17bd:	data_out=16'h4f;
17'h17be:	data_out=16'h92;
17'h17bf:	data_out=16'h518;
17'h17c0:	data_out=16'h242;
17'h17c1:	data_out=16'h306;
17'h17c2:	data_out=16'h2f2;
17'h17c3:	data_out=16'h15d;
17'h17c4:	data_out=16'h289;
17'h17c5:	data_out=16'h34;
17'h17c6:	data_out=16'h39c;
17'h17c7:	data_out=16'h80fb;
17'h17c8:	data_out=16'h808e;
17'h17c9:	data_out=16'h1af;
17'h17ca:	data_out=16'h2e5;
17'h17cb:	data_out=16'h587;
17'h17cc:	data_out=16'h1b6;
17'h17cd:	data_out=16'h16d;
17'h17ce:	data_out=16'h194;
17'h17cf:	data_out=16'h15c;
17'h17d0:	data_out=16'h137;
17'h17d1:	data_out=16'h1c9;
17'h17d2:	data_out=16'h35;
17'h17d3:	data_out=16'h3f6;
17'h17d4:	data_out=16'h2fa;
17'h17d5:	data_out=16'h1c5;
17'h17d6:	data_out=16'h59;
17'h17d7:	data_out=16'h801d;
17'h17d8:	data_out=16'h213;
17'h17d9:	data_out=16'h284;
17'h17da:	data_out=16'h216;
17'h17db:	data_out=16'h2de;
17'h17dc:	data_out=16'h300;
17'h17dd:	data_out=16'h35c;
17'h17de:	data_out=16'h4bc;
17'h17df:	data_out=16'h2e;
17'h17e0:	data_out=16'he4;
17'h17e1:	data_out=16'h3d9;
17'h17e2:	data_out=16'h129;
17'h17e3:	data_out=16'h80a2;
17'h17e4:	data_out=16'hab;
17'h17e5:	data_out=16'h434;
17'h17e6:	data_out=16'h234;
17'h17e7:	data_out=16'h80c2;
17'h17e8:	data_out=16'h7d;
17'h17e9:	data_out=16'h1ee;
17'h17ea:	data_out=16'h6a;
17'h17eb:	data_out=16'h4cd;
17'h17ec:	data_out=16'h340;
17'h17ed:	data_out=16'h80a5;
17'h17ee:	data_out=16'h6d;
17'h17ef:	data_out=16'h72f;
17'h17f0:	data_out=16'h77;
17'h17f1:	data_out=16'h82d5;
17'h17f2:	data_out=16'h4e4;
17'h17f3:	data_out=16'h4a3;
17'h17f4:	data_out=16'h829;
17'h17f5:	data_out=16'h4d7;
17'h17f6:	data_out=16'h816a;
17'h17f7:	data_out=16'h20f;
17'h17f8:	data_out=16'h266;
17'h17f9:	data_out=16'h34;
17'h17fa:	data_out=16'h8050;
17'h17fb:	data_out=16'h91;
17'h17fc:	data_out=16'h8076;
17'h17fd:	data_out=16'h47;
17'h17fe:	data_out=16'h80ce;
17'h17ff:	data_out=16'h1e9;
17'h1800:	data_out=16'h1e2;
17'h1801:	data_out=16'h380;
17'h1802:	data_out=16'h21e;
17'h1803:	data_out=16'h356;
17'h1804:	data_out=16'h496;
17'h1805:	data_out=16'h4e3;
17'h1806:	data_out=16'h88;
17'h1807:	data_out=16'hc2;
17'h1808:	data_out=16'h280;
17'h1809:	data_out=16'h812d;
17'h180a:	data_out=16'h3ee;
17'h180b:	data_out=16'h308;
17'h180c:	data_out=16'h492;
17'h180d:	data_out=16'h203;
17'h180e:	data_out=16'h84;
17'h180f:	data_out=16'h100;
17'h1810:	data_out=16'h13a;
17'h1811:	data_out=16'h46d;
17'h1812:	data_out=16'h8023;
17'h1813:	data_out=16'h37a;
17'h1814:	data_out=16'h12f;
17'h1815:	data_out=16'h125;
17'h1816:	data_out=16'h29a;
17'h1817:	data_out=16'h21a;
17'h1818:	data_out=16'h8023;
17'h1819:	data_out=16'h1ca;
17'h181a:	data_out=16'h50c;
17'h181b:	data_out=16'h392;
17'h181c:	data_out=16'h40c;
17'h181d:	data_out=16'h40b;
17'h181e:	data_out=16'h109;
17'h181f:	data_out=16'h1;
17'h1820:	data_out=16'h2f8;
17'h1821:	data_out=16'h92;
17'h1822:	data_out=16'h138;
17'h1823:	data_out=16'h18;
17'h1824:	data_out=16'h19;
17'h1825:	data_out=16'h178;
17'h1826:	data_out=16'hc9;
17'h1827:	data_out=16'h3df;
17'h1828:	data_out=16'h9c;
17'h1829:	data_out=16'h1f0;
17'h182a:	data_out=16'hd2;
17'h182b:	data_out=16'h16e;
17'h182c:	data_out=16'h2e4;
17'h182d:	data_out=16'h415;
17'h182e:	data_out=16'h123;
17'h182f:	data_out=16'h442;
17'h1830:	data_out=16'h64b;
17'h1831:	data_out=16'h383;
17'h1832:	data_out=16'h652;
17'h1833:	data_out=16'hae;
17'h1834:	data_out=16'h2c6;
17'h1835:	data_out=16'h5a6;
17'h1836:	data_out=16'h256;
17'h1837:	data_out=16'h25b;
17'h1838:	data_out=16'h209;
17'h1839:	data_out=16'h3;
17'h183a:	data_out=16'h80e3;
17'h183b:	data_out=16'h3dc;
17'h183c:	data_out=16'h502;
17'h183d:	data_out=16'h190;
17'h183e:	data_out=16'ha1;
17'h183f:	data_out=16'h4e1;
17'h1840:	data_out=16'h1a3;
17'h1841:	data_out=16'h3a0;
17'h1842:	data_out=16'h2b3;
17'h1843:	data_out=16'h155;
17'h1844:	data_out=16'h371;
17'h1845:	data_out=16'haf;
17'h1846:	data_out=16'h481;
17'h1847:	data_out=16'h80ce;
17'h1848:	data_out=16'h806d;
17'h1849:	data_out=16'h181;
17'h184a:	data_out=16'h254;
17'h184b:	data_out=16'h449;
17'h184c:	data_out=16'h168;
17'h184d:	data_out=16'h176;
17'h184e:	data_out=16'h276;
17'h184f:	data_out=16'h12b;
17'h1850:	data_out=16'hde;
17'h1851:	data_out=16'h2a3;
17'h1852:	data_out=16'h3a;
17'h1853:	data_out=16'h4d4;
17'h1854:	data_out=16'h3e1;
17'h1855:	data_out=16'h2dc;
17'h1856:	data_out=16'h116;
17'h1857:	data_out=16'h4a;
17'h1858:	data_out=16'h326;
17'h1859:	data_out=16'h22b;
17'h185a:	data_out=16'h30d;
17'h185b:	data_out=16'h3d2;
17'h185c:	data_out=16'h3c9;
17'h185d:	data_out=16'h395;
17'h185e:	data_out=16'h4b5;
17'h185f:	data_out=16'h75;
17'h1860:	data_out=16'h22b;
17'h1861:	data_out=16'h480;
17'h1862:	data_out=16'h232;
17'h1863:	data_out=16'hd8;
17'h1864:	data_out=16'h17a;
17'h1865:	data_out=16'h313;
17'h1866:	data_out=16'h18b;
17'h1867:	data_out=16'h8014;
17'h1868:	data_out=16'h93;
17'h1869:	data_out=16'h2f9;
17'h186a:	data_out=16'h86;
17'h186b:	data_out=16'h460;
17'h186c:	data_out=16'h429;
17'h186d:	data_out=16'hd6;
17'h186e:	data_out=16'h76;
17'h186f:	data_out=16'h566;
17'h1870:	data_out=16'h7a;
17'h1871:	data_out=16'h8181;
17'h1872:	data_out=16'h4ce;
17'h1873:	data_out=16'h4a0;
17'h1874:	data_out=16'h656;
17'h1875:	data_out=16'h593;
17'h1876:	data_out=16'h20;
17'h1877:	data_out=16'h220;
17'h1878:	data_out=16'h20d;
17'h1879:	data_out=16'h15f;
17'h187a:	data_out=16'h11f;
17'h187b:	data_out=16'h98;
17'h187c:	data_out=16'h8016;
17'h187d:	data_out=16'h6c;
17'h187e:	data_out=16'h8033;
17'h187f:	data_out=16'h198;
17'h1880:	data_out=16'h93;
17'h1881:	data_out=16'h144;
17'h1882:	data_out=16'h5e;
17'h1883:	data_out=16'h155;
17'h1884:	data_out=16'h30d;
17'h1885:	data_out=16'h2d3;
17'h1886:	data_out=16'h806b;
17'h1887:	data_out=16'h807c;
17'h1888:	data_out=16'he0;
17'h1889:	data_out=16'h814b;
17'h188a:	data_out=16'h19f;
17'h188b:	data_out=16'h1ed;
17'h188c:	data_out=16'h30b;
17'h188d:	data_out=16'he4;
17'h188e:	data_out=16'hf;
17'h188f:	data_out=16'h8031;
17'h1890:	data_out=16'ha3;
17'h1891:	data_out=16'h28a;
17'h1892:	data_out=16'h80b6;
17'h1893:	data_out=16'h1a7;
17'h1894:	data_out=16'h1;
17'h1895:	data_out=16'h6;
17'h1896:	data_out=16'he3;
17'h1897:	data_out=16'h84;
17'h1898:	data_out=16'h8065;
17'h1899:	data_out=16'h161;
17'h189a:	data_out=16'h360;
17'h189b:	data_out=16'h19f;
17'h189c:	data_out=16'h190;
17'h189d:	data_out=16'h166;
17'h189e:	data_out=16'h8020;
17'h189f:	data_out=16'h80e5;
17'h18a0:	data_out=16'h10f;
17'h18a1:	data_out=16'h10;
17'h18a2:	data_out=16'h8024;
17'h18a3:	data_out=16'h80c3;
17'h18a4:	data_out=16'h80c0;
17'h18a5:	data_out=16'h11e;
17'h18a6:	data_out=16'h802a;
17'h18a7:	data_out=16'h15c;
17'h18a8:	data_out=16'h16;
17'h18a9:	data_out=16'h122;
17'h18aa:	data_out=16'h800b;
17'h18ab:	data_out=16'h70;
17'h18ac:	data_out=16'h162;
17'h18ad:	data_out=16'h2a5;
17'h18ae:	data_out=16'h25;
17'h18af:	data_out=16'h1a5;
17'h18b0:	data_out=16'h40c;
17'h18b1:	data_out=16'h1f7;
17'h18b2:	data_out=16'h40d;
17'h18b3:	data_out=16'h805a;
17'h18b4:	data_out=16'h17b;
17'h18b5:	data_out=16'h3b7;
17'h18b6:	data_out=16'ha9;
17'h18b7:	data_out=16'h82;
17'h18b8:	data_out=16'h90;
17'h18b9:	data_out=16'h80a8;
17'h18ba:	data_out=16'h815a;
17'h18bb:	data_out=16'h23f;
17'h18bc:	data_out=16'h214;
17'h18bd:	data_out=16'h7f;
17'h18be:	data_out=16'h1b;
17'h18bf:	data_out=16'h34e;
17'h18c0:	data_out=16'h78;
17'h18c1:	data_out=16'h13f;
17'h18c2:	data_out=16'h257;
17'h18c3:	data_out=16'h87;
17'h18c4:	data_out=16'h283;
17'h18c5:	data_out=16'h8027;
17'h18c6:	data_out=16'h1bb;
17'h18c7:	data_out=16'h815d;
17'h18c8:	data_out=16'h80ac;
17'h18c9:	data_out=16'hed;
17'h18ca:	data_out=16'h198;
17'h18cb:	data_out=16'h325;
17'h18cc:	data_out=16'hde;
17'h18cd:	data_out=16'h801a;
17'h18ce:	data_out=16'h1d3;
17'h18cf:	data_out=16'h107;
17'h18d0:	data_out=16'h8005;
17'h18d1:	data_out=16'hd0;
17'h18d2:	data_out=16'h80ae;
17'h18d3:	data_out=16'h1e9;
17'h18d4:	data_out=16'h1a3;
17'h18d5:	data_out=16'hd1;
17'h18d6:	data_out=16'h8031;
17'h18d7:	data_out=16'h80ac;
17'h18d8:	data_out=16'h110;
17'h18d9:	data_out=16'h98;
17'h18da:	data_out=16'h132;
17'h18db:	data_out=16'h182;
17'h18dc:	data_out=16'h210;
17'h18dd:	data_out=16'h181;
17'h18de:	data_out=16'h27f;
17'h18df:	data_out=16'h8062;
17'h18e0:	data_out=16'h15f;
17'h18e1:	data_out=16'h278;
17'h18e2:	data_out=16'h43;
17'h18e3:	data_out=16'h800b;
17'h18e4:	data_out=16'h89;
17'h18e5:	data_out=16'h22c;
17'h18e6:	data_out=16'h143;
17'h18e7:	data_out=16'h8085;
17'h18e8:	data_out=16'hb;
17'h18e9:	data_out=16'h119;
17'h18ea:	data_out=16'h14;
17'h18eb:	data_out=16'h223;
17'h18ec:	data_out=16'h1a2;
17'h18ed:	data_out=16'h803a;
17'h18ee:	data_out=16'hd;
17'h18ef:	data_out=16'h2aa;
17'h18f0:	data_out=16'h5;
17'h18f1:	data_out=16'h8156;
17'h18f2:	data_out=16'h28c;
17'h18f3:	data_out=16'h236;
17'h18f4:	data_out=16'h412;
17'h18f5:	data_out=16'h39b;
17'h18f6:	data_out=16'h8073;
17'h18f7:	data_out=16'h1d1;
17'h18f8:	data_out=16'hcf;
17'h18f9:	data_out=16'h43;
17'h18fa:	data_out=16'h800c;
17'h18fb:	data_out=16'h13;
17'h18fc:	data_out=16'h80e7;
17'h18fd:	data_out=16'h8090;
17'h18fe:	data_out=16'h80cc;
17'h18ff:	data_out=16'he7;
17'h1900:	data_out=16'h801e;
17'h1901:	data_out=16'h1b;
17'h1902:	data_out=16'h80fb;
17'h1903:	data_out=16'h3f;
17'h1904:	data_out=16'h298;
17'h1905:	data_out=16'h18f;
17'h1906:	data_out=16'h8101;
17'h1907:	data_out=16'h80f5;
17'h1908:	data_out=16'h805a;
17'h1909:	data_out=16'h8116;
17'h190a:	data_out=16'hcc;
17'h190b:	data_out=16'hbe;
17'h190c:	data_out=16'h338;
17'h190d:	data_out=16'h8014;
17'h190e:	data_out=16'h803f;
17'h190f:	data_out=16'h8162;
17'h1910:	data_out=16'h8022;
17'h1911:	data_out=16'h1c4;
17'h1912:	data_out=16'h817b;
17'h1913:	data_out=16'ha7;
17'h1914:	data_out=16'h8168;
17'h1915:	data_out=16'h805e;
17'h1916:	data_out=16'h4;
17'h1917:	data_out=16'h8127;
17'h1918:	data_out=16'h8099;
17'h1919:	data_out=16'h18d;
17'h191a:	data_out=16'h354;
17'h191b:	data_out=16'h47;
17'h191c:	data_out=16'h3d;
17'h191d:	data_out=16'h20;
17'h191e:	data_out=16'h8172;
17'h191f:	data_out=16'h816f;
17'h1920:	data_out=16'h58;
17'h1921:	data_out=16'h803a;
17'h1922:	data_out=16'h8098;
17'h1923:	data_out=16'h8109;
17'h1924:	data_out=16'h8109;
17'h1925:	data_out=16'h88;
17'h1926:	data_out=16'h8134;
17'h1927:	data_out=16'h21;
17'h1928:	data_out=16'h8038;
17'h1929:	data_out=16'h6e;
17'h192a:	data_out=16'h814b;
17'h192b:	data_out=16'h19;
17'h192c:	data_out=16'h75;
17'h192d:	data_out=16'h1c6;
17'h192e:	data_out=16'h80cf;
17'h192f:	data_out=16'h88;
17'h1930:	data_out=16'h379;
17'h1931:	data_out=16'h130;
17'h1932:	data_out=16'h37a;
17'h1933:	data_out=16'h819e;
17'h1934:	data_out=16'hb3;
17'h1935:	data_out=16'h34a;
17'h1936:	data_out=16'h80b3;
17'h1937:	data_out=16'h8100;
17'h1938:	data_out=16'h8015;
17'h1939:	data_out=16'h81a5;
17'h193a:	data_out=16'h8170;
17'h193b:	data_out=16'h15c;
17'h193c:	data_out=16'h2e;
17'h193d:	data_out=16'h8000;
17'h193e:	data_out=16'h802e;
17'h193f:	data_out=16'h2a9;
17'h1940:	data_out=16'h1b;
17'h1941:	data_out=16'h8042;
17'h1942:	data_out=16'h1a4;
17'h1943:	data_out=16'h28;
17'h1944:	data_out=16'h1e7;
17'h1945:	data_out=16'h808c;
17'h1946:	data_out=16'hc;
17'h1947:	data_out=16'h814b;
17'h1948:	data_out=16'h80d1;
17'h1949:	data_out=16'h67;
17'h194a:	data_out=16'hf6;
17'h194b:	data_out=16'h28a;
17'h194c:	data_out=16'h5e;
17'h194d:	data_out=16'h80ac;
17'h194e:	data_out=16'ha2;
17'h194f:	data_out=16'hb0;
17'h1950:	data_out=16'h8067;
17'h1951:	data_out=16'h806d;
17'h1952:	data_out=16'h8101;
17'h1953:	data_out=16'h4f;
17'h1954:	data_out=16'h93;
17'h1955:	data_out=16'h80b4;
17'h1956:	data_out=16'h812d;
17'h1957:	data_out=16'h8135;
17'h1958:	data_out=16'h8088;
17'h1959:	data_out=16'h8045;
17'h195a:	data_out=16'h8023;
17'h195b:	data_out=16'h4d;
17'h195c:	data_out=16'hef;
17'h195d:	data_out=16'ha8;
17'h195e:	data_out=16'h183;
17'h195f:	data_out=16'h80c8;
17'h1960:	data_out=16'h19;
17'h1961:	data_out=16'h169;
17'h1962:	data_out=16'h8132;
17'h1963:	data_out=16'h8150;
17'h1964:	data_out=16'h8004;
17'h1965:	data_out=16'h20f;
17'h1966:	data_out=16'h173;
17'h1967:	data_out=16'h80c1;
17'h1968:	data_out=16'h8033;
17'h1969:	data_out=16'h8045;
17'h196a:	data_out=16'h8044;
17'h196b:	data_out=16'h1d9;
17'h196c:	data_out=16'h43;
17'h196d:	data_out=16'h8185;
17'h196e:	data_out=16'h8048;
17'h196f:	data_out=16'h1c1;
17'h1970:	data_out=16'h803f;
17'h1971:	data_out=16'h8222;
17'h1972:	data_out=16'h199;
17'h1973:	data_out=16'h13e;
17'h1974:	data_out=16'h37c;
17'h1975:	data_out=16'h218;
17'h1976:	data_out=16'h80a5;
17'h1977:	data_out=16'h165;
17'h1978:	data_out=16'h30;
17'h1979:	data_out=16'h813f;
17'h197a:	data_out=16'h816f;
17'h197b:	data_out=16'h803c;
17'h197c:	data_out=16'h8155;
17'h197d:	data_out=16'h8129;
17'h197e:	data_out=16'h810a;
17'h197f:	data_out=16'h46;
17'h1980:	data_out=16'h8059;
17'h1981:	data_out=16'h804e;
17'h1982:	data_out=16'h8104;
17'h1983:	data_out=16'h802a;
17'h1984:	data_out=16'h18c;
17'h1985:	data_out=16'h95;
17'h1986:	data_out=16'h8084;
17'h1987:	data_out=16'h8086;
17'h1988:	data_out=16'h8070;
17'h1989:	data_out=16'h809e;
17'h198a:	data_out=16'h2c;
17'h198b:	data_out=16'h801d;
17'h198c:	data_out=16'h268;
17'h198d:	data_out=16'h8048;
17'h198e:	data_out=16'h8033;
17'h198f:	data_out=16'h813f;
17'h1990:	data_out=16'h8051;
17'h1991:	data_out=16'hae;
17'h1992:	data_out=16'h813d;
17'h1993:	data_out=16'he;
17'h1994:	data_out=16'h813d;
17'h1995:	data_out=16'h8059;
17'h1996:	data_out=16'h803b;
17'h1997:	data_out=16'h8125;
17'h1998:	data_out=16'h8074;
17'h1999:	data_out=16'h101;
17'h199a:	data_out=16'h226;
17'h199b:	data_out=16'h8045;
17'h199c:	data_out=16'h804f;
17'h199d:	data_out=16'h8046;
17'h199e:	data_out=16'h8140;
17'h199f:	data_out=16'h80f7;
17'h19a0:	data_out=16'h8012;
17'h19a1:	data_out=16'h802a;
17'h19a2:	data_out=16'h806c;
17'h19a3:	data_out=16'h809a;
17'h19a4:	data_out=16'h8094;
17'h19a5:	data_out=16'h2b;
17'h19a6:	data_out=16'h80f1;
17'h19a7:	data_out=16'h8054;
17'h19a8:	data_out=16'h8035;
17'h19a9:	data_out=16'h4;
17'h19aa:	data_out=16'h8145;
17'h19ab:	data_out=16'h803c;
17'h19ac:	data_out=16'hb;
17'h19ad:	data_out=16'hda;
17'h19ae:	data_out=16'h80c6;
17'h19af:	data_out=16'hd;
17'h19b0:	data_out=16'h277;
17'h19b1:	data_out=16'h57;
17'h19b2:	data_out=16'h276;
17'h19b3:	data_out=16'h8155;
17'h19b4:	data_out=16'h24;
17'h19b5:	data_out=16'h208;
17'h19b6:	data_out=16'h80c3;
17'h19b7:	data_out=16'h8106;
17'h19b8:	data_out=16'h804e;
17'h19b9:	data_out=16'h8155;
17'h19ba:	data_out=16'h80db;
17'h19bb:	data_out=16'ha6;
17'h19bc:	data_out=16'h8068;
17'h19bd:	data_out=16'h8028;
17'h19be:	data_out=16'h8029;
17'h19bf:	data_out=16'h179;
17'h19c0:	data_out=16'h1b;
17'h19c1:	data_out=16'h8093;
17'h19c2:	data_out=16'h141;
17'h19c3:	data_out=16'h23;
17'h19c4:	data_out=16'hc8;
17'h19c5:	data_out=16'h8078;
17'h19c6:	data_out=16'h807f;
17'h19c7:	data_out=16'h80c9;
17'h19c8:	data_out=16'h808c;
17'h19c9:	data_out=16'h23;
17'h19ca:	data_out=16'h84;
17'h19cb:	data_out=16'h172;
17'h19cc:	data_out=16'h35;
17'h19cd:	data_out=16'h8077;
17'h19ce:	data_out=16'h4e;
17'h19cf:	data_out=16'h55;
17'h19d0:	data_out=16'h8052;
17'h19d1:	data_out=16'h80a6;
17'h19d2:	data_out=16'h808b;
17'h19d3:	data_out=16'h8043;
17'h19d4:	data_out=16'h0;
17'h19d5:	data_out=16'h80c8;
17'h19d6:	data_out=16'h811c;
17'h19d7:	data_out=16'h80db;
17'h19d8:	data_out=16'h80cc;
17'h19d9:	data_out=16'h803b;
17'h19da:	data_out=16'h809b;
17'h19db:	data_out=16'h8037;
17'h19dc:	data_out=16'h1a;
17'h19dd:	data_out=16'h1c;
17'h19de:	data_out=16'hac;
17'h19df:	data_out=16'h807e;
17'h19e0:	data_out=16'h806d;
17'h19e1:	data_out=16'h64;
17'h19e2:	data_out=16'h812b;
17'h19e3:	data_out=16'h8131;
17'h19e4:	data_out=16'h8070;
17'h19e5:	data_out=16'h152;
17'h19e6:	data_out=16'h10c;
17'h19e7:	data_out=16'h80a9;
17'h19e8:	data_out=16'h8037;
17'h19e9:	data_out=16'h806c;
17'h19ea:	data_out=16'h8039;
17'h19eb:	data_out=16'h113;
17'h19ec:	data_out=16'h8034;
17'h19ed:	data_out=16'h814b;
17'h19ee:	data_out=16'h8035;
17'h19ef:	data_out=16'h120;
17'h19f0:	data_out=16'h803c;
17'h19f1:	data_out=16'h81a5;
17'h19f2:	data_out=16'ha2;
17'h19f3:	data_out=16'h65;
17'h19f4:	data_out=16'h279;
17'h19f5:	data_out=16'hf1;
17'h19f6:	data_out=16'h8068;
17'h19f7:	data_out=16'hb7;
17'h19f8:	data_out=16'h2;
17'h19f9:	data_out=16'h8135;
17'h19fa:	data_out=16'h8144;
17'h19fb:	data_out=16'h802b;
17'h19fc:	data_out=16'h80b4;
17'h19fd:	data_out=16'h80be;
17'h19fe:	data_out=16'h808e;
17'h19ff:	data_out=16'h800c;
17'h1a00:	data_out=16'h8;
17'h1a01:	data_out=16'h8005;
17'h1a02:	data_out=16'h2;
17'h1a03:	data_out=16'h8007;
17'h1a04:	data_out=16'h5;
17'h1a05:	data_out=16'h0;
17'h1a06:	data_out=16'h7;
17'h1a07:	data_out=16'h9;
17'h1a08:	data_out=16'h8007;
17'h1a09:	data_out=16'h8005;
17'h1a0a:	data_out=16'h8008;
17'h1a0b:	data_out=16'h8008;
17'h1a0c:	data_out=16'h7;
17'h1a0d:	data_out=16'h1;
17'h1a0e:	data_out=16'h8009;
17'h1a0f:	data_out=16'h8;
17'h1a10:	data_out=16'h8009;
17'h1a11:	data_out=16'h2;
17'h1a12:	data_out=16'h8001;
17'h1a13:	data_out=16'h8004;
17'h1a14:	data_out=16'h8005;
17'h1a15:	data_out=16'h8008;
17'h1a16:	data_out=16'h4;
17'h1a17:	data_out=16'h8;
17'h1a18:	data_out=16'h9;
17'h1a19:	data_out=16'h8001;
17'h1a1a:	data_out=16'h4;
17'h1a1b:	data_out=16'h9;
17'h1a1c:	data_out=16'h7;
17'h1a1d:	data_out=16'h8001;
17'h1a1e:	data_out=16'h8006;
17'h1a1f:	data_out=16'h6;
17'h1a20:	data_out=16'h4;
17'h1a21:	data_out=16'h5;
17'h1a22:	data_out=16'h8;
17'h1a23:	data_out=16'h8001;
17'h1a24:	data_out=16'h8004;
17'h1a25:	data_out=16'h7;
17'h1a26:	data_out=16'h8001;
17'h1a27:	data_out=16'h8001;
17'h1a28:	data_out=16'h8008;
17'h1a29:	data_out=16'h8001;
17'h1a2a:	data_out=16'h8000;
17'h1a2b:	data_out=16'h8;
17'h1a2c:	data_out=16'h8008;
17'h1a2d:	data_out=16'h8000;
17'h1a2e:	data_out=16'h7;
17'h1a2f:	data_out=16'h8008;
17'h1a30:	data_out=16'h8007;
17'h1a31:	data_out=16'h8004;
17'h1a32:	data_out=16'h8003;
17'h1a33:	data_out=16'h8003;
17'h1a34:	data_out=16'h8002;
17'h1a35:	data_out=16'h8008;
17'h1a36:	data_out=16'h8004;
17'h1a37:	data_out=16'h8002;
17'h1a38:	data_out=16'h8000;
17'h1a39:	data_out=16'h8009;
17'h1a3a:	data_out=16'h8003;
17'h1a3b:	data_out=16'h8002;
17'h1a3c:	data_out=16'h8001;
17'h1a3d:	data_out=16'h0;
17'h1a3e:	data_out=16'h8006;
17'h1a3f:	data_out=16'h8006;
17'h1a40:	data_out=16'h8004;
17'h1a41:	data_out=16'h8006;
17'h1a42:	data_out=16'h2;
17'h1a43:	data_out=16'h2;
17'h1a44:	data_out=16'h8009;
17'h1a45:	data_out=16'h8008;
17'h1a46:	data_out=16'h8009;
17'h1a47:	data_out=16'h8008;
17'h1a48:	data_out=16'h1;
17'h1a49:	data_out=16'h0;
17'h1a4a:	data_out=16'h8009;
17'h1a4b:	data_out=16'h1;
17'h1a4c:	data_out=16'h8009;
17'h1a4d:	data_out=16'h8;
17'h1a4e:	data_out=16'h3;
17'h1a4f:	data_out=16'h8007;
17'h1a50:	data_out=16'h8005;
17'h1a51:	data_out=16'h9;
17'h1a52:	data_out=16'h8001;
17'h1a53:	data_out=16'h2;
17'h1a54:	data_out=16'h8008;
17'h1a55:	data_out=16'h5;
17'h1a56:	data_out=16'h9;
17'h1a57:	data_out=16'h0;
17'h1a58:	data_out=16'h5;
17'h1a59:	data_out=16'h8003;
17'h1a5a:	data_out=16'h7;
17'h1a5b:	data_out=16'h8005;
17'h1a5c:	data_out=16'h6;
17'h1a5d:	data_out=16'h8008;
17'h1a5e:	data_out=16'h8002;
17'h1a5f:	data_out=16'h8007;
17'h1a60:	data_out=16'h8005;
17'h1a61:	data_out=16'h8008;
17'h1a62:	data_out=16'h5;
17'h1a63:	data_out=16'h8005;
17'h1a64:	data_out=16'h8007;
17'h1a65:	data_out=16'h5;
17'h1a66:	data_out=16'h8003;
17'h1a67:	data_out=16'h2;
17'h1a68:	data_out=16'h8004;
17'h1a69:	data_out=16'h8003;
17'h1a6a:	data_out=16'h8005;
17'h1a6b:	data_out=16'h8003;
17'h1a6c:	data_out=16'h8004;
17'h1a6d:	data_out=16'h7;
17'h1a6e:	data_out=16'h8001;
17'h1a6f:	data_out=16'h8000;
17'h1a70:	data_out=16'h6;
17'h1a71:	data_out=16'h8;
17'h1a72:	data_out=16'h8007;
17'h1a73:	data_out=16'h7;
17'h1a74:	data_out=16'h3;
17'h1a75:	data_out=16'h8007;
17'h1a76:	data_out=16'h8002;
17'h1a77:	data_out=16'h8001;
17'h1a78:	data_out=16'h8001;
17'h1a79:	data_out=16'h8004;
17'h1a7a:	data_out=16'h4;
17'h1a7b:	data_out=16'h8004;
17'h1a7c:	data_out=16'h8003;
17'h1a7d:	data_out=16'h8007;
17'h1a7e:	data_out=16'h8002;
17'h1a7f:	data_out=16'h2;
17'h1a80:	data_out=16'h8006;
17'h1a81:	data_out=16'h8006;
17'h1a82:	data_out=16'h6;
17'h1a83:	data_out=16'h8004;
17'h1a84:	data_out=16'h8;
17'h1a85:	data_out=16'h8007;
17'h1a86:	data_out=16'h7;
17'h1a87:	data_out=16'h8005;
17'h1a88:	data_out=16'h8000;
17'h1a89:	data_out=16'h8007;
17'h1a8a:	data_out=16'h1;
17'h1a8b:	data_out=16'h5;
17'h1a8c:	data_out=16'h9;
17'h1a8d:	data_out=16'h8009;
17'h1a8e:	data_out=16'h8005;
17'h1a8f:	data_out=16'h6;
17'h1a90:	data_out=16'h8;
17'h1a91:	data_out=16'h8002;
17'h1a92:	data_out=16'h4;
17'h1a93:	data_out=16'h2;
17'h1a94:	data_out=16'h8000;
17'h1a95:	data_out=16'h8007;
17'h1a96:	data_out=16'h8008;
17'h1a97:	data_out=16'h8;
17'h1a98:	data_out=16'h8002;
17'h1a99:	data_out=16'h6;
17'h1a9a:	data_out=16'h8006;
17'h1a9b:	data_out=16'h4;
17'h1a9c:	data_out=16'h8;
17'h1a9d:	data_out=16'h2;
17'h1a9e:	data_out=16'h8003;
17'h1a9f:	data_out=16'h8007;
17'h1aa0:	data_out=16'h5;
17'h1aa1:	data_out=16'h8007;
17'h1aa2:	data_out=16'h8002;
17'h1aa3:	data_out=16'h4;
17'h1aa4:	data_out=16'h8004;
17'h1aa5:	data_out=16'h8004;
17'h1aa6:	data_out=16'h8;
17'h1aa7:	data_out=16'h5;
17'h1aa8:	data_out=16'h8002;
17'h1aa9:	data_out=16'h0;
17'h1aaa:	data_out=16'h1;
17'h1aab:	data_out=16'h8002;
17'h1aac:	data_out=16'h1;
17'h1aad:	data_out=16'h5;
17'h1aae:	data_out=16'h8005;
17'h1aaf:	data_out=16'h8001;
17'h1ab0:	data_out=16'h8006;
17'h1ab1:	data_out=16'h7;
17'h1ab2:	data_out=16'h8007;
17'h1ab3:	data_out=16'h2;
17'h1ab4:	data_out=16'h8009;
17'h1ab5:	data_out=16'h8006;
17'h1ab6:	data_out=16'h1;
17'h1ab7:	data_out=16'h8002;
17'h1ab8:	data_out=16'h9;
17'h1ab9:	data_out=16'h4;
17'h1aba:	data_out=16'h8007;
17'h1abb:	data_out=16'h8;
17'h1abc:	data_out=16'h8003;
17'h1abd:	data_out=16'h8001;
17'h1abe:	data_out=16'h8008;
17'h1abf:	data_out=16'h8007;
17'h1ac0:	data_out=16'h1;
17'h1ac1:	data_out=16'h8001;
17'h1ac2:	data_out=16'h5;
17'h1ac3:	data_out=16'h7;
17'h1ac4:	data_out=16'h4;
17'h1ac5:	data_out=16'h4;
17'h1ac6:	data_out=16'h2;
17'h1ac7:	data_out=16'h8006;
17'h1ac8:	data_out=16'h8005;
17'h1ac9:	data_out=16'h8006;
17'h1aca:	data_out=16'h1;
17'h1acb:	data_out=16'h5;
17'h1acc:	data_out=16'h8;
17'h1acd:	data_out=16'h4;
17'h1ace:	data_out=16'h8004;
17'h1acf:	data_out=16'h8007;
17'h1ad0:	data_out=16'h2;
17'h1ad1:	data_out=16'h8003;
17'h1ad2:	data_out=16'h4;
17'h1ad3:	data_out=16'h2;
17'h1ad4:	data_out=16'h1;
17'h1ad5:	data_out=16'h8004;
17'h1ad6:	data_out=16'h8009;
17'h1ad7:	data_out=16'h0;
17'h1ad8:	data_out=16'h8009;
17'h1ad9:	data_out=16'h8007;
17'h1ada:	data_out=16'h8001;
17'h1adb:	data_out=16'h8003;
17'h1adc:	data_out=16'h1;
17'h1add:	data_out=16'h8000;
17'h1ade:	data_out=16'h8001;
17'h1adf:	data_out=16'h8007;
17'h1ae0:	data_out=16'h8;
17'h1ae1:	data_out=16'h8005;
17'h1ae2:	data_out=16'h9;
17'h1ae3:	data_out=16'h3;
17'h1ae4:	data_out=16'h9;
17'h1ae5:	data_out=16'h2;
17'h1ae6:	data_out=16'h6;
17'h1ae7:	data_out=16'h8005;
17'h1ae8:	data_out=16'h5;
17'h1ae9:	data_out=16'h8003;
17'h1aea:	data_out=16'h8009;
17'h1aeb:	data_out=16'h4;
17'h1aec:	data_out=16'h8008;
17'h1aed:	data_out=16'h8004;
17'h1aee:	data_out=16'h6;
17'h1aef:	data_out=16'h3;
17'h1af0:	data_out=16'h2;
17'h1af1:	data_out=16'h1;
17'h1af2:	data_out=16'h8003;
17'h1af3:	data_out=16'h8006;
17'h1af4:	data_out=16'h6;
17'h1af5:	data_out=16'h8003;
17'h1af6:	data_out=16'h3;
17'h1af7:	data_out=16'h7;
17'h1af8:	data_out=16'h8001;
17'h1af9:	data_out=16'h8007;
17'h1afa:	data_out=16'h8005;
17'h1afb:	data_out=16'h9;
17'h1afc:	data_out=16'h2;
17'h1afd:	data_out=16'h3;
17'h1afe:	data_out=16'h8007;
17'h1aff:	data_out=16'h1;
17'h1b00:	data_out=16'h8;
17'h1b01:	data_out=16'h8007;
17'h1b02:	data_out=16'h8006;
17'h1b03:	data_out=16'h7;
17'h1b04:	data_out=16'h4;
17'h1b05:	data_out=16'h9;
17'h1b06:	data_out=16'h8006;
17'h1b07:	data_out=16'h8000;
17'h1b08:	data_out=16'h8003;
17'h1b09:	data_out=16'h8006;
17'h1b0a:	data_out=16'h8005;
17'h1b0b:	data_out=16'h8002;
17'h1b0c:	data_out=16'h8001;
17'h1b0d:	data_out=16'h8008;
17'h1b0e:	data_out=16'h8008;
17'h1b0f:	data_out=16'h8007;
17'h1b10:	data_out=16'h2;
17'h1b11:	data_out=16'h8002;
17'h1b12:	data_out=16'h8004;
17'h1b13:	data_out=16'h8001;
17'h1b14:	data_out=16'h4;
17'h1b15:	data_out=16'h8;
17'h1b16:	data_out=16'h8003;
17'h1b17:	data_out=16'h8006;
17'h1b18:	data_out=16'h8008;
17'h1b19:	data_out=16'h1;
17'h1b1a:	data_out=16'h8006;
17'h1b1b:	data_out=16'h3;
17'h1b1c:	data_out=16'h8005;
17'h1b1d:	data_out=16'h8004;
17'h1b1e:	data_out=16'h8005;
17'h1b1f:	data_out=16'h8007;
17'h1b20:	data_out=16'h8002;
17'h1b21:	data_out=16'h8002;
17'h1b22:	data_out=16'h8009;
17'h1b23:	data_out=16'h8007;
17'h1b24:	data_out=16'h8002;
17'h1b25:	data_out=16'h8006;
17'h1b26:	data_out=16'h2;
17'h1b27:	data_out=16'h4;
17'h1b28:	data_out=16'h8003;
17'h1b29:	data_out=16'h6;
17'h1b2a:	data_out=16'h8008;
17'h1b2b:	data_out=16'h5;
17'h1b2c:	data_out=16'h7;
17'h1b2d:	data_out=16'h8006;
17'h1b2e:	data_out=16'h7;
17'h1b2f:	data_out=16'h8000;
17'h1b30:	data_out=16'h1;
17'h1b31:	data_out=16'h8006;
17'h1b32:	data_out=16'h8;
17'h1b33:	data_out=16'h8004;
17'h1b34:	data_out=16'h8008;
17'h1b35:	data_out=16'h8004;
17'h1b36:	data_out=16'h8001;
17'h1b37:	data_out=16'h8006;
17'h1b38:	data_out=16'h5;
17'h1b39:	data_out=16'h2;
17'h1b3a:	data_out=16'h6;
17'h1b3b:	data_out=16'h9;
17'h1b3c:	data_out=16'h7;
17'h1b3d:	data_out=16'h8009;
17'h1b3e:	data_out=16'h8007;
17'h1b3f:	data_out=16'h8004;
17'h1b40:	data_out=16'h8001;
17'h1b41:	data_out=16'h8007;
17'h1b42:	data_out=16'h8003;
17'h1b43:	data_out=16'h6;
17'h1b44:	data_out=16'h8003;
17'h1b45:	data_out=16'h8;
17'h1b46:	data_out=16'h0;
17'h1b47:	data_out=16'h3;
17'h1b48:	data_out=16'h5;
17'h1b49:	data_out=16'h2;
17'h1b4a:	data_out=16'h8001;
17'h1b4b:	data_out=16'h2;
17'h1b4c:	data_out=16'h5;
17'h1b4d:	data_out=16'h8003;
17'h1b4e:	data_out=16'h8007;
17'h1b4f:	data_out=16'h8004;
17'h1b50:	data_out=16'h8000;
17'h1b51:	data_out=16'h8008;
17'h1b52:	data_out=16'h1;
17'h1b53:	data_out=16'h1;
17'h1b54:	data_out=16'h8004;
17'h1b55:	data_out=16'h9;
17'h1b56:	data_out=16'h4;
17'h1b57:	data_out=16'h8007;
17'h1b58:	data_out=16'h2;
17'h1b59:	data_out=16'h1;
17'h1b5a:	data_out=16'h8007;
17'h1b5b:	data_out=16'h8001;
17'h1b5c:	data_out=16'h2;
17'h1b5d:	data_out=16'h8005;
17'h1b5e:	data_out=16'h4;
17'h1b5f:	data_out=16'h8009;
17'h1b60:	data_out=16'h8003;
17'h1b61:	data_out=16'h8008;
17'h1b62:	data_out=16'h6;
17'h1b63:	data_out=16'h3;
17'h1b64:	data_out=16'h8009;
17'h1b65:	data_out=16'h8003;
17'h1b66:	data_out=16'h8003;
17'h1b67:	data_out=16'h5;
17'h1b68:	data_out=16'h7;
17'h1b69:	data_out=16'h5;
17'h1b6a:	data_out=16'h8002;
17'h1b6b:	data_out=16'h3;
17'h1b6c:	data_out=16'h8007;
17'h1b6d:	data_out=16'h8000;
17'h1b6e:	data_out=16'h8;
17'h1b6f:	data_out=16'h2;
17'h1b70:	data_out=16'h1;
17'h1b71:	data_out=16'h0;
17'h1b72:	data_out=16'h8006;
17'h1b73:	data_out=16'h6;
17'h1b74:	data_out=16'h0;
17'h1b75:	data_out=16'h8;
17'h1b76:	data_out=16'h8;
17'h1b77:	data_out=16'h8007;
17'h1b78:	data_out=16'h8001;
17'h1b79:	data_out=16'h8009;
17'h1b7a:	data_out=16'h1;
17'h1b7b:	data_out=16'h8008;
17'h1b7c:	data_out=16'h8005;
17'h1b7d:	data_out=16'h8004;
17'h1b7e:	data_out=16'h8008;
17'h1b7f:	data_out=16'h2;
17'h1b80:	data_out=16'h8003;
17'h1b81:	data_out=16'h7;
17'h1b82:	data_out=16'h8004;
17'h1b83:	data_out=16'h8002;
17'h1b84:	data_out=16'h8006;
17'h1b85:	data_out=16'h2;
17'h1b86:	data_out=16'h8006;
17'h1b87:	data_out=16'h8008;
17'h1b88:	data_out=16'h8002;
17'h1b89:	data_out=16'h1;
17'h1b8a:	data_out=16'h4;
17'h1b8b:	data_out=16'h0;
17'h1b8c:	data_out=16'h8009;
17'h1b8d:	data_out=16'h3;
17'h1b8e:	data_out=16'h8007;
17'h1b8f:	data_out=16'h1;
17'h1b90:	data_out=16'h8005;
17'h1b91:	data_out=16'h8004;
17'h1b92:	data_out=16'h8002;
17'h1b93:	data_out=16'h4;
17'h1b94:	data_out=16'h8005;
17'h1b95:	data_out=16'h8003;
17'h1b96:	data_out=16'h5;
17'h1b97:	data_out=16'h3;
17'h1b98:	data_out=16'h8003;
17'h1b99:	data_out=16'h8003;
17'h1b9a:	data_out=16'h4;
17'h1b9b:	data_out=16'h2;
17'h1b9c:	data_out=16'h2;
17'h1b9d:	data_out=16'h5;
17'h1b9e:	data_out=16'h8006;
17'h1b9f:	data_out=16'h9;
17'h1ba0:	data_out=16'h3;
17'h1ba1:	data_out=16'h8000;
17'h1ba2:	data_out=16'h8003;
17'h1ba3:	data_out=16'h6;
17'h1ba4:	data_out=16'h8008;
17'h1ba5:	data_out=16'h0;
17'h1ba6:	data_out=16'h7;
17'h1ba7:	data_out=16'h8001;
17'h1ba8:	data_out=16'h8008;
17'h1ba9:	data_out=16'h3;
17'h1baa:	data_out=16'h9;
17'h1bab:	data_out=16'h8008;
17'h1bac:	data_out=16'h8003;
17'h1bad:	data_out=16'h8008;
17'h1bae:	data_out=16'h2;
17'h1baf:	data_out=16'h1;
17'h1bb0:	data_out=16'h8002;
17'h1bb1:	data_out=16'h8009;
17'h1bb2:	data_out=16'h8005;
17'h1bb3:	data_out=16'h2;
17'h1bb4:	data_out=16'h8003;
17'h1bb5:	data_out=16'h8008;
17'h1bb6:	data_out=16'h8004;
17'h1bb7:	data_out=16'h3;
17'h1bb8:	data_out=16'h8002;
17'h1bb9:	data_out=16'h9;
17'h1bba:	data_out=16'h8004;
17'h1bbb:	data_out=16'h8009;
17'h1bbc:	data_out=16'h5;
17'h1bbd:	data_out=16'h8001;
17'h1bbe:	data_out=16'h8009;
17'h1bbf:	data_out=16'h8001;
17'h1bc0:	data_out=16'h8;
17'h1bc1:	data_out=16'h8002;
17'h1bc2:	data_out=16'h8005;
17'h1bc3:	data_out=16'h8009;
17'h1bc4:	data_out=16'h7;
17'h1bc5:	data_out=16'h8006;
17'h1bc6:	data_out=16'h8000;
17'h1bc7:	data_out=16'h7;
17'h1bc8:	data_out=16'h6;
17'h1bc9:	data_out=16'h8001;
17'h1bca:	data_out=16'h9;
17'h1bcb:	data_out=16'h8006;
17'h1bcc:	data_out=16'h1;
17'h1bcd:	data_out=16'h2;
17'h1bce:	data_out=16'h3;
17'h1bcf:	data_out=16'h8;
17'h1bd0:	data_out=16'h2;
17'h1bd1:	data_out=16'h8;
17'h1bd2:	data_out=16'h1;
17'h1bd3:	data_out=16'h8;
17'h1bd4:	data_out=16'h9;
17'h1bd5:	data_out=16'h6;
17'h1bd6:	data_out=16'h2;
17'h1bd7:	data_out=16'h8002;
17'h1bd8:	data_out=16'h5;
17'h1bd9:	data_out=16'h7;
17'h1bda:	data_out=16'h8002;
17'h1bdb:	data_out=16'h1;
17'h1bdc:	data_out=16'h8003;
17'h1bdd:	data_out=16'h8002;
17'h1bde:	data_out=16'h8009;
17'h1bdf:	data_out=16'h8004;
17'h1be0:	data_out=16'h5;
17'h1be1:	data_out=16'h8005;
17'h1be2:	data_out=16'h8004;
17'h1be3:	data_out=16'h3;
17'h1be4:	data_out=16'h8002;
17'h1be5:	data_out=16'h5;
17'h1be6:	data_out=16'h1;
17'h1be7:	data_out=16'h8005;
17'h1be8:	data_out=16'h8004;
17'h1be9:	data_out=16'h0;
17'h1bea:	data_out=16'h8003;
17'h1beb:	data_out=16'h6;
17'h1bec:	data_out=16'h8007;
17'h1bed:	data_out=16'h8008;
17'h1bee:	data_out=16'h5;
17'h1bef:	data_out=16'h3;
17'h1bf0:	data_out=16'h9;
17'h1bf1:	data_out=16'h8004;
17'h1bf2:	data_out=16'h2;
17'h1bf3:	data_out=16'h8;
17'h1bf4:	data_out=16'h8008;
17'h1bf5:	data_out=16'h8005;
17'h1bf6:	data_out=16'h8003;
17'h1bf7:	data_out=16'h7;
17'h1bf8:	data_out=16'h8008;
17'h1bf9:	data_out=16'h4;
17'h1bfa:	data_out=16'h8001;
17'h1bfb:	data_out=16'h8001;
17'h1bfc:	data_out=16'h8007;
17'h1bfd:	data_out=16'h8001;
17'h1bfe:	data_out=16'h4;
17'h1bff:	data_out=16'h7;
17'h1c00:	data_out=16'h4;
17'h1c01:	data_out=16'h8009;
17'h1c02:	data_out=16'h1;
17'h1c03:	data_out=16'h8007;
17'h1c04:	data_out=16'h6;
17'h1c05:	data_out=16'h8008;
17'h1c06:	data_out=16'h8003;
17'h1c07:	data_out=16'h8008;
17'h1c08:	data_out=16'h2;
17'h1c09:	data_out=16'h4;
17'h1c0a:	data_out=16'h7;
17'h1c0b:	data_out=16'h3;
17'h1c0c:	data_out=16'h5;
17'h1c0d:	data_out=16'h3;
17'h1c0e:	data_out=16'h8002;
17'h1c0f:	data_out=16'h4;
17'h1c10:	data_out=16'h8;
17'h1c11:	data_out=16'h9;
17'h1c12:	data_out=16'h3;
17'h1c13:	data_out=16'h8009;
17'h1c14:	data_out=16'h8006;
17'h1c15:	data_out=16'h8009;
17'h1c16:	data_out=16'h7;
17'h1c17:	data_out=16'h8004;
17'h1c18:	data_out=16'h4;
17'h1c19:	data_out=16'h8003;
17'h1c1a:	data_out=16'h4;
17'h1c1b:	data_out=16'h6;
17'h1c1c:	data_out=16'h6;
17'h1c1d:	data_out=16'h8002;
17'h1c1e:	data_out=16'h5;
17'h1c1f:	data_out=16'h1;
17'h1c20:	data_out=16'h8002;
17'h1c21:	data_out=16'h8004;
17'h1c22:	data_out=16'h3;
17'h1c23:	data_out=16'h8005;
17'h1c24:	data_out=16'h8002;
17'h1c25:	data_out=16'h8009;
17'h1c26:	data_out=16'h8004;
17'h1c27:	data_out=16'h8;
17'h1c28:	data_out=16'h4;
17'h1c29:	data_out=16'h8006;
17'h1c2a:	data_out=16'h3;
17'h1c2b:	data_out=16'h8000;
17'h1c2c:	data_out=16'h6;
17'h1c2d:	data_out=16'h8009;
17'h1c2e:	data_out=16'h8005;
17'h1c2f:	data_out=16'h5;
17'h1c30:	data_out=16'h9;
17'h1c31:	data_out=16'h7;
17'h1c32:	data_out=16'h5;
17'h1c33:	data_out=16'h8006;
17'h1c34:	data_out=16'h8;
17'h1c35:	data_out=16'h3;
17'h1c36:	data_out=16'h8001;
17'h1c37:	data_out=16'h3;
17'h1c38:	data_out=16'h8009;
17'h1c39:	data_out=16'h8007;
17'h1c3a:	data_out=16'h8000;
17'h1c3b:	data_out=16'h7;
17'h1c3c:	data_out=16'h1;
17'h1c3d:	data_out=16'h8005;
17'h1c3e:	data_out=16'h8002;
17'h1c3f:	data_out=16'h8;
17'h1c40:	data_out=16'h1;
17'h1c41:	data_out=16'h8008;
17'h1c42:	data_out=16'h8006;
17'h1c43:	data_out=16'h8;
17'h1c44:	data_out=16'h8007;
17'h1c45:	data_out=16'h8000;
17'h1c46:	data_out=16'h7;
17'h1c47:	data_out=16'h6;
17'h1c48:	data_out=16'h3;
17'h1c49:	data_out=16'h0;
17'h1c4a:	data_out=16'h8004;
17'h1c4b:	data_out=16'h0;
17'h1c4c:	data_out=16'h0;
17'h1c4d:	data_out=16'h0;
17'h1c4e:	data_out=16'h8004;
17'h1c4f:	data_out=16'h0;
17'h1c50:	data_out=16'h8001;
17'h1c51:	data_out=16'h8008;
17'h1c52:	data_out=16'h3;
17'h1c53:	data_out=16'h8003;
17'h1c54:	data_out=16'h4;
17'h1c55:	data_out=16'h8007;
17'h1c56:	data_out=16'h9;
17'h1c57:	data_out=16'h5;
17'h1c58:	data_out=16'h8005;
17'h1c59:	data_out=16'h8000;
17'h1c5a:	data_out=16'h2;
17'h1c5b:	data_out=16'h5;
17'h1c5c:	data_out=16'h4;
17'h1c5d:	data_out=16'h8008;
17'h1c5e:	data_out=16'h4;
17'h1c5f:	data_out=16'h8004;
17'h1c60:	data_out=16'h8007;
17'h1c61:	data_out=16'h7;
17'h1c62:	data_out=16'h8006;
17'h1c63:	data_out=16'h8005;
17'h1c64:	data_out=16'h8002;
17'h1c65:	data_out=16'h8008;
17'h1c66:	data_out=16'h8009;
17'h1c67:	data_out=16'h8008;
17'h1c68:	data_out=16'h2;
17'h1c69:	data_out=16'h8003;
17'h1c6a:	data_out=16'h1;
17'h1c6b:	data_out=16'h8007;
17'h1c6c:	data_out=16'h7;
17'h1c6d:	data_out=16'h6;
17'h1c6e:	data_out=16'h2;
17'h1c6f:	data_out=16'h8004;
17'h1c70:	data_out=16'h7;
17'h1c71:	data_out=16'h8004;
17'h1c72:	data_out=16'h3;
17'h1c73:	data_out=16'h3;
17'h1c74:	data_out=16'h8002;
17'h1c75:	data_out=16'h2;
17'h1c76:	data_out=16'h8002;
17'h1c77:	data_out=16'h2;
17'h1c78:	data_out=16'h8007;
17'h1c79:	data_out=16'h8008;
17'h1c7a:	data_out=16'h8002;
17'h1c7b:	data_out=16'h7;
17'h1c7c:	data_out=16'h8008;
17'h1c7d:	data_out=16'h8007;
17'h1c7e:	data_out=16'h8007;
17'h1c7f:	data_out=16'h8005;
17'h1c80:	data_out=16'h9;
17'h1c81:	data_out=16'h8003;
17'h1c82:	data_out=16'h8002;
17'h1c83:	data_out=16'h8003;
17'h1c84:	data_out=16'h8002;
17'h1c85:	data_out=16'h8001;
17'h1c86:	data_out=16'h8002;
17'h1c87:	data_out=16'h9;
17'h1c88:	data_out=16'h5;
17'h1c89:	data_out=16'h9;
17'h1c8a:	data_out=16'h8007;
17'h1c8b:	data_out=16'h3;
17'h1c8c:	data_out=16'h6;
17'h1c8d:	data_out=16'h4;
17'h1c8e:	data_out=16'h8;
17'h1c8f:	data_out=16'h4;
17'h1c90:	data_out=16'h8009;
17'h1c91:	data_out=16'h2;
17'h1c92:	data_out=16'h8003;
17'h1c93:	data_out=16'h8002;
17'h1c94:	data_out=16'h8005;
17'h1c95:	data_out=16'h5;
17'h1c96:	data_out=16'h8008;
17'h1c97:	data_out=16'h8003;
17'h1c98:	data_out=16'h6;
17'h1c99:	data_out=16'h8001;
17'h1c9a:	data_out=16'h8005;
17'h1c9b:	data_out=16'h7;
17'h1c9c:	data_out=16'h1;
17'h1c9d:	data_out=16'h8003;
17'h1c9e:	data_out=16'h8007;
17'h1c9f:	data_out=16'h1;
17'h1ca0:	data_out=16'h3;
17'h1ca1:	data_out=16'h0;
17'h1ca2:	data_out=16'h8;
17'h1ca3:	data_out=16'h8008;
17'h1ca4:	data_out=16'h8;
17'h1ca5:	data_out=16'h8003;
17'h1ca6:	data_out=16'h8008;
17'h1ca7:	data_out=16'h5;
17'h1ca8:	data_out=16'h8004;
17'h1ca9:	data_out=16'h8006;
17'h1caa:	data_out=16'h8002;
17'h1cab:	data_out=16'h8007;
17'h1cac:	data_out=16'h7;
17'h1cad:	data_out=16'h8003;
17'h1cae:	data_out=16'h6;
17'h1caf:	data_out=16'h8;
17'h1cb0:	data_out=16'h8;
17'h1cb1:	data_out=16'h8006;
17'h1cb2:	data_out=16'h8003;
17'h1cb3:	data_out=16'h8006;
17'h1cb4:	data_out=16'h8;
17'h1cb5:	data_out=16'h8002;
17'h1cb6:	data_out=16'h1;
17'h1cb7:	data_out=16'h5;
17'h1cb8:	data_out=16'h6;
17'h1cb9:	data_out=16'h4;
17'h1cba:	data_out=16'h3;
17'h1cbb:	data_out=16'h8002;
17'h1cbc:	data_out=16'h8008;
17'h1cbd:	data_out=16'h5;
17'h1cbe:	data_out=16'h8;
17'h1cbf:	data_out=16'h5;
17'h1cc0:	data_out=16'h8004;
17'h1cc1:	data_out=16'h7;
17'h1cc2:	data_out=16'h6;
17'h1cc3:	data_out=16'h8005;
17'h1cc4:	data_out=16'h8006;
17'h1cc5:	data_out=16'h7;
17'h1cc6:	data_out=16'h9;
17'h1cc7:	data_out=16'h8001;
17'h1cc8:	data_out=16'h8007;
17'h1cc9:	data_out=16'h8002;
17'h1cca:	data_out=16'h1;
17'h1ccb:	data_out=16'h9;
17'h1ccc:	data_out=16'h4;
17'h1ccd:	data_out=16'h8002;
17'h1cce:	data_out=16'h8;
17'h1ccf:	data_out=16'h4;
17'h1cd0:	data_out=16'h1;
17'h1cd1:	data_out=16'h8004;
17'h1cd2:	data_out=16'h7;
17'h1cd3:	data_out=16'h8000;
17'h1cd4:	data_out=16'h3;
17'h1cd5:	data_out=16'h8002;
17'h1cd6:	data_out=16'h8004;
17'h1cd7:	data_out=16'h8000;
17'h1cd8:	data_out=16'h8006;
17'h1cd9:	data_out=16'h8;
17'h1cda:	data_out=16'h7;
17'h1cdb:	data_out=16'h8005;
17'h1cdc:	data_out=16'h3;
17'h1cdd:	data_out=16'h6;
17'h1cde:	data_out=16'h8009;
17'h1cdf:	data_out=16'h9;
17'h1ce0:	data_out=16'h3;
17'h1ce1:	data_out=16'h6;
17'h1ce2:	data_out=16'h8005;
17'h1ce3:	data_out=16'h6;
17'h1ce4:	data_out=16'h5;
17'h1ce5:	data_out=16'h8005;
17'h1ce6:	data_out=16'h8003;
17'h1ce7:	data_out=16'h6;
17'h1ce8:	data_out=16'h2;
17'h1ce9:	data_out=16'h7;
17'h1cea:	data_out=16'h6;
17'h1ceb:	data_out=16'h8003;
17'h1cec:	data_out=16'h8004;
17'h1ced:	data_out=16'h5;
17'h1cee:	data_out=16'h8008;
17'h1cef:	data_out=16'h6;
17'h1cf0:	data_out=16'h8009;
17'h1cf1:	data_out=16'h8;
17'h1cf2:	data_out=16'h8003;
17'h1cf3:	data_out=16'h3;
17'h1cf4:	data_out=16'h8003;
17'h1cf5:	data_out=16'h1;
17'h1cf6:	data_out=16'h8007;
17'h1cf7:	data_out=16'h8000;
17'h1cf8:	data_out=16'h8000;
17'h1cf9:	data_out=16'h8009;
17'h1cfa:	data_out=16'h4;
17'h1cfb:	data_out=16'h8006;
17'h1cfc:	data_out=16'h6;
17'h1cfd:	data_out=16'h4;
17'h1cfe:	data_out=16'h8006;
17'h1cff:	data_out=16'h8000;
17'h1d00:	data_out=16'h6;
17'h1d01:	data_out=16'h9;
17'h1d02:	data_out=16'ha;
17'h1d03:	data_out=16'hb;
17'h1d04:	data_out=16'hc;
17'h1d05:	data_out=16'h13;
17'h1d06:	data_out=16'h6;
17'h1d07:	data_out=16'h3;
17'h1d08:	data_out=16'h8;
17'h1d09:	data_out=16'hd;
17'h1d0a:	data_out=16'ha;
17'h1d0b:	data_out=16'h10;
17'h1d0c:	data_out=16'hc;
17'h1d0d:	data_out=16'he;
17'h1d0e:	data_out=16'h6;
17'h1d0f:	data_out=16'h11;
17'h1d10:	data_out=16'h9;
17'h1d11:	data_out=16'h11;
17'h1d12:	data_out=16'hd;
17'h1d13:	data_out=16'h15;
17'h1d14:	data_out=16'h12;
17'h1d15:	data_out=16'h9;
17'h1d16:	data_out=16'h9;
17'h1d17:	data_out=16'h1c;
17'h1d18:	data_out=16'h6;
17'h1d19:	data_out=16'h8005;
17'h1d1a:	data_out=16'h4;
17'h1d1b:	data_out=16'hc;
17'h1d1c:	data_out=16'h16;
17'h1d1d:	data_out=16'hb;
17'h1d1e:	data_out=16'h16;
17'h1d1f:	data_out=16'hb;
17'h1d20:	data_out=16'h13;
17'h1d21:	data_out=16'h8001;
17'h1d22:	data_out=16'h12;
17'h1d23:	data_out=16'h8000;
17'h1d24:	data_out=16'hb;
17'h1d25:	data_out=16'he;
17'h1d26:	data_out=16'h4;
17'h1d27:	data_out=16'hc;
17'h1d28:	data_out=16'hb;
17'h1d29:	data_out=16'h12;
17'h1d2a:	data_out=16'h5;
17'h1d2b:	data_out=16'h7;
17'h1d2c:	data_out=16'he;
17'h1d2d:	data_out=16'hb;
17'h1d2e:	data_out=16'hd;
17'h1d2f:	data_out=16'h8;
17'h1d30:	data_out=16'h17;
17'h1d31:	data_out=16'hc;
17'h1d32:	data_out=16'h1b;
17'h1d33:	data_out=16'hb;
17'h1d34:	data_out=16'h5;
17'h1d35:	data_out=16'h4;
17'h1d36:	data_out=16'h6;
17'h1d37:	data_out=16'h6;
17'h1d38:	data_out=16'h3;
17'h1d39:	data_out=16'h6;
17'h1d3a:	data_out=16'h8;
17'h1d3b:	data_out=16'h8001;
17'h1d3c:	data_out=16'h12;
17'h1d3d:	data_out=16'h3;
17'h1d3e:	data_out=16'h4;
17'h1d3f:	data_out=16'h8;
17'h1d40:	data_out=16'hd;
17'h1d41:	data_out=16'ha;
17'h1d42:	data_out=16'h5;
17'h1d43:	data_out=16'h8;
17'h1d44:	data_out=16'h0;
17'h1d45:	data_out=16'he;
17'h1d46:	data_out=16'h11;
17'h1d47:	data_out=16'h10;
17'h1d48:	data_out=16'h14;
17'h1d49:	data_out=16'he;
17'h1d4a:	data_out=16'h7;
17'h1d4b:	data_out=16'h5;
17'h1d4c:	data_out=16'h8;
17'h1d4d:	data_out=16'h16;
17'h1d4e:	data_out=16'ha;
17'h1d4f:	data_out=16'h1;
17'h1d50:	data_out=16'he;
17'h1d51:	data_out=16'ha;
17'h1d52:	data_out=16'h5;
17'h1d53:	data_out=16'hd;
17'h1d54:	data_out=16'h13;
17'h1d55:	data_out=16'h11;
17'h1d56:	data_out=16'ha;
17'h1d57:	data_out=16'h14;
17'h1d58:	data_out=16'h15;
17'h1d59:	data_out=16'hf;
17'h1d5a:	data_out=16'h5;
17'h1d5b:	data_out=16'he;
17'h1d5c:	data_out=16'h11;
17'h1d5d:	data_out=16'he;
17'h1d5e:	data_out=16'h17;
17'h1d5f:	data_out=16'h5;
17'h1d60:	data_out=16'hb;
17'h1d61:	data_out=16'ha;
17'h1d62:	data_out=16'h13;
17'h1d63:	data_out=16'h15;
17'h1d64:	data_out=16'h2;
17'h1d65:	data_out=16'h6;
17'h1d66:	data_out=16'h7;
17'h1d67:	data_out=16'h4;
17'h1d68:	data_out=16'h8001;
17'h1d69:	data_out=16'h4;
17'h1d6a:	data_out=16'h5;
17'h1d6b:	data_out=16'h10;
17'h1d6c:	data_out=16'h5;
17'h1d6d:	data_out=16'h9;
17'h1d6e:	data_out=16'h8003;
17'h1d6f:	data_out=16'h18;
17'h1d70:	data_out=16'h3;
17'h1d71:	data_out=16'hd;
17'h1d72:	data_out=16'h18;
17'h1d73:	data_out=16'h6;
17'h1d74:	data_out=16'hf;
17'h1d75:	data_out=16'h6;
17'h1d76:	data_out=16'he;
17'h1d77:	data_out=16'h1;
17'h1d78:	data_out=16'hc;
17'h1d79:	data_out=16'h6;
17'h1d7a:	data_out=16'h15;
17'h1d7b:	data_out=16'h7;
17'h1d7c:	data_out=16'h9;
17'h1d7d:	data_out=16'hb;
17'h1d7e:	data_out=16'hf;
17'h1d7f:	data_out=16'h4;
17'h1d80:	data_out=16'h39;
17'h1d81:	data_out=16'h2;
17'h1d82:	data_out=16'h8050;
17'h1d83:	data_out=16'h8077;
17'h1d84:	data_out=16'h8023;
17'h1d85:	data_out=16'h8075;
17'h1d86:	data_out=16'h8064;
17'h1d87:	data_out=16'h8006;
17'h1d88:	data_out=16'h1f;
17'h1d89:	data_out=16'hd;
17'h1d8a:	data_out=16'h4f;
17'h1d8b:	data_out=16'h8019;
17'h1d8c:	data_out=16'h62;
17'h1d8d:	data_out=16'h8085;
17'h1d8e:	data_out=16'h801b;
17'h1d8f:	data_out=16'h8088;
17'h1d90:	data_out=16'h8014;
17'h1d91:	data_out=16'h23;
17'h1d92:	data_out=16'h8040;
17'h1d93:	data_out=16'h8069;
17'h1d94:	data_out=16'h8092;
17'h1d95:	data_out=16'h803b;
17'h1d96:	data_out=16'h804c;
17'h1d97:	data_out=16'h8096;
17'h1d98:	data_out=16'h802e;
17'h1d99:	data_out=16'h45;
17'h1d9a:	data_out=16'h802c;
17'h1d9b:	data_out=16'h8084;
17'h1d9c:	data_out=16'h8090;
17'h1d9d:	data_out=16'h10;
17'h1d9e:	data_out=16'h808e;
17'h1d9f:	data_out=16'h8080;
17'h1da0:	data_out=16'h8063;
17'h1da1:	data_out=16'h8016;
17'h1da2:	data_out=16'h8024;
17'h1da3:	data_out=16'h41;
17'h1da4:	data_out=16'h3c;
17'h1da5:	data_out=16'h800c;
17'h1da6:	data_out=16'h19;
17'h1da7:	data_out=16'h4;
17'h1da8:	data_out=16'h801f;
17'h1da9:	data_out=16'h8073;
17'h1daa:	data_out=16'h802b;
17'h1dab:	data_out=16'h17;
17'h1dac:	data_out=16'h803c;
17'h1dad:	data_out=16'h23;
17'h1dae:	data_out=16'h8076;
17'h1daf:	data_out=16'h8065;
17'h1db0:	data_out=16'h8018;
17'h1db1:	data_out=16'h5d;
17'h1db2:	data_out=16'h8017;
17'h1db3:	data_out=16'h809e;
17'h1db4:	data_out=16'h47;
17'h1db5:	data_out=16'h23;
17'h1db6:	data_out=16'h8034;
17'h1db7:	data_out=16'h8067;
17'h1db8:	data_out=16'h805b;
17'h1db9:	data_out=16'h8084;
17'h1dba:	data_out=16'h8020;
17'h1dbb:	data_out=16'h59;
17'h1dbc:	data_out=16'h8041;
17'h1dbd:	data_out=16'h8044;
17'h1dbe:	data_out=16'h8019;
17'h1dbf:	data_out=16'h806d;
17'h1dc0:	data_out=16'h8062;
17'h1dc1:	data_out=16'h805c;
17'h1dc2:	data_out=16'h2a;
17'h1dc3:	data_out=16'h8083;
17'h1dc4:	data_out=16'h8007;
17'h1dc5:	data_out=16'h803b;
17'h1dc6:	data_out=16'h8032;
17'h1dc7:	data_out=16'h8016;
17'h1dc8:	data_out=16'h804e;
17'h1dc9:	data_out=16'h8023;
17'h1dca:	data_out=16'h8016;
17'h1dcb:	data_out=16'h2a;
17'h1dcc:	data_out=16'h8015;
17'h1dcd:	data_out=16'h803e;
17'h1dce:	data_out=16'h8031;
17'h1dcf:	data_out=16'h8016;
17'h1dd0:	data_out=16'h807c;
17'h1dd1:	data_out=16'h8078;
17'h1dd2:	data_out=16'h22;
17'h1dd3:	data_out=16'h804e;
17'h1dd4:	data_out=16'h8061;
17'h1dd5:	data_out=16'h8063;
17'h1dd6:	data_out=16'h805b;
17'h1dd7:	data_out=16'h804a;
17'h1dd8:	data_out=16'h8048;
17'h1dd9:	data_out=16'h8048;
17'h1dda:	data_out=16'h8064;
17'h1ddb:	data_out=16'h8054;
17'h1ddc:	data_out=16'h802c;
17'h1ddd:	data_out=16'h804e;
17'h1dde:	data_out=16'h806b;
17'h1ddf:	data_out=16'h8030;
17'h1de0:	data_out=16'h8003;
17'h1de1:	data_out=16'h804a;
17'h1de2:	data_out=16'h808e;
17'h1de3:	data_out=16'h8091;
17'h1de4:	data_out=16'h33;
17'h1de5:	data_out=16'h19;
17'h1de6:	data_out=16'h2f;
17'h1de7:	data_out=16'h8040;
17'h1de8:	data_out=16'h8026;
17'h1de9:	data_out=16'h1;
17'h1dea:	data_out=16'h801a;
17'h1deb:	data_out=16'h803f;
17'h1dec:	data_out=16'h2c;
17'h1ded:	data_out=16'h8093;
17'h1dee:	data_out=16'h8021;
17'h1def:	data_out=16'h8066;
17'h1df0:	data_out=16'h8021;
17'h1df1:	data_out=16'h8058;
17'h1df2:	data_out=16'h8070;
17'h1df3:	data_out=16'h806d;
17'h1df4:	data_out=16'h801d;
17'h1df5:	data_out=16'h8076;
17'h1df6:	data_out=16'h37;
17'h1df7:	data_out=16'h8060;
17'h1df8:	data_out=16'h8055;
17'h1df9:	data_out=16'h8072;
17'h1dfa:	data_out=16'h8091;
17'h1dfb:	data_out=16'h8022;
17'h1dfc:	data_out=16'h802b;
17'h1dfd:	data_out=16'h808e;
17'h1dfe:	data_out=16'h9;
17'h1dff:	data_out=16'h8066;
17'h1e00:	data_out=16'h39;
17'h1e01:	data_out=16'h77;
17'h1e02:	data_out=16'h4c;
17'h1e03:	data_out=16'h32;
17'h1e04:	data_out=16'h66;
17'h1e05:	data_out=16'h62;
17'h1e06:	data_out=16'h1d;
17'h1e07:	data_out=16'h28;
17'h1e08:	data_out=16'h45;
17'h1e09:	data_out=16'h3;
17'h1e0a:	data_out=16'h9d;
17'h1e0b:	data_out=16'h89;
17'h1e0c:	data_out=16'h8d;
17'h1e0d:	data_out=16'h16;
17'h1e0e:	data_out=16'h14;
17'h1e0f:	data_out=16'h11;
17'h1e10:	data_out=16'h2b;
17'h1e11:	data_out=16'h78;
17'h1e12:	data_out=16'h19;
17'h1e13:	data_out=16'h45;
17'h1e14:	data_out=16'h40;
17'h1e15:	data_out=16'he;
17'h1e16:	data_out=16'h2c;
17'h1e17:	data_out=16'h52;
17'h1e18:	data_out=16'h3;
17'h1e19:	data_out=16'h3c;
17'h1e1a:	data_out=16'h5b;
17'h1e1b:	data_out=16'h4a;
17'h1e1c:	data_out=16'h4c;
17'h1e1d:	data_out=16'h9e;
17'h1e1e:	data_out=16'h20;
17'h1e1f:	data_out=16'h800b;
17'h1e20:	data_out=16'h57;
17'h1e21:	data_out=16'h12;
17'h1e22:	data_out=16'h34;
17'h1e23:	data_out=16'h30;
17'h1e24:	data_out=16'h2d;
17'h1e25:	data_out=16'h38;
17'h1e26:	data_out=16'h2d;
17'h1e27:	data_out=16'h85;
17'h1e28:	data_out=16'hc;
17'h1e29:	data_out=16'h18;
17'h1e2a:	data_out=16'h35;
17'h1e2b:	data_out=16'h49;
17'h1e2c:	data_out=16'h5e;
17'h1e2d:	data_out=16'ha9;
17'h1e2e:	data_out=16'h2c;
17'h1e2f:	data_out=16'h5f;
17'h1e30:	data_out=16'hb6;
17'h1e31:	data_out=16'h71;
17'h1e32:	data_out=16'hb6;
17'h1e33:	data_out=16'h2a;
17'h1e34:	data_out=16'h6b;
17'h1e35:	data_out=16'hb0;
17'h1e36:	data_out=16'h60;
17'h1e37:	data_out=16'h49;
17'h1e38:	data_out=16'h1e;
17'h1e39:	data_out=16'h8;
17'h1e3a:	data_out=16'h13;
17'h1e3b:	data_out=16'h6b;
17'h1e3c:	data_out=16'h92;
17'h1e3d:	data_out=16'h2f;
17'h1e3e:	data_out=16'hc;
17'h1e3f:	data_out=16'h72;
17'h1e40:	data_out=16'h31;
17'h1e41:	data_out=16'h5e;
17'h1e42:	data_out=16'h84;
17'h1e43:	data_out=16'h24;
17'h1e44:	data_out=16'h78;
17'h1e45:	data_out=16'hb;
17'h1e46:	data_out=16'h78;
17'h1e47:	data_out=16'hf;
17'h1e48:	data_out=16'hb;
17'h1e49:	data_out=16'h39;
17'h1e4a:	data_out=16'h3f;
17'h1e4b:	data_out=16'h8e;
17'h1e4c:	data_out=16'h31;
17'h1e4d:	data_out=16'h22;
17'h1e4e:	data_out=16'h4c;
17'h1e4f:	data_out=16'h39;
17'h1e50:	data_out=16'he;
17'h1e51:	data_out=16'h17;
17'h1e52:	data_out=16'h2d;
17'h1e53:	data_out=16'h86;
17'h1e54:	data_out=16'h69;
17'h1e55:	data_out=16'h50;
17'h1e56:	data_out=16'h43;
17'h1e57:	data_out=16'h1f;
17'h1e58:	data_out=16'h5b;
17'h1e59:	data_out=16'h54;
17'h1e5a:	data_out=16'h44;
17'h1e5b:	data_out=16'h62;
17'h1e5c:	data_out=16'h63;
17'h1e5d:	data_out=16'h4b;
17'h1e5e:	data_out=16'h75;
17'h1e5f:	data_out=16'h17;
17'h1e60:	data_out=16'h55;
17'h1e61:	data_out=16'h70;
17'h1e62:	data_out=16'h4a;
17'h1e63:	data_out=16'h3b;
17'h1e64:	data_out=16'h64;
17'h1e65:	data_out=16'h6b;
17'h1e66:	data_out=16'h3a;
17'h1e67:	data_out=16'h15;
17'h1e68:	data_out=16'h12;
17'h1e69:	data_out=16'h5e;
17'h1e6a:	data_out=16'hf;
17'h1e6b:	data_out=16'h2d;
17'h1e6c:	data_out=16'h93;
17'h1e6d:	data_out=16'h26;
17'h1e6e:	data_out=16'h16;
17'h1e6f:	data_out=16'h5a;
17'h1e70:	data_out=16'h13;
17'h1e71:	data_out=16'h8008;
17'h1e72:	data_out=16'h60;
17'h1e73:	data_out=16'h45;
17'h1e74:	data_out=16'hc7;
17'h1e75:	data_out=16'h8b;
17'h1e76:	data_out=16'h30;
17'h1e77:	data_out=16'h4f;
17'h1e78:	data_out=16'h13;
17'h1e79:	data_out=16'h39;
17'h1e7a:	data_out=16'h37;
17'h1e7b:	data_out=16'hb;
17'h1e7c:	data_out=16'h8;
17'h1e7d:	data_out=16'he;
17'h1e7e:	data_out=16'h14;
17'h1e7f:	data_out=16'h1f;
17'h1e80:	data_out=16'h8011;
17'h1e81:	data_out=16'ha;
17'h1e82:	data_out=16'h12;
17'h1e83:	data_out=16'h32;
17'h1e84:	data_out=16'h4d;
17'h1e85:	data_out=16'h45;
17'h1e86:	data_out=16'h1a;
17'h1e87:	data_out=16'h1f;
17'h1e88:	data_out=16'h800f;
17'h1e89:	data_out=16'h6;
17'h1e8a:	data_out=16'h1d;
17'h1e8b:	data_out=16'h3d;
17'h1e8c:	data_out=16'h44;
17'h1e8d:	data_out=16'h2a;
17'h1e8e:	data_out=16'hb;
17'h1e8f:	data_out=16'h8008;
17'h1e90:	data_out=16'hf;
17'h1e91:	data_out=16'h37;
17'h1e92:	data_out=16'h6;
17'h1e93:	data_out=16'h37;
17'h1e94:	data_out=16'h14;
17'h1e95:	data_out=16'h11;
17'h1e96:	data_out=16'h1e;
17'h1e97:	data_out=16'h24;
17'h1e98:	data_out=16'h6;
17'h1e99:	data_out=16'h2b;
17'h1e9a:	data_out=16'h63;
17'h1e9b:	data_out=16'h24;
17'h1e9c:	data_out=16'h27;
17'h1e9d:	data_out=16'h16;
17'h1e9e:	data_out=16'h6;
17'h1e9f:	data_out=16'h1f;
17'h1ea0:	data_out=16'h25;
17'h1ea1:	data_out=16'h15;
17'h1ea2:	data_out=16'h38;
17'h1ea3:	data_out=16'h8006;
17'h1ea4:	data_out=16'h8008;
17'h1ea5:	data_out=16'h20;
17'h1ea6:	data_out=16'h800f;
17'h1ea7:	data_out=16'h1d;
17'h1ea8:	data_out=16'h15;
17'h1ea9:	data_out=16'h18;
17'h1eaa:	data_out=16'h8004;
17'h1eab:	data_out=16'h14;
17'h1eac:	data_out=16'h2a;
17'h1ead:	data_out=16'h48;
17'h1eae:	data_out=16'h17;
17'h1eaf:	data_out=16'h39;
17'h1eb0:	data_out=16'ha5;
17'h1eb1:	data_out=16'ha;
17'h1eb2:	data_out=16'h9d;
17'h1eb3:	data_out=16'h16;
17'h1eb4:	data_out=16'h3;
17'h1eb5:	data_out=16'h57;
17'h1eb6:	data_out=16'h15;
17'h1eb7:	data_out=16'h21;
17'h1eb8:	data_out=16'h800c;
17'h1eb9:	data_out=16'h800f;
17'h1eba:	data_out=16'h12;
17'h1ebb:	data_out=16'h28;
17'h1ebc:	data_out=16'h1e;
17'h1ebd:	data_out=16'h8;
17'h1ebe:	data_out=16'he;
17'h1ebf:	data_out=16'h5e;
17'h1ec0:	data_out=16'h47;
17'h1ec1:	data_out=16'h27;
17'h1ec2:	data_out=16'h45;
17'h1ec3:	data_out=16'h33;
17'h1ec4:	data_out=16'h32;
17'h1ec5:	data_out=16'h1;
17'h1ec6:	data_out=16'h21;
17'h1ec7:	data_out=16'h18;
17'h1ec8:	data_out=16'h1b;
17'h1ec9:	data_out=16'h1d;
17'h1eca:	data_out=16'h3b;
17'h1ecb:	data_out=16'h4c;
17'h1ecc:	data_out=16'h33;
17'h1ecd:	data_out=16'h25;
17'h1ece:	data_out=16'h2d;
17'h1ecf:	data_out=16'h2b;
17'h1ed0:	data_out=16'h33;
17'h1ed1:	data_out=16'h8000;
17'h1ed2:	data_out=16'h8002;
17'h1ed3:	data_out=16'h31;
17'h1ed4:	data_out=16'h30;
17'h1ed5:	data_out=16'h16;
17'h1ed6:	data_out=16'h21;
17'h1ed7:	data_out=16'h12;
17'h1ed8:	data_out=16'h7;
17'h1ed9:	data_out=16'h38;
17'h1eda:	data_out=16'h8;
17'h1edb:	data_out=16'h15;
17'h1edc:	data_out=16'h16;
17'h1edd:	data_out=16'h30;
17'h1ede:	data_out=16'h4d;
17'h1edf:	data_out=16'h12;
17'h1ee0:	data_out=16'h8;
17'h1ee1:	data_out=16'h3f;
17'h1ee2:	data_out=16'h6;
17'h1ee3:	data_out=16'h17;
17'h1ee4:	data_out=16'h8008;
17'h1ee5:	data_out=16'h42;
17'h1ee6:	data_out=16'h20;
17'h1ee7:	data_out=16'h14;
17'h1ee8:	data_out=16'hd;
17'h1ee9:	data_out=16'hd;
17'h1eea:	data_out=16'h7;
17'h1eeb:	data_out=16'h3f;
17'h1eec:	data_out=16'h17;
17'h1eed:	data_out=16'h8;
17'h1eee:	data_out=16'hf;
17'h1eef:	data_out=16'h74;
17'h1ef0:	data_out=16'h7;
17'h1ef1:	data_out=16'h8011;
17'h1ef2:	data_out=16'h51;
17'h1ef3:	data_out=16'h37;
17'h1ef4:	data_out=16'h9a;
17'h1ef5:	data_out=16'h34;
17'h1ef6:	data_out=16'h6;
17'h1ef7:	data_out=16'h47;
17'h1ef8:	data_out=16'h18;
17'h1ef9:	data_out=16'h12;
17'h1efa:	data_out=16'h1c;
17'h1efb:	data_out=16'h10;
17'h1efc:	data_out=16'h8001;
17'h1efd:	data_out=16'h18;
17'h1efe:	data_out=16'ha;
17'h1eff:	data_out=16'h2b;
17'h1f00:	data_out=16'h82e3;
17'h1f01:	data_out=16'h82d7;
17'h1f02:	data_out=16'h81fe;
17'h1f03:	data_out=16'h8071;
17'h1f04:	data_out=16'h36b;
17'h1f05:	data_out=16'h195;
17'h1f06:	data_out=16'h8035;
17'h1f07:	data_out=16'h8041;
17'h1f08:	data_out=16'h8293;
17'h1f09:	data_out=16'h80b5;
17'h1f0a:	data_out=16'h81d5;
17'h1f0b:	data_out=16'h7a;
17'h1f0c:	data_out=16'h32a;
17'h1f0d:	data_out=16'h805f;
17'h1f0e:	data_out=16'h8021;
17'h1f0f:	data_out=16'h823e;
17'h1f10:	data_out=16'h8062;
17'h1f11:	data_out=16'h149;
17'h1f12:	data_out=16'h8137;
17'h1f13:	data_out=16'h35;
17'h1f14:	data_out=16'h82b7;
17'h1f15:	data_out=16'h8154;
17'h1f16:	data_out=16'h80f7;
17'h1f17:	data_out=16'h823e;
17'h1f18:	data_out=16'h80d3;
17'h1f19:	data_out=16'h182;
17'h1f1a:	data_out=16'h434;
17'h1f1b:	data_out=16'h8165;
17'h1f1c:	data_out=16'h8249;
17'h1f1d:	data_out=16'h828e;
17'h1f1e:	data_out=16'h8329;
17'h1f1f:	data_out=16'h80f7;
17'h1f20:	data_out=16'h8190;
17'h1f21:	data_out=16'h8022;
17'h1f22:	data_out=16'h18;
17'h1f23:	data_out=16'h8172;
17'h1f24:	data_out=16'h8172;
17'h1f25:	data_out=16'h154;
17'h1f26:	data_out=16'h8279;
17'h1f27:	data_out=16'h82c7;
17'h1f28:	data_out=16'h801d;
17'h1f29:	data_out=16'h8145;
17'h1f2a:	data_out=16'h81e3;
17'h1f2b:	data_out=16'h8141;
17'h1f2c:	data_out=16'h8028;
17'h1f2d:	data_out=16'h1bb;
17'h1f2e:	data_out=16'h80e4;
17'h1f2f:	data_out=16'h80ab;
17'h1f30:	data_out=16'h4ca;
17'h1f31:	data_out=16'h826b;
17'h1f32:	data_out=16'h4bc;
17'h1f33:	data_out=16'h8311;
17'h1f34:	data_out=16'h81f6;
17'h1f35:	data_out=16'h27b;
17'h1f36:	data_out=16'h81f6;
17'h1f37:	data_out=16'h81b9;
17'h1f38:	data_out=16'h8345;
17'h1f39:	data_out=16'h8390;
17'h1f3a:	data_out=16'h8101;
17'h1f3b:	data_out=16'hb7;
17'h1f3c:	data_out=16'h820d;
17'h1f3d:	data_out=16'h8172;
17'h1f3e:	data_out=16'h8015;
17'h1f3f:	data_out=16'h28e;
17'h1f40:	data_out=16'h2e3;
17'h1f41:	data_out=16'h80ff;
17'h1f42:	data_out=16'h31d;
17'h1f43:	data_out=16'hdc;
17'h1f44:	data_out=16'h2c;
17'h1f45:	data_out=16'h8152;
17'h1f46:	data_out=16'h819f;
17'h1f47:	data_out=16'h8057;
17'h1f48:	data_out=16'h23;
17'h1f49:	data_out=16'h125;
17'h1f4a:	data_out=16'h1d6;
17'h1f4b:	data_out=16'h26c;
17'h1f4c:	data_out=16'h1d8;
17'h1f4d:	data_out=16'h8072;
17'h1f4e:	data_out=16'hd;
17'h1f4f:	data_out=16'h1a3;
17'h1f50:	data_out=16'h17c;
17'h1f51:	data_out=16'h8227;
17'h1f52:	data_out=16'h815d;
17'h1f53:	data_out=16'h8208;
17'h1f54:	data_out=16'h8152;
17'h1f55:	data_out=16'h82ab;
17'h1f56:	data_out=16'h814b;
17'h1f57:	data_out=16'h81a3;
17'h1f58:	data_out=16'h8271;
17'h1f59:	data_out=16'h13b;
17'h1f5a:	data_out=16'h8282;
17'h1f5b:	data_out=16'h82db;
17'h1f5c:	data_out=16'h80f5;
17'h1f5d:	data_out=16'h800f;
17'h1f5e:	data_out=16'h108;
17'h1f5f:	data_out=16'h80d6;
17'h1f60:	data_out=16'h8162;
17'h1f61:	data_out=16'h804c;
17'h1f62:	data_out=16'h82b6;
17'h1f63:	data_out=16'h82b3;
17'h1f64:	data_out=16'h8251;
17'h1f65:	data_out=16'h2e5;
17'h1f66:	data_out=16'h1c3;
17'h1f67:	data_out=16'h807b;
17'h1f68:	data_out=16'h8024;
17'h1f69:	data_out=16'h81f2;
17'h1f6a:	data_out=16'h802f;
17'h1f6b:	data_out=16'h228;
17'h1f6c:	data_out=16'h8228;
17'h1f6d:	data_out=16'h830c;
17'h1f6e:	data_out=16'h802f;
17'h1f6f:	data_out=16'h3ad;
17'h1f70:	data_out=16'h8024;
17'h1f71:	data_out=16'h8255;
17'h1f72:	data_out=16'h1ad;
17'h1f73:	data_out=16'hab;
17'h1f74:	data_out=16'h4d6;
17'h1f75:	data_out=16'h8046;
17'h1f76:	data_out=16'h81a6;
17'h1f77:	data_out=16'h28e;
17'h1f78:	data_out=16'h95;
17'h1f79:	data_out=16'h81ca;
17'h1f7a:	data_out=16'h82ba;
17'h1f7b:	data_out=16'h8015;
17'h1f7c:	data_out=16'h819c;
17'h1f7d:	data_out=16'h80a9;
17'h1f7e:	data_out=16'h8088;
17'h1f7f:	data_out=16'h19c;
17'h1f80:	data_out=16'h83a0;
17'h1f81:	data_out=16'h8289;
17'h1f82:	data_out=16'h8289;
17'h1f83:	data_out=16'h171;
17'h1f84:	data_out=16'h889;
17'h1f85:	data_out=16'h5b9;
17'h1f86:	data_out=16'hc7;
17'h1f87:	data_out=16'hc7;
17'h1f88:	data_out=16'h8284;
17'h1f89:	data_out=16'h814e;
17'h1f8a:	data_out=16'h8118;
17'h1f8b:	data_out=16'h98;
17'h1f8c:	data_out=16'h7c6;
17'h1f8d:	data_out=16'h81a6;
17'h1f8e:	data_out=16'h8077;
17'h1f8f:	data_out=16'h8396;
17'h1f90:	data_out=16'h127;
17'h1f91:	data_out=16'h4cb;
17'h1f92:	data_out=16'h8234;
17'h1f93:	data_out=16'had;
17'h1f94:	data_out=16'h8690;
17'h1f95:	data_out=16'h8148;
17'h1f96:	data_out=16'h19;
17'h1f97:	data_out=16'h84fe;
17'h1f98:	data_out=16'h82f8;
17'h1f99:	data_out=16'h386;
17'h1f9a:	data_out=16'h978;
17'h1f9b:	data_out=16'h8274;
17'h1f9c:	data_out=16'h8268;
17'h1f9d:	data_out=16'h8289;
17'h1f9e:	data_out=16'h85fd;
17'h1f9f:	data_out=16'h82ec;
17'h1fa0:	data_out=16'h8310;
17'h1fa1:	data_out=16'h8064;
17'h1fa2:	data_out=16'h8078;
17'h1fa3:	data_out=16'h81cf;
17'h1fa4:	data_out=16'h81cf;
17'h1fa5:	data_out=16'h2b6;
17'h1fa6:	data_out=16'h83af;
17'h1fa7:	data_out=16'h832d;
17'h1fa8:	data_out=16'h8041;
17'h1fa9:	data_out=16'h82f1;
17'h1faa:	data_out=16'h830b;
17'h1fab:	data_out=16'h822a;
17'h1fac:	data_out=16'he9;
17'h1fad:	data_out=16'h4bc;
17'h1fae:	data_out=16'h81d4;
17'h1faf:	data_out=16'h189;
17'h1fb0:	data_out=16'ha00;
17'h1fb1:	data_out=16'h82e6;
17'h1fb2:	data_out=16'ha00;
17'h1fb3:	data_out=16'h8762;
17'h1fb4:	data_out=16'h82d3;
17'h1fb5:	data_out=16'h65d;
17'h1fb6:	data_out=16'h8210;
17'h1fb7:	data_out=16'h8290;
17'h1fb8:	data_out=16'h84e5;
17'h1fb9:	data_out=16'h876d;
17'h1fba:	data_out=16'h813f;
17'h1fbb:	data_out=16'h550;
17'h1fbc:	data_out=16'h8071;
17'h1fbd:	data_out=16'h8268;
17'h1fbe:	data_out=16'h8042;
17'h1fbf:	data_out=16'h629;
17'h1fc0:	data_out=16'h72e;
17'h1fc1:	data_out=16'h8063;
17'h1fc2:	data_out=16'h850;
17'h1fc3:	data_out=16'h8016;
17'h1fc4:	data_out=16'hd0;
17'h1fc5:	data_out=16'h813b;
17'h1fc6:	data_out=16'h80dc;
17'h1fc7:	data_out=16'h80af;
17'h1fc8:	data_out=16'h8051;
17'h1fc9:	data_out=16'h2f2;
17'h1fca:	data_out=16'h336;
17'h1fcb:	data_out=16'h519;
17'h1fcc:	data_out=16'h2dd;
17'h1fcd:	data_out=16'h807b;
17'h1fce:	data_out=16'h7d;
17'h1fcf:	data_out=16'h25c;
17'h1fd0:	data_out=16'h311;
17'h1fd1:	data_out=16'h827f;
17'h1fd2:	data_out=16'h817f;
17'h1fd3:	data_out=16'h825b;
17'h1fd4:	data_out=16'h819f;
17'h1fd5:	data_out=16'h8398;
17'h1fd6:	data_out=16'h833d;
17'h1fd7:	data_out=16'h833c;
17'h1fd8:	data_out=16'h8295;
17'h1fd9:	data_out=16'h481;
17'h1fda:	data_out=16'h83ad;
17'h1fdb:	data_out=16'h8326;
17'h1fdc:	data_out=16'h68;
17'h1fdd:	data_out=16'h163;
17'h1fde:	data_out=16'h251;
17'h1fdf:	data_out=16'h8214;
17'h1fe0:	data_out=16'h81f5;
17'h1fe1:	data_out=16'h8058;
17'h1fe2:	data_out=16'h84f9;
17'h1fe3:	data_out=16'h86a0;
17'h1fe4:	data_out=16'h8434;
17'h1fe5:	data_out=16'h71d;
17'h1fe6:	data_out=16'h2fb;
17'h1fe7:	data_out=16'h8169;
17'h1fe8:	data_out=16'h8062;
17'h1fe9:	data_out=16'h8252;
17'h1fea:	data_out=16'h8088;
17'h1feb:	data_out=16'h5d7;
17'h1fec:	data_out=16'h8111;
17'h1fed:	data_out=16'h871f;
17'h1fee:	data_out=16'h8082;
17'h1fef:	data_out=16'ha00;
17'h1ff0:	data_out=16'h8070;
17'h1ff1:	data_out=16'h86bd;
17'h1ff2:	data_out=16'h507;
17'h1ff3:	data_out=16'h3f3;
17'h1ff4:	data_out=16'ha00;
17'h1ff5:	data_out=16'hab;
17'h1ff6:	data_out=16'h828b;
17'h1ff7:	data_out=16'h480;
17'h1ff8:	data_out=16'h140;
17'h1ff9:	data_out=16'h8337;
17'h1ffa:	data_out=16'h86a5;
17'h1ffb:	data_out=16'h803f;
17'h1ffc:	data_out=16'h82b9;
17'h1ffd:	data_out=16'h8131;
17'h1ffe:	data_out=16'h802e;
17'h1fff:	data_out=16'h313;
17'h2000:	data_out=16'h8688;
17'h2001:	data_out=16'h83de;
17'h2002:	data_out=16'h81aa;
17'h2003:	data_out=16'h56a;
17'h2004:	data_out=16'ha00;
17'h2005:	data_out=16'ha00;
17'h2006:	data_out=16'h3a5;
17'h2007:	data_out=16'h28b;
17'h2008:	data_out=16'h82cf;
17'h2009:	data_out=16'h800d;
17'h200a:	data_out=16'h830e;
17'h200b:	data_out=16'hdf;
17'h200c:	data_out=16'ha00;
17'h200d:	data_out=16'h8082;
17'h200e:	data_out=16'he0;
17'h200f:	data_out=16'h82c9;
17'h2010:	data_out=16'h46d;
17'h2011:	data_out=16'h783;
17'h2012:	data_out=16'h8102;
17'h2013:	data_out=16'h408;
17'h2014:	data_out=16'h85fd;
17'h2015:	data_out=16'h80f9;
17'h2016:	data_out=16'h190;
17'h2017:	data_out=16'h838d;
17'h2018:	data_out=16'h83af;
17'h2019:	data_out=16'h439;
17'h201a:	data_out=16'ha00;
17'h201b:	data_out=16'h8121;
17'h201c:	data_out=16'h81ab;
17'h201d:	data_out=16'h8365;
17'h201e:	data_out=16'h8680;
17'h201f:	data_out=16'h80da;
17'h2020:	data_out=16'h821f;
17'h2021:	data_out=16'hed;
17'h2022:	data_out=16'h2f5;
17'h2023:	data_out=16'h8240;
17'h2024:	data_out=16'h8240;
17'h2025:	data_out=16'h58f;
17'h2026:	data_out=16'h8488;
17'h2027:	data_out=16'h843d;
17'h2028:	data_out=16'h127;
17'h2029:	data_out=16'h83ff;
17'h202a:	data_out=16'h8188;
17'h202b:	data_out=16'h81f2;
17'h202c:	data_out=16'h20d;
17'h202d:	data_out=16'h665;
17'h202e:	data_out=16'ha7;
17'h202f:	data_out=16'h4bf;
17'h2030:	data_out=16'ha00;
17'h2031:	data_out=16'h860c;
17'h2032:	data_out=16'ha00;
17'h2033:	data_out=16'h87ca;
17'h2034:	data_out=16'h866b;
17'h2035:	data_out=16'h9d2;
17'h2036:	data_out=16'h823e;
17'h2037:	data_out=16'h81a8;
17'h2038:	data_out=16'h84b5;
17'h2039:	data_out=16'h88d4;
17'h203a:	data_out=16'h52;
17'h203b:	data_out=16'h6d3;
17'h203c:	data_out=16'h123;
17'h203d:	data_out=16'h8250;
17'h203e:	data_out=16'h12b;
17'h203f:	data_out=16'ha00;
17'h2040:	data_out=16'ha00;
17'h2041:	data_out=16'he8;
17'h2042:	data_out=16'ha00;
17'h2043:	data_out=16'h32b;
17'h2044:	data_out=16'h1f;
17'h2045:	data_out=16'h80dd;
17'h2046:	data_out=16'h3f;
17'h2047:	data_out=16'h82;
17'h2048:	data_out=16'h32a;
17'h2049:	data_out=16'h5ce;
17'h204a:	data_out=16'h5ff;
17'h204b:	data_out=16'h87d;
17'h204c:	data_out=16'h533;
17'h204d:	data_out=16'h26e;
17'h204e:	data_out=16'h32a;
17'h204f:	data_out=16'h449;
17'h2050:	data_out=16'h853;
17'h2051:	data_out=16'h80c4;
17'h2052:	data_out=16'h81ba;
17'h2053:	data_out=16'h810d;
17'h2054:	data_out=16'h8083;
17'h2055:	data_out=16'h833c;
17'h2056:	data_out=16'h8159;
17'h2057:	data_out=16'h81e3;
17'h2058:	data_out=16'h8243;
17'h2059:	data_out=16'h96b;
17'h205a:	data_out=16'h82ef;
17'h205b:	data_out=16'h83cd;
17'h205c:	data_out=16'h139;
17'h205d:	data_out=16'h440;
17'h205e:	data_out=16'h66e;
17'h205f:	data_out=16'h81dd;
17'h2060:	data_out=16'h845e;
17'h2061:	data_out=16'ha7;
17'h2062:	data_out=16'h8553;
17'h2063:	data_out=16'h86d3;
17'h2064:	data_out=16'h8842;
17'h2065:	data_out=16'h9dd;
17'h2066:	data_out=16'h3cb;
17'h2067:	data_out=16'h162;
17'h2068:	data_out=16'h105;
17'h2069:	data_out=16'h82e7;
17'h206a:	data_out=16'hb3;
17'h206b:	data_out=16'ha00;
17'h206c:	data_out=16'h821c;
17'h206d:	data_out=16'h8789;
17'h206e:	data_out=16'hc3;
17'h206f:	data_out=16'ha00;
17'h2070:	data_out=16'hcd;
17'h2071:	data_out=16'h875c;
17'h2072:	data_out=16'h8e8;
17'h2073:	data_out=16'h86d;
17'h2074:	data_out=16'ha00;
17'h2075:	data_out=16'h204;
17'h2076:	data_out=16'h8298;
17'h2077:	data_out=16'h9f1;
17'h2078:	data_out=16'h592;
17'h2079:	data_out=16'h80f1;
17'h207a:	data_out=16'h8621;
17'h207b:	data_out=16'h126;
17'h207c:	data_out=16'h8353;
17'h207d:	data_out=16'h10f;
17'h207e:	data_out=16'h1a9;
17'h207f:	data_out=16'h6bb;
17'h2080:	data_out=16'h85e0;
17'h2081:	data_out=16'h8110;
17'h2082:	data_out=16'h8135;
17'h2083:	data_out=16'h9ff;
17'h2084:	data_out=16'ha00;
17'h2085:	data_out=16'ha00;
17'h2086:	data_out=16'h873;
17'h2087:	data_out=16'h573;
17'h2088:	data_out=16'h842d;
17'h2089:	data_out=16'h373;
17'h208a:	data_out=16'h8162;
17'h208b:	data_out=16'h31;
17'h208c:	data_out=16'ha00;
17'h208d:	data_out=16'h21c;
17'h208e:	data_out=16'h25d;
17'h208f:	data_out=16'h82f1;
17'h2090:	data_out=16'h904;
17'h2091:	data_out=16'h91d;
17'h2092:	data_out=16'h8107;
17'h2093:	data_out=16'h9f5;
17'h2094:	data_out=16'h84b0;
17'h2095:	data_out=16'hf1;
17'h2096:	data_out=16'h4a7;
17'h2097:	data_out=16'h81af;
17'h2098:	data_out=16'h84a8;
17'h2099:	data_out=16'h710;
17'h209a:	data_out=16'ha00;
17'h209b:	data_out=16'h35e;
17'h209c:	data_out=16'h6a9;
17'h209d:	data_out=16'h80a5;
17'h209e:	data_out=16'h84de;
17'h209f:	data_out=16'h351;
17'h20a0:	data_out=16'h561;
17'h20a1:	data_out=16'h263;
17'h20a2:	data_out=16'h981;
17'h20a3:	data_out=16'h831a;
17'h20a4:	data_out=16'h8319;
17'h20a5:	data_out=16'ha00;
17'h20a6:	data_out=16'h855b;
17'h20a7:	data_out=16'h8114;
17'h20a8:	data_out=16'h264;
17'h20a9:	data_out=16'h83ca;
17'h20aa:	data_out=16'h83a1;
17'h20ab:	data_out=16'h162;
17'h20ac:	data_out=16'h53a;
17'h20ad:	data_out=16'h9eb;
17'h20ae:	data_out=16'h10b;
17'h20af:	data_out=16'ha00;
17'h20b0:	data_out=16'ha00;
17'h20b1:	data_out=16'h83d5;
17'h20b2:	data_out=16'ha00;
17'h20b3:	data_out=16'h8631;
17'h20b4:	data_out=16'h8586;
17'h20b5:	data_out=16'h9f6;
17'h20b6:	data_out=16'h834f;
17'h20b7:	data_out=16'h8112;
17'h20b8:	data_out=16'h59a;
17'h20b9:	data_out=16'h87c0;
17'h20ba:	data_out=16'h2aa;
17'h20bb:	data_out=16'ha00;
17'h20bc:	data_out=16'h4e9;
17'h20bd:	data_out=16'h667;
17'h20be:	data_out=16'h263;
17'h20bf:	data_out=16'ha00;
17'h20c0:	data_out=16'ha00;
17'h20c1:	data_out=16'h244;
17'h20c2:	data_out=16'ha00;
17'h20c3:	data_out=16'h858;
17'h20c4:	data_out=16'h25e;
17'h20c5:	data_out=16'h125;
17'h20c6:	data_out=16'h22e;
17'h20c7:	data_out=16'h22f;
17'h20c8:	data_out=16'h491;
17'h20c9:	data_out=16'ha00;
17'h20ca:	data_out=16'ha00;
17'h20cb:	data_out=16'ha00;
17'h20cc:	data_out=16'h96e;
17'h20cd:	data_out=16'h9ce;
17'h20ce:	data_out=16'h40b;
17'h20cf:	data_out=16'h7c0;
17'h20d0:	data_out=16'ha00;
17'h20d1:	data_out=16'h300;
17'h20d2:	data_out=16'h823b;
17'h20d3:	data_out=16'h529;
17'h20d4:	data_out=16'h7ac;
17'h20d5:	data_out=16'h831c;
17'h20d6:	data_out=16'h15f;
17'h20d7:	data_out=16'h1e2;
17'h20d8:	data_out=16'h82ba;
17'h20d9:	data_out=16'ha00;
17'h20da:	data_out=16'h99;
17'h20db:	data_out=16'h9c;
17'h20dc:	data_out=16'h4c9;
17'h20dd:	data_out=16'h9a4;
17'h20de:	data_out=16'ha00;
17'h20df:	data_out=16'h81c5;
17'h20e0:	data_out=16'h8867;
17'h20e1:	data_out=16'h6c4;
17'h20e2:	data_out=16'h85e1;
17'h20e3:	data_out=16'h8571;
17'h20e4:	data_out=16'h88fb;
17'h20e5:	data_out=16'ha00;
17'h20e6:	data_out=16'h603;
17'h20e7:	data_out=16'h2cb;
17'h20e8:	data_out=16'h267;
17'h20e9:	data_out=16'h84e7;
17'h20ea:	data_out=16'h259;
17'h20eb:	data_out=16'ha00;
17'h20ec:	data_out=16'h820d;
17'h20ed:	data_out=16'h85a2;
17'h20ee:	data_out=16'h259;
17'h20ef:	data_out=16'ha00;
17'h20f0:	data_out=16'h25b;
17'h20f1:	data_out=16'h899c;
17'h20f2:	data_out=16'ha00;
17'h20f3:	data_out=16'ha00;
17'h20f4:	data_out=16'h9ff;
17'h20f5:	data_out=16'h5bc;
17'h20f6:	data_out=16'h80f2;
17'h20f7:	data_out=16'ha00;
17'h20f8:	data_out=16'ha00;
17'h20f9:	data_out=16'h81ae;
17'h20fa:	data_out=16'h84b2;
17'h20fb:	data_out=16'h261;
17'h20fc:	data_out=16'h8407;
17'h20fd:	data_out=16'h63a;
17'h20fe:	data_out=16'h666;
17'h20ff:	data_out=16'ha00;
17'h2100:	data_out=16'h871e;
17'h2101:	data_out=16'h1da;
17'h2102:	data_out=16'h814d;
17'h2103:	data_out=16'h9fd;
17'h2104:	data_out=16'ha00;
17'h2105:	data_out=16'ha00;
17'h2106:	data_out=16'ha00;
17'h2107:	data_out=16'h824;
17'h2108:	data_out=16'h82d8;
17'h2109:	data_out=16'h4;
17'h210a:	data_out=16'h281;
17'h210b:	data_out=16'h469;
17'h210c:	data_out=16'h9ff;
17'h210d:	data_out=16'h474;
17'h210e:	data_out=16'h1ae;
17'h210f:	data_out=16'h855c;
17'h2110:	data_out=16'ha00;
17'h2111:	data_out=16'h8f3;
17'h2112:	data_out=16'h86c6;
17'h2113:	data_out=16'h9f9;
17'h2114:	data_out=16'h895a;
17'h2115:	data_out=16'h262;
17'h2116:	data_out=16'ha00;
17'h2117:	data_out=16'h83d0;
17'h2118:	data_out=16'h8824;
17'h2119:	data_out=16'ha00;
17'h211a:	data_out=16'ha00;
17'h211b:	data_out=16'h814;
17'h211c:	data_out=16'h9f7;
17'h211d:	data_out=16'h451;
17'h211e:	data_out=16'h8829;
17'h211f:	data_out=16'h2c8;
17'h2120:	data_out=16'h921;
17'h2121:	data_out=16'h1c0;
17'h2122:	data_out=16'ha00;
17'h2123:	data_out=16'h83f4;
17'h2124:	data_out=16'h83ef;
17'h2125:	data_out=16'ha00;
17'h2126:	data_out=16'h8877;
17'h2127:	data_out=16'h418;
17'h2128:	data_out=16'h1da;
17'h2129:	data_out=16'h861d;
17'h212a:	data_out=16'h87c8;
17'h212b:	data_out=16'h8088;
17'h212c:	data_out=16'ha00;
17'h212d:	data_out=16'h9b6;
17'h212e:	data_out=16'h8111;
17'h212f:	data_out=16'ha00;
17'h2130:	data_out=16'ha00;
17'h2131:	data_out=16'h81ec;
17'h2132:	data_out=16'ha00;
17'h2133:	data_out=16'h89fc;
17'h2134:	data_out=16'h8893;
17'h2135:	data_out=16'h9fe;
17'h2136:	data_out=16'h84ed;
17'h2137:	data_out=16'h8118;
17'h2138:	data_out=16'h6f4;
17'h2139:	data_out=16'h89fb;
17'h213a:	data_out=16'h826e;
17'h213b:	data_out=16'ha00;
17'h213c:	data_out=16'h9fa;
17'h213d:	data_out=16'h823;
17'h213e:	data_out=16'h1da;
17'h213f:	data_out=16'ha00;
17'h2140:	data_out=16'ha00;
17'h2141:	data_out=16'h77e;
17'h2142:	data_out=16'h9fd;
17'h2143:	data_out=16'ha00;
17'h2144:	data_out=16'h7af;
17'h2145:	data_out=16'h2c3;
17'h2146:	data_out=16'h601;
17'h2147:	data_out=16'h90;
17'h2148:	data_out=16'h441;
17'h2149:	data_out=16'ha00;
17'h214a:	data_out=16'ha00;
17'h214b:	data_out=16'ha00;
17'h214c:	data_out=16'ha00;
17'h214d:	data_out=16'ha00;
17'h214e:	data_out=16'h329;
17'h214f:	data_out=16'h8be;
17'h2150:	data_out=16'ha00;
17'h2151:	data_out=16'h7a4;
17'h2152:	data_out=16'h82cd;
17'h2153:	data_out=16'ha00;
17'h2154:	data_out=16'ha00;
17'h2155:	data_out=16'h8105;
17'h2156:	data_out=16'h81c5;
17'h2157:	data_out=16'h81a5;
17'h2158:	data_out=16'h8085;
17'h2159:	data_out=16'ha00;
17'h215a:	data_out=16'h61e;
17'h215b:	data_out=16'h629;
17'h215c:	data_out=16'h9fc;
17'h215d:	data_out=16'ha00;
17'h215e:	data_out=16'ha00;
17'h215f:	data_out=16'h8336;
17'h2160:	data_out=16'h87f7;
17'h2161:	data_out=16'ha00;
17'h2162:	data_out=16'h859d;
17'h2163:	data_out=16'h89cb;
17'h2164:	data_out=16'h89fb;
17'h2165:	data_out=16'ha00;
17'h2166:	data_out=16'h996;
17'h2167:	data_out=16'h19f;
17'h2168:	data_out=16'h1cb;
17'h2169:	data_out=16'h84b8;
17'h216a:	data_out=16'h1a3;
17'h216b:	data_out=16'ha00;
17'h216c:	data_out=16'h1fb;
17'h216d:	data_out=16'h89d2;
17'h216e:	data_out=16'h1a3;
17'h216f:	data_out=16'ha00;
17'h2170:	data_out=16'h1aa;
17'h2171:	data_out=16'h89ff;
17'h2172:	data_out=16'ha00;
17'h2173:	data_out=16'ha00;
17'h2174:	data_out=16'h9ff;
17'h2175:	data_out=16'h9fd;
17'h2176:	data_out=16'h83ce;
17'h2177:	data_out=16'ha00;
17'h2178:	data_out=16'ha00;
17'h2179:	data_out=16'h8519;
17'h217a:	data_out=16'h893f;
17'h217b:	data_out=16'h1d9;
17'h217c:	data_out=16'h86c2;
17'h217d:	data_out=16'h881;
17'h217e:	data_out=16'h54d;
17'h217f:	data_out=16'ha00;
17'h2180:	data_out=16'h86b3;
17'h2181:	data_out=16'h813;
17'h2182:	data_out=16'hd7;
17'h2183:	data_out=16'h9ff;
17'h2184:	data_out=16'ha00;
17'h2185:	data_out=16'ha00;
17'h2186:	data_out=16'ha00;
17'h2187:	data_out=16'ha00;
17'h2188:	data_out=16'h1e9;
17'h2189:	data_out=16'h819b;
17'h218a:	data_out=16'ha00;
17'h218b:	data_out=16'h8ef;
17'h218c:	data_out=16'ha00;
17'h218d:	data_out=16'h56f;
17'h218e:	data_out=16'h129;
17'h218f:	data_out=16'h855f;
17'h2190:	data_out=16'ha00;
17'h2191:	data_out=16'h782;
17'h2192:	data_out=16'h892b;
17'h2193:	data_out=16'h9f6;
17'h2194:	data_out=16'h8996;
17'h2195:	data_out=16'h3ee;
17'h2196:	data_out=16'ha00;
17'h2197:	data_out=16'h8417;
17'h2198:	data_out=16'h8a00;
17'h2199:	data_out=16'ha00;
17'h219a:	data_out=16'ha00;
17'h219b:	data_out=16'h9f8;
17'h219c:	data_out=16'h9fb;
17'h219d:	data_out=16'h9f4;
17'h219e:	data_out=16'h88ea;
17'h219f:	data_out=16'h80cc;
17'h21a0:	data_out=16'ha00;
17'h21a1:	data_out=16'h145;
17'h21a2:	data_out=16'ha00;
17'h21a3:	data_out=16'h84be;
17'h21a4:	data_out=16'h84b9;
17'h21a5:	data_out=16'ha00;
17'h21a6:	data_out=16'h87a4;
17'h21a7:	data_out=16'h9f5;
17'h21a8:	data_out=16'h192;
17'h21a9:	data_out=16'h866e;
17'h21aa:	data_out=16'h87c4;
17'h21ab:	data_out=16'h323;
17'h21ac:	data_out=16'ha00;
17'h21ad:	data_out=16'h94b;
17'h21ae:	data_out=16'h109;
17'h21af:	data_out=16'ha00;
17'h21b0:	data_out=16'ha00;
17'h21b1:	data_out=16'h130;
17'h21b2:	data_out=16'ha00;
17'h21b3:	data_out=16'h89fe;
17'h21b4:	data_out=16'h8864;
17'h21b5:	data_out=16'ha00;
17'h21b6:	data_out=16'h822a;
17'h21b7:	data_out=16'h136;
17'h21b8:	data_out=16'h6c8;
17'h21b9:	data_out=16'h89fe;
17'h21ba:	data_out=16'h8638;
17'h21bb:	data_out=16'ha00;
17'h21bc:	data_out=16'h9fe;
17'h21bd:	data_out=16'h9d9;
17'h21be:	data_out=16'h197;
17'h21bf:	data_out=16'ha00;
17'h21c0:	data_out=16'ha00;
17'h21c1:	data_out=16'h9fc;
17'h21c2:	data_out=16'h9fe;
17'h21c3:	data_out=16'ha00;
17'h21c4:	data_out=16'h9f8;
17'h21c5:	data_out=16'h54c;
17'h21c6:	data_out=16'h78a;
17'h21c7:	data_out=16'h80cb;
17'h21c8:	data_out=16'h568;
17'h21c9:	data_out=16'ha00;
17'h21ca:	data_out=16'ha00;
17'h21cb:	data_out=16'ha00;
17'h21cc:	data_out=16'ha00;
17'h21cd:	data_out=16'ha00;
17'h21ce:	data_out=16'h8df;
17'h21cf:	data_out=16'h9dc;
17'h21d0:	data_out=16'ha00;
17'h21d1:	data_out=16'h517;
17'h21d2:	data_out=16'h830c;
17'h21d3:	data_out=16'ha00;
17'h21d4:	data_out=16'ha00;
17'h21d5:	data_out=16'h314;
17'h21d6:	data_out=16'h851d;
17'h21d7:	data_out=16'h8559;
17'h21d8:	data_out=16'h3dc;
17'h21d9:	data_out=16'ha00;
17'h21da:	data_out=16'h77f;
17'h21db:	data_out=16'h9f8;
17'h21dc:	data_out=16'ha00;
17'h21dd:	data_out=16'ha00;
17'h21de:	data_out=16'ha00;
17'h21df:	data_out=16'h843a;
17'h21e0:	data_out=16'h880b;
17'h21e1:	data_out=16'ha00;
17'h21e2:	data_out=16'h839e;
17'h21e3:	data_out=16'h89f9;
17'h21e4:	data_out=16'h89fc;
17'h21e5:	data_out=16'ha00;
17'h21e6:	data_out=16'ha00;
17'h21e7:	data_out=16'h539;
17'h21e8:	data_out=16'h157;
17'h21e9:	data_out=16'h8143;
17'h21ea:	data_out=16'h112;
17'h21eb:	data_out=16'ha00;
17'h21ec:	data_out=16'h8a4;
17'h21ed:	data_out=16'h89fd;
17'h21ee:	data_out=16'h113;
17'h21ef:	data_out=16'ha00;
17'h21f0:	data_out=16'h120;
17'h21f1:	data_out=16'h8a00;
17'h21f2:	data_out=16'ha00;
17'h21f3:	data_out=16'ha00;
17'h21f4:	data_out=16'ha00;
17'h21f5:	data_out=16'h9ff;
17'h21f6:	data_out=16'h8276;
17'h21f7:	data_out=16'ha00;
17'h21f8:	data_out=16'ha00;
17'h21f9:	data_out=16'h83e8;
17'h21fa:	data_out=16'h8982;
17'h21fb:	data_out=16'h198;
17'h21fc:	data_out=16'h8902;
17'h21fd:	data_out=16'h8c0;
17'h21fe:	data_out=16'h703;
17'h21ff:	data_out=16'ha00;
17'h2200:	data_out=16'h8125;
17'h2201:	data_out=16'h9f3;
17'h2202:	data_out=16'h8299;
17'h2203:	data_out=16'h9ff;
17'h2204:	data_out=16'ha00;
17'h2205:	data_out=16'ha00;
17'h2206:	data_out=16'ha00;
17'h2207:	data_out=16'ha00;
17'h2208:	data_out=16'h81f2;
17'h2209:	data_out=16'h8015;
17'h220a:	data_out=16'h9fb;
17'h220b:	data_out=16'h7d6;
17'h220c:	data_out=16'ha00;
17'h220d:	data_out=16'h85a;
17'h220e:	data_out=16'hfa;
17'h220f:	data_out=16'h897f;
17'h2210:	data_out=16'ha00;
17'h2211:	data_out=16'h89d;
17'h2212:	data_out=16'h8a00;
17'h2213:	data_out=16'h9e4;
17'h2214:	data_out=16'h89a8;
17'h2215:	data_out=16'h943;
17'h2216:	data_out=16'ha00;
17'h2217:	data_out=16'h83e0;
17'h2218:	data_out=16'h8a00;
17'h2219:	data_out=16'ha00;
17'h221a:	data_out=16'ha00;
17'h221b:	data_out=16'h8c8;
17'h221c:	data_out=16'h9f1;
17'h221d:	data_out=16'h9eb;
17'h221e:	data_out=16'h883b;
17'h221f:	data_out=16'h81fd;
17'h2220:	data_out=16'h9f7;
17'h2221:	data_out=16'h141;
17'h2222:	data_out=16'ha00;
17'h2223:	data_out=16'h89d9;
17'h2224:	data_out=16'h89d2;
17'h2225:	data_out=16'ha00;
17'h2226:	data_out=16'h8a00;
17'h2227:	data_out=16'h9ef;
17'h2228:	data_out=16'h1a7;
17'h2229:	data_out=16'h8473;
17'h222a:	data_out=16'h88d8;
17'h222b:	data_out=16'h515;
17'h222c:	data_out=16'ha00;
17'h222d:	data_out=16'h725;
17'h222e:	data_out=16'h8065;
17'h222f:	data_out=16'ha00;
17'h2230:	data_out=16'ha00;
17'h2231:	data_out=16'h5c3;
17'h2232:	data_out=16'ha00;
17'h2233:	data_out=16'h8a00;
17'h2234:	data_out=16'h88b7;
17'h2235:	data_out=16'h9f9;
17'h2236:	data_out=16'h8426;
17'h2237:	data_out=16'h81da;
17'h2238:	data_out=16'h9b1;
17'h2239:	data_out=16'h89ff;
17'h223a:	data_out=16'h85a0;
17'h223b:	data_out=16'ha00;
17'h223c:	data_out=16'h9f5;
17'h223d:	data_out=16'h9f9;
17'h223e:	data_out=16'h1ab;
17'h223f:	data_out=16'ha00;
17'h2240:	data_out=16'ha00;
17'h2241:	data_out=16'h9f5;
17'h2242:	data_out=16'h9fe;
17'h2243:	data_out=16'ha00;
17'h2244:	data_out=16'h9f0;
17'h2245:	data_out=16'ha00;
17'h2246:	data_out=16'h3b3;
17'h2247:	data_out=16'h807f;
17'h2248:	data_out=16'h8b0;
17'h2249:	data_out=16'ha00;
17'h224a:	data_out=16'ha00;
17'h224b:	data_out=16'ha00;
17'h224c:	data_out=16'ha00;
17'h224d:	data_out=16'ha00;
17'h224e:	data_out=16'h8b9;
17'h224f:	data_out=16'ha00;
17'h2250:	data_out=16'ha00;
17'h2251:	data_out=16'h198;
17'h2252:	data_out=16'h872e;
17'h2253:	data_out=16'h9f8;
17'h2254:	data_out=16'h9f7;
17'h2255:	data_out=16'h1ac;
17'h2256:	data_out=16'h8796;
17'h2257:	data_out=16'h8550;
17'h2258:	data_out=16'h1ad;
17'h2259:	data_out=16'ha00;
17'h225a:	data_out=16'h495;
17'h225b:	data_out=16'h9ee;
17'h225c:	data_out=16'h9f7;
17'h225d:	data_out=16'ha00;
17'h225e:	data_out=16'ha00;
17'h225f:	data_out=16'h8429;
17'h2260:	data_out=16'h89ff;
17'h2261:	data_out=16'ha00;
17'h2262:	data_out=16'h8577;
17'h2263:	data_out=16'h89fa;
17'h2264:	data_out=16'h89fd;
17'h2265:	data_out=16'ha00;
17'h2266:	data_out=16'ha00;
17'h2267:	data_out=16'h9fa;
17'h2268:	data_out=16'h165;
17'h2269:	data_out=16'h8588;
17'h226a:	data_out=16'hcd;
17'h226b:	data_out=16'ha00;
17'h226c:	data_out=16'h950;
17'h226d:	data_out=16'h89fe;
17'h226e:	data_out=16'hce;
17'h226f:	data_out=16'ha00;
17'h2270:	data_out=16'he4;
17'h2271:	data_out=16'h8a00;
17'h2272:	data_out=16'ha00;
17'h2273:	data_out=16'ha00;
17'h2274:	data_out=16'ha00;
17'h2275:	data_out=16'h9fe;
17'h2276:	data_out=16'h80f9;
17'h2277:	data_out=16'ha00;
17'h2278:	data_out=16'ha00;
17'h2279:	data_out=16'h870e;
17'h227a:	data_out=16'h8996;
17'h227b:	data_out=16'h1ad;
17'h227c:	data_out=16'h8a00;
17'h227d:	data_out=16'h9fa;
17'h227e:	data_out=16'ha00;
17'h227f:	data_out=16'ha00;
17'h2280:	data_out=16'h8ce;
17'h2281:	data_out=16'h9dd;
17'h2282:	data_out=16'h84ac;
17'h2283:	data_out=16'ha00;
17'h2284:	data_out=16'ha00;
17'h2285:	data_out=16'ha00;
17'h2286:	data_out=16'ha00;
17'h2287:	data_out=16'ha00;
17'h2288:	data_out=16'h8a00;
17'h2289:	data_out=16'h82b7;
17'h228a:	data_out=16'h9f1;
17'h228b:	data_out=16'h727;
17'h228c:	data_out=16'ha00;
17'h228d:	data_out=16'h9e6;
17'h228e:	data_out=16'h68;
17'h228f:	data_out=16'h8922;
17'h2290:	data_out=16'ha00;
17'h2291:	data_out=16'h7d3;
17'h2292:	data_out=16'h8a00;
17'h2293:	data_out=16'h9f0;
17'h2294:	data_out=16'h851c;
17'h2295:	data_out=16'ha00;
17'h2296:	data_out=16'ha00;
17'h2297:	data_out=16'h7fe;
17'h2298:	data_out=16'h8a00;
17'h2299:	data_out=16'ha00;
17'h229a:	data_out=16'ha00;
17'h229b:	data_out=16'h7c6;
17'h229c:	data_out=16'h9db;
17'h229d:	data_out=16'h9a8;
17'h229e:	data_out=16'h2a4;
17'h229f:	data_out=16'h1be;
17'h22a0:	data_out=16'h9f7;
17'h22a1:	data_out=16'hbf;
17'h22a2:	data_out=16'ha00;
17'h22a3:	data_out=16'h89f1;
17'h22a4:	data_out=16'h89f1;
17'h22a5:	data_out=16'h9ff;
17'h22a6:	data_out=16'h8a00;
17'h22a7:	data_out=16'h9de;
17'h22a8:	data_out=16'h11d;
17'h22a9:	data_out=16'h20a;
17'h22aa:	data_out=16'h88f9;
17'h22ab:	data_out=16'h85f0;
17'h22ac:	data_out=16'ha00;
17'h22ad:	data_out=16'h3e0;
17'h22ae:	data_out=16'h6a;
17'h22af:	data_out=16'ha00;
17'h22b0:	data_out=16'ha00;
17'h22b1:	data_out=16'h9d9;
17'h22b2:	data_out=16'ha00;
17'h22b3:	data_out=16'h88b0;
17'h22b4:	data_out=16'h873c;
17'h22b5:	data_out=16'h9fa;
17'h22b6:	data_out=16'h872e;
17'h22b7:	data_out=16'h82d6;
17'h22b8:	data_out=16'h9b8;
17'h22b9:	data_out=16'h8979;
17'h22ba:	data_out=16'h84a9;
17'h22bb:	data_out=16'ha00;
17'h22bc:	data_out=16'h9e5;
17'h22bd:	data_out=16'h9fd;
17'h22be:	data_out=16'h122;
17'h22bf:	data_out=16'ha00;
17'h22c0:	data_out=16'ha00;
17'h22c1:	data_out=16'h9f2;
17'h22c2:	data_out=16'h9fe;
17'h22c3:	data_out=16'ha00;
17'h22c4:	data_out=16'h9e0;
17'h22c5:	data_out=16'ha00;
17'h22c6:	data_out=16'h81a5;
17'h22c7:	data_out=16'h8052;
17'h22c8:	data_out=16'h778;
17'h22c9:	data_out=16'ha00;
17'h22ca:	data_out=16'ha00;
17'h22cb:	data_out=16'ha00;
17'h22cc:	data_out=16'h9ff;
17'h22cd:	data_out=16'ha00;
17'h22ce:	data_out=16'h7f0;
17'h22cf:	data_out=16'h9ff;
17'h22d0:	data_out=16'ha00;
17'h22d1:	data_out=16'h4ca;
17'h22d2:	data_out=16'h897e;
17'h22d3:	data_out=16'h9f4;
17'h22d4:	data_out=16'h9f0;
17'h22d5:	data_out=16'h63d;
17'h22d6:	data_out=16'h8854;
17'h22d7:	data_out=16'h85a5;
17'h22d8:	data_out=16'h146;
17'h22d9:	data_out=16'ha00;
17'h22da:	data_out=16'h4a6;
17'h22db:	data_out=16'h9e3;
17'h22dc:	data_out=16'h9e6;
17'h22dd:	data_out=16'ha00;
17'h22de:	data_out=16'ha00;
17'h22df:	data_out=16'h838a;
17'h22e0:	data_out=16'h8a00;
17'h22e1:	data_out=16'ha00;
17'h22e2:	data_out=16'h1dd;
17'h22e3:	data_out=16'h873d;
17'h22e4:	data_out=16'h89ff;
17'h22e5:	data_out=16'ha00;
17'h22e6:	data_out=16'ha00;
17'h22e7:	data_out=16'ha00;
17'h22e8:	data_out=16'hec;
17'h22e9:	data_out=16'h8a00;
17'h22ea:	data_out=16'h2c;
17'h22eb:	data_out=16'ha00;
17'h22ec:	data_out=16'h9d3;
17'h22ed:	data_out=16'h86ed;
17'h22ee:	data_out=16'h2e;
17'h22ef:	data_out=16'ha00;
17'h22f0:	data_out=16'h4a;
17'h22f1:	data_out=16'h89ff;
17'h22f2:	data_out=16'ha00;
17'h22f3:	data_out=16'ha00;
17'h22f4:	data_out=16'ha00;
17'h22f5:	data_out=16'h9fa;
17'h22f6:	data_out=16'h8709;
17'h22f7:	data_out=16'ha00;
17'h22f8:	data_out=16'ha00;
17'h22f9:	data_out=16'h8536;
17'h22fa:	data_out=16'h85a1;
17'h22fb:	data_out=16'h124;
17'h22fc:	data_out=16'h8a00;
17'h22fd:	data_out=16'ha00;
17'h22fe:	data_out=16'h9f0;
17'h22ff:	data_out=16'ha00;
17'h2300:	data_out=16'h7c1;
17'h2301:	data_out=16'h9e6;
17'h2302:	data_out=16'h3cb;
17'h2303:	data_out=16'ha00;
17'h2304:	data_out=16'ha00;
17'h2305:	data_out=16'ha00;
17'h2306:	data_out=16'ha00;
17'h2307:	data_out=16'ha00;
17'h2308:	data_out=16'h8a00;
17'h2309:	data_out=16'h809e;
17'h230a:	data_out=16'h9fc;
17'h230b:	data_out=16'h923;
17'h230c:	data_out=16'ha00;
17'h230d:	data_out=16'h9fb;
17'h230e:	data_out=16'h1e2;
17'h230f:	data_out=16'h226;
17'h2310:	data_out=16'ha00;
17'h2311:	data_out=16'h7cb;
17'h2312:	data_out=16'h8894;
17'h2313:	data_out=16'h9fc;
17'h2314:	data_out=16'h856;
17'h2315:	data_out=16'ha00;
17'h2316:	data_out=16'ha00;
17'h2317:	data_out=16'h9fc;
17'h2318:	data_out=16'h8a00;
17'h2319:	data_out=16'ha00;
17'h231a:	data_out=16'ha00;
17'h231b:	data_out=16'h9d9;
17'h231c:	data_out=16'h9ef;
17'h231d:	data_out=16'h99d;
17'h231e:	data_out=16'h9f5;
17'h231f:	data_out=16'h9f4;
17'h2320:	data_out=16'h9fa;
17'h2321:	data_out=16'h234;
17'h2322:	data_out=16'ha00;
17'h2323:	data_out=16'h89fc;
17'h2324:	data_out=16'h89fb;
17'h2325:	data_out=16'ha00;
17'h2326:	data_out=16'h8a00;
17'h2327:	data_out=16'h9ec;
17'h2328:	data_out=16'h2a4;
17'h2329:	data_out=16'h3c3;
17'h232a:	data_out=16'h8201;
17'h232b:	data_out=16'h8a00;
17'h232c:	data_out=16'ha00;
17'h232d:	data_out=16'h311;
17'h232e:	data_out=16'h7ce;
17'h232f:	data_out=16'ha00;
17'h2330:	data_out=16'ha00;
17'h2331:	data_out=16'h9e8;
17'h2332:	data_out=16'ha00;
17'h2333:	data_out=16'h4bc;
17'h2334:	data_out=16'h8796;
17'h2335:	data_out=16'ha00;
17'h2336:	data_out=16'h85fb;
17'h2337:	data_out=16'h59e;
17'h2338:	data_out=16'h82d;
17'h2339:	data_out=16'h347;
17'h233a:	data_out=16'h8364;
17'h233b:	data_out=16'ha00;
17'h233c:	data_out=16'h9f5;
17'h233d:	data_out=16'h9fc;
17'h233e:	data_out=16'h2ab;
17'h233f:	data_out=16'ha00;
17'h2340:	data_out=16'ha00;
17'h2341:	data_out=16'h9f9;
17'h2342:	data_out=16'h9fe;
17'h2343:	data_out=16'ha00;
17'h2344:	data_out=16'h9ee;
17'h2345:	data_out=16'ha00;
17'h2346:	data_out=16'h874a;
17'h2347:	data_out=16'h269;
17'h2348:	data_out=16'ha00;
17'h2349:	data_out=16'ha00;
17'h234a:	data_out=16'ha00;
17'h234b:	data_out=16'ha00;
17'h234c:	data_out=16'ha00;
17'h234d:	data_out=16'ha00;
17'h234e:	data_out=16'h81d;
17'h234f:	data_out=16'h9fe;
17'h2350:	data_out=16'ha00;
17'h2351:	data_out=16'h7a4;
17'h2352:	data_out=16'h8980;
17'h2353:	data_out=16'h9fc;
17'h2354:	data_out=16'h9f7;
17'h2355:	data_out=16'h9f5;
17'h2356:	data_out=16'h81ee;
17'h2357:	data_out=16'h4c;
17'h2358:	data_out=16'h4a9;
17'h2359:	data_out=16'ha00;
17'h235a:	data_out=16'h7ca;
17'h235b:	data_out=16'h9e8;
17'h235c:	data_out=16'h9f8;
17'h235d:	data_out=16'ha00;
17'h235e:	data_out=16'ha00;
17'h235f:	data_out=16'h823b;
17'h2360:	data_out=16'h8a00;
17'h2361:	data_out=16'ha00;
17'h2362:	data_out=16'h9fd;
17'h2363:	data_out=16'h629;
17'h2364:	data_out=16'h8a00;
17'h2365:	data_out=16'ha00;
17'h2366:	data_out=16'ha00;
17'h2367:	data_out=16'ha00;
17'h2368:	data_out=16'h263;
17'h2369:	data_out=16'h8a00;
17'h236a:	data_out=16'h1a9;
17'h236b:	data_out=16'ha00;
17'h236c:	data_out=16'h93f;
17'h236d:	data_out=16'h676;
17'h236e:	data_out=16'h1ab;
17'h236f:	data_out=16'ha00;
17'h2370:	data_out=16'h1c9;
17'h2371:	data_out=16'h89e4;
17'h2372:	data_out=16'ha00;
17'h2373:	data_out=16'ha00;
17'h2374:	data_out=16'ha00;
17'h2375:	data_out=16'h9ff;
17'h2376:	data_out=16'h89fc;
17'h2377:	data_out=16'ha00;
17'h2378:	data_out=16'ha00;
17'h2379:	data_out=16'h573;
17'h237a:	data_out=16'h7b3;
17'h237b:	data_out=16'h2ae;
17'h237c:	data_out=16'h8a00;
17'h237d:	data_out=16'ha00;
17'h237e:	data_out=16'h9f5;
17'h237f:	data_out=16'ha00;
17'h2380:	data_out=16'h9f4;
17'h2381:	data_out=16'h9ff;
17'h2382:	data_out=16'h4ed;
17'h2383:	data_out=16'ha00;
17'h2384:	data_out=16'ha00;
17'h2385:	data_out=16'ha00;
17'h2386:	data_out=16'ha00;
17'h2387:	data_out=16'h9d7;
17'h2388:	data_out=16'h89f0;
17'h2389:	data_out=16'h83f6;
17'h238a:	data_out=16'ha00;
17'h238b:	data_out=16'h9aa;
17'h238c:	data_out=16'ha00;
17'h238d:	data_out=16'ha00;
17'h238e:	data_out=16'h23d;
17'h238f:	data_out=16'h3dd;
17'h2390:	data_out=16'ha00;
17'h2391:	data_out=16'h89f;
17'h2392:	data_out=16'h8674;
17'h2393:	data_out=16'ha00;
17'h2394:	data_out=16'ha00;
17'h2395:	data_out=16'ha00;
17'h2396:	data_out=16'ha00;
17'h2397:	data_out=16'ha00;
17'h2398:	data_out=16'h8a00;
17'h2399:	data_out=16'ha00;
17'h239a:	data_out=16'ha00;
17'h239b:	data_out=16'h9ff;
17'h239c:	data_out=16'ha00;
17'h239d:	data_out=16'h9fb;
17'h239e:	data_out=16'ha00;
17'h239f:	data_out=16'h9fe;
17'h23a0:	data_out=16'ha00;
17'h23a1:	data_out=16'h286;
17'h23a2:	data_out=16'ha00;
17'h23a3:	data_out=16'h8a00;
17'h23a4:	data_out=16'h8a00;
17'h23a5:	data_out=16'h676;
17'h23a6:	data_out=16'h89fa;
17'h23a7:	data_out=16'h9ff;
17'h23a8:	data_out=16'h2e0;
17'h23a9:	data_out=16'h228;
17'h23aa:	data_out=16'h81e2;
17'h23ab:	data_out=16'h89fc;
17'h23ac:	data_out=16'ha00;
17'h23ad:	data_out=16'h6d;
17'h23ae:	data_out=16'h84a;
17'h23af:	data_out=16'ha00;
17'h23b0:	data_out=16'ha00;
17'h23b1:	data_out=16'h9ff;
17'h23b2:	data_out=16'ha00;
17'h23b3:	data_out=16'h9fe;
17'h23b4:	data_out=16'h8361;
17'h23b5:	data_out=16'ha00;
17'h23b6:	data_out=16'h8834;
17'h23b7:	data_out=16'h6c8;
17'h23b8:	data_out=16'h983;
17'h23b9:	data_out=16'h9fd;
17'h23ba:	data_out=16'h867d;
17'h23bb:	data_out=16'ha00;
17'h23bc:	data_out=16'ha00;
17'h23bd:	data_out=16'ha00;
17'h23be:	data_out=16'h2e5;
17'h23bf:	data_out=16'ha00;
17'h23c0:	data_out=16'ha00;
17'h23c1:	data_out=16'ha00;
17'h23c2:	data_out=16'ha00;
17'h23c3:	data_out=16'ha00;
17'h23c4:	data_out=16'h9ff;
17'h23c5:	data_out=16'ha00;
17'h23c6:	data_out=16'h8757;
17'h23c7:	data_out=16'h85f3;
17'h23c8:	data_out=16'h6be;
17'h23c9:	data_out=16'h6e2;
17'h23ca:	data_out=16'ha00;
17'h23cb:	data_out=16'ha00;
17'h23cc:	data_out=16'h8111;
17'h23cd:	data_out=16'ha00;
17'h23ce:	data_out=16'h8e3;
17'h23cf:	data_out=16'h83a7;
17'h23d0:	data_out=16'ha00;
17'h23d1:	data_out=16'h9fd;
17'h23d2:	data_out=16'h89f3;
17'h23d3:	data_out=16'h9ff;
17'h23d4:	data_out=16'h9ff;
17'h23d5:	data_out=16'h9ff;
17'h23d6:	data_out=16'h84d9;
17'h23d7:	data_out=16'h8209;
17'h23d8:	data_out=16'h879;
17'h23d9:	data_out=16'ha00;
17'h23da:	data_out=16'h9fc;
17'h23db:	data_out=16'h9fc;
17'h23dc:	data_out=16'ha00;
17'h23dd:	data_out=16'ha00;
17'h23de:	data_out=16'ha00;
17'h23df:	data_out=16'h81ee;
17'h23e0:	data_out=16'h89f2;
17'h23e1:	data_out=16'ha00;
17'h23e2:	data_out=16'ha00;
17'h23e3:	data_out=16'h9ff;
17'h23e4:	data_out=16'h89f8;
17'h23e5:	data_out=16'ha00;
17'h23e6:	data_out=16'h9ff;
17'h23e7:	data_out=16'h844;
17'h23e8:	data_out=16'h2ae;
17'h23e9:	data_out=16'h8a00;
17'h23ea:	data_out=16'h207;
17'h23eb:	data_out=16'ha00;
17'h23ec:	data_out=16'h9fd;
17'h23ed:	data_out=16'h9ff;
17'h23ee:	data_out=16'h208;
17'h23ef:	data_out=16'ha00;
17'h23f0:	data_out=16'h226;
17'h23f1:	data_out=16'h88c7;
17'h23f2:	data_out=16'ha00;
17'h23f3:	data_out=16'ha00;
17'h23f4:	data_out=16'ha00;
17'h23f5:	data_out=16'ha00;
17'h23f6:	data_out=16'h89fb;
17'h23f7:	data_out=16'ha00;
17'h23f8:	data_out=16'ha00;
17'h23f9:	data_out=16'h5de;
17'h23fa:	data_out=16'ha00;
17'h23fb:	data_out=16'h2e8;
17'h23fc:	data_out=16'h8a00;
17'h23fd:	data_out=16'ha00;
17'h23fe:	data_out=16'h9e6;
17'h23ff:	data_out=16'ha00;
17'h2400:	data_out=16'h9f1;
17'h2401:	data_out=16'ha00;
17'h2402:	data_out=16'h9ff;
17'h2403:	data_out=16'ha00;
17'h2404:	data_out=16'ha00;
17'h2405:	data_out=16'ha00;
17'h2406:	data_out=16'ha00;
17'h2407:	data_out=16'h9ff;
17'h2408:	data_out=16'h6df;
17'h2409:	data_out=16'h83e9;
17'h240a:	data_out=16'ha00;
17'h240b:	data_out=16'h9fe;
17'h240c:	data_out=16'ha00;
17'h240d:	data_out=16'ha00;
17'h240e:	data_out=16'h3ef;
17'h240f:	data_out=16'ha00;
17'h2410:	data_out=16'ha00;
17'h2411:	data_out=16'h92b;
17'h2412:	data_out=16'h2e;
17'h2413:	data_out=16'ha00;
17'h2414:	data_out=16'ha00;
17'h2415:	data_out=16'ha00;
17'h2416:	data_out=16'ha00;
17'h2417:	data_out=16'ha00;
17'h2418:	data_out=16'h8a00;
17'h2419:	data_out=16'ha00;
17'h241a:	data_out=16'ha00;
17'h241b:	data_out=16'ha00;
17'h241c:	data_out=16'ha00;
17'h241d:	data_out=16'ha00;
17'h241e:	data_out=16'ha00;
17'h241f:	data_out=16'ha00;
17'h2420:	data_out=16'ha00;
17'h2421:	data_out=16'h43b;
17'h2422:	data_out=16'ha00;
17'h2423:	data_out=16'h89ff;
17'h2424:	data_out=16'h89ff;
17'h2425:	data_out=16'h9f7;
17'h2426:	data_out=16'h3c9;
17'h2427:	data_out=16'ha00;
17'h2428:	data_out=16'h4b1;
17'h2429:	data_out=16'h3fa;
17'h242a:	data_out=16'ha00;
17'h242b:	data_out=16'h81b3;
17'h242c:	data_out=16'ha00;
17'h242d:	data_out=16'h4f1;
17'h242e:	data_out=16'ha00;
17'h242f:	data_out=16'ha00;
17'h2430:	data_out=16'ha00;
17'h2431:	data_out=16'ha00;
17'h2432:	data_out=16'ha00;
17'h2433:	data_out=16'ha00;
17'h2434:	data_out=16'h98;
17'h2435:	data_out=16'ha00;
17'h2436:	data_out=16'h992;
17'h2437:	data_out=16'h9ff;
17'h2438:	data_out=16'h9c1;
17'h2439:	data_out=16'ha00;
17'h243a:	data_out=16'h85fc;
17'h243b:	data_out=16'ha00;
17'h243c:	data_out=16'ha00;
17'h243d:	data_out=16'ha00;
17'h243e:	data_out=16'h4b7;
17'h243f:	data_out=16'ha00;
17'h2440:	data_out=16'ha00;
17'h2441:	data_out=16'ha00;
17'h2442:	data_out=16'h9ff;
17'h2443:	data_out=16'ha00;
17'h2444:	data_out=16'ha00;
17'h2445:	data_out=16'ha00;
17'h2446:	data_out=16'h399;
17'h2447:	data_out=16'h1a8;
17'h2448:	data_out=16'ha00;
17'h2449:	data_out=16'h9e9;
17'h244a:	data_out=16'ha00;
17'h244b:	data_out=16'h9ff;
17'h244c:	data_out=16'h625;
17'h244d:	data_out=16'ha00;
17'h244e:	data_out=16'h9ee;
17'h244f:	data_out=16'h346;
17'h2450:	data_out=16'ha00;
17'h2451:	data_out=16'ha00;
17'h2452:	data_out=16'h899b;
17'h2453:	data_out=16'ha00;
17'h2454:	data_out=16'ha00;
17'h2455:	data_out=16'ha00;
17'h2456:	data_out=16'h608;
17'h2457:	data_out=16'h443;
17'h2458:	data_out=16'ha00;
17'h2459:	data_out=16'ha00;
17'h245a:	data_out=16'ha00;
17'h245b:	data_out=16'h9ff;
17'h245c:	data_out=16'ha00;
17'h245d:	data_out=16'ha00;
17'h245e:	data_out=16'ha00;
17'h245f:	data_out=16'h22;
17'h2460:	data_out=16'h82b8;
17'h2461:	data_out=16'ha00;
17'h2462:	data_out=16'ha00;
17'h2463:	data_out=16'ha00;
17'h2464:	data_out=16'h8a00;
17'h2465:	data_out=16'ha00;
17'h2466:	data_out=16'ha00;
17'h2467:	data_out=16'h9dc;
17'h2468:	data_out=16'h468;
17'h2469:	data_out=16'hd0;
17'h246a:	data_out=16'h3b5;
17'h246b:	data_out=16'ha00;
17'h246c:	data_out=16'ha00;
17'h246d:	data_out=16'ha00;
17'h246e:	data_out=16'h3b7;
17'h246f:	data_out=16'ha00;
17'h2470:	data_out=16'h3d8;
17'h2471:	data_out=16'h8498;
17'h2472:	data_out=16'ha00;
17'h2473:	data_out=16'ha00;
17'h2474:	data_out=16'ha00;
17'h2475:	data_out=16'ha00;
17'h2476:	data_out=16'h8a00;
17'h2477:	data_out=16'ha00;
17'h2478:	data_out=16'ha00;
17'h2479:	data_out=16'h9c9;
17'h247a:	data_out=16'ha00;
17'h247b:	data_out=16'h4ba;
17'h247c:	data_out=16'h89b2;
17'h247d:	data_out=16'h9ff;
17'h247e:	data_out=16'h9fe;
17'h247f:	data_out=16'ha00;
17'h2480:	data_out=16'h9cd;
17'h2481:	data_out=16'ha00;
17'h2482:	data_out=16'ha00;
17'h2483:	data_out=16'ha00;
17'h2484:	data_out=16'ha00;
17'h2485:	data_out=16'ha00;
17'h2486:	data_out=16'ha00;
17'h2487:	data_out=16'ha00;
17'h2488:	data_out=16'ha00;
17'h2489:	data_out=16'hdc;
17'h248a:	data_out=16'ha00;
17'h248b:	data_out=16'h9fc;
17'h248c:	data_out=16'ha00;
17'h248d:	data_out=16'ha00;
17'h248e:	data_out=16'h610;
17'h248f:	data_out=16'ha00;
17'h2490:	data_out=16'ha00;
17'h2491:	data_out=16'h9b0;
17'h2492:	data_out=16'h848;
17'h2493:	data_out=16'ha00;
17'h2494:	data_out=16'ha00;
17'h2495:	data_out=16'ha00;
17'h2496:	data_out=16'ha00;
17'h2497:	data_out=16'ha00;
17'h2498:	data_out=16'h8583;
17'h2499:	data_out=16'h9c3;
17'h249a:	data_out=16'ha00;
17'h249b:	data_out=16'ha00;
17'h249c:	data_out=16'ha00;
17'h249d:	data_out=16'ha00;
17'h249e:	data_out=16'ha00;
17'h249f:	data_out=16'h9fb;
17'h24a0:	data_out=16'h9ff;
17'h24a1:	data_out=16'h651;
17'h24a2:	data_out=16'ha00;
17'h24a3:	data_out=16'h8373;
17'h24a4:	data_out=16'h8379;
17'h24a5:	data_out=16'ha00;
17'h24a6:	data_out=16'ha00;
17'h24a7:	data_out=16'ha00;
17'h24a8:	data_out=16'h6f9;
17'h24a9:	data_out=16'h80a;
17'h24aa:	data_out=16'ha00;
17'h24ab:	data_out=16'h8072;
17'h24ac:	data_out=16'ha00;
17'h24ad:	data_out=16'h758;
17'h24ae:	data_out=16'ha00;
17'h24af:	data_out=16'ha00;
17'h24b0:	data_out=16'ha00;
17'h24b1:	data_out=16'ha00;
17'h24b2:	data_out=16'ha00;
17'h24b3:	data_out=16'ha00;
17'h24b4:	data_out=16'h3ea;
17'h24b5:	data_out=16'ha00;
17'h24b6:	data_out=16'ha00;
17'h24b7:	data_out=16'ha00;
17'h24b8:	data_out=16'h9c8;
17'h24b9:	data_out=16'h96c;
17'h24ba:	data_out=16'h83bd;
17'h24bb:	data_out=16'ha00;
17'h24bc:	data_out=16'ha00;
17'h24bd:	data_out=16'h9ff;
17'h24be:	data_out=16'h702;
17'h24bf:	data_out=16'ha00;
17'h24c0:	data_out=16'ha00;
17'h24c1:	data_out=16'ha00;
17'h24c2:	data_out=16'ha00;
17'h24c3:	data_out=16'ha00;
17'h24c4:	data_out=16'ha00;
17'h24c5:	data_out=16'ha00;
17'h24c6:	data_out=16'ha00;
17'h24c7:	data_out=16'h6ab;
17'h24c8:	data_out=16'ha00;
17'h24c9:	data_out=16'ha00;
17'h24ca:	data_out=16'ha00;
17'h24cb:	data_out=16'ha00;
17'h24cc:	data_out=16'h9fc;
17'h24cd:	data_out=16'ha00;
17'h24ce:	data_out=16'ha00;
17'h24cf:	data_out=16'h9da;
17'h24d0:	data_out=16'ha00;
17'h24d1:	data_out=16'ha00;
17'h24d2:	data_out=16'h80a0;
17'h24d3:	data_out=16'ha00;
17'h24d4:	data_out=16'ha00;
17'h24d5:	data_out=16'ha00;
17'h24d6:	data_out=16'ha00;
17'h24d7:	data_out=16'h754;
17'h24d8:	data_out=16'ha00;
17'h24d9:	data_out=16'ha00;
17'h24da:	data_out=16'ha00;
17'h24db:	data_out=16'h9fa;
17'h24dc:	data_out=16'ha00;
17'h24dd:	data_out=16'ha00;
17'h24de:	data_out=16'ha00;
17'h24df:	data_out=16'h2e1;
17'h24e0:	data_out=16'ha00;
17'h24e1:	data_out=16'ha00;
17'h24e2:	data_out=16'ha00;
17'h24e3:	data_out=16'ha00;
17'h24e4:	data_out=16'h880c;
17'h24e5:	data_out=16'ha00;
17'h24e6:	data_out=16'ha00;
17'h24e7:	data_out=16'h977;
17'h24e8:	data_out=16'h683;
17'h24e9:	data_out=16'h911;
17'h24ea:	data_out=16'h5e2;
17'h24eb:	data_out=16'ha00;
17'h24ec:	data_out=16'ha00;
17'h24ed:	data_out=16'ha00;
17'h24ee:	data_out=16'h5e3;
17'h24ef:	data_out=16'ha00;
17'h24f0:	data_out=16'h5ff;
17'h24f1:	data_out=16'h2c6;
17'h24f2:	data_out=16'ha00;
17'h24f3:	data_out=16'ha00;
17'h24f4:	data_out=16'ha00;
17'h24f5:	data_out=16'ha00;
17'h24f6:	data_out=16'h8945;
17'h24f7:	data_out=16'ha00;
17'h24f8:	data_out=16'ha00;
17'h24f9:	data_out=16'ha00;
17'h24fa:	data_out=16'ha00;
17'h24fb:	data_out=16'h706;
17'h24fc:	data_out=16'h852a;
17'h24fd:	data_out=16'h97f;
17'h24fe:	data_out=16'h9ff;
17'h24ff:	data_out=16'ha00;
17'h2500:	data_out=16'h10b;
17'h2501:	data_out=16'ha00;
17'h2502:	data_out=16'ha00;
17'h2503:	data_out=16'ha00;
17'h2504:	data_out=16'ha00;
17'h2505:	data_out=16'ha00;
17'h2506:	data_out=16'ha00;
17'h2507:	data_out=16'ha00;
17'h2508:	data_out=16'ha00;
17'h2509:	data_out=16'h19d;
17'h250a:	data_out=16'ha00;
17'h250b:	data_out=16'h9ff;
17'h250c:	data_out=16'ha00;
17'h250d:	data_out=16'ha00;
17'h250e:	data_out=16'h68e;
17'h250f:	data_out=16'ha00;
17'h2510:	data_out=16'h9fe;
17'h2511:	data_out=16'h9f8;
17'h2512:	data_out=16'h7fd;
17'h2513:	data_out=16'ha00;
17'h2514:	data_out=16'ha00;
17'h2515:	data_out=16'ha00;
17'h2516:	data_out=16'ha00;
17'h2517:	data_out=16'ha00;
17'h2518:	data_out=16'h8306;
17'h2519:	data_out=16'h9b4;
17'h251a:	data_out=16'ha00;
17'h251b:	data_out=16'ha00;
17'h251c:	data_out=16'ha00;
17'h251d:	data_out=16'ha00;
17'h251e:	data_out=16'ha00;
17'h251f:	data_out=16'h9fe;
17'h2520:	data_out=16'h9fc;
17'h2521:	data_out=16'h6bb;
17'h2522:	data_out=16'h9ff;
17'h2523:	data_out=16'h4be;
17'h2524:	data_out=16'h4b7;
17'h2525:	data_out=16'h9fe;
17'h2526:	data_out=16'ha00;
17'h2527:	data_out=16'ha00;
17'h2528:	data_out=16'h73a;
17'h2529:	data_out=16'ha00;
17'h252a:	data_out=16'ha00;
17'h252b:	data_out=16'h8a00;
17'h252c:	data_out=16'ha00;
17'h252d:	data_out=16'h892;
17'h252e:	data_out=16'ha00;
17'h252f:	data_out=16'ha00;
17'h2530:	data_out=16'ha00;
17'h2531:	data_out=16'h841;
17'h2532:	data_out=16'ha00;
17'h2533:	data_out=16'h6c8;
17'h2534:	data_out=16'h30e;
17'h2535:	data_out=16'ha00;
17'h2536:	data_out=16'ha00;
17'h2537:	data_out=16'ha00;
17'h2538:	data_out=16'h9d0;
17'h2539:	data_out=16'h596;
17'h253a:	data_out=16'h5b;
17'h253b:	data_out=16'ha00;
17'h253c:	data_out=16'ha00;
17'h253d:	data_out=16'h9fd;
17'h253e:	data_out=16'h741;
17'h253f:	data_out=16'ha00;
17'h2540:	data_out=16'ha00;
17'h2541:	data_out=16'ha00;
17'h2542:	data_out=16'ha00;
17'h2543:	data_out=16'ha00;
17'h2544:	data_out=16'ha00;
17'h2545:	data_out=16'ha00;
17'h2546:	data_out=16'ha00;
17'h2547:	data_out=16'h680;
17'h2548:	data_out=16'ha00;
17'h2549:	data_out=16'h9fe;
17'h254a:	data_out=16'ha00;
17'h254b:	data_out=16'ha00;
17'h254c:	data_out=16'h9fe;
17'h254d:	data_out=16'h9ff;
17'h254e:	data_out=16'ha00;
17'h254f:	data_out=16'h9fc;
17'h2550:	data_out=16'ha00;
17'h2551:	data_out=16'ha00;
17'h2552:	data_out=16'h721;
17'h2553:	data_out=16'ha00;
17'h2554:	data_out=16'ha00;
17'h2555:	data_out=16'ha00;
17'h2556:	data_out=16'ha00;
17'h2557:	data_out=16'h88c;
17'h2558:	data_out=16'ha00;
17'h2559:	data_out=16'ha00;
17'h255a:	data_out=16'ha00;
17'h255b:	data_out=16'h9fd;
17'h255c:	data_out=16'ha00;
17'h255d:	data_out=16'ha00;
17'h255e:	data_out=16'ha00;
17'h255f:	data_out=16'h31f;
17'h2560:	data_out=16'ha00;
17'h2561:	data_out=16'ha00;
17'h2562:	data_out=16'ha00;
17'h2563:	data_out=16'h94d;
17'h2564:	data_out=16'h8869;
17'h2565:	data_out=16'ha00;
17'h2566:	data_out=16'h9ff;
17'h2567:	data_out=16'h808;
17'h2568:	data_out=16'h6dc;
17'h2569:	data_out=16'h91e;
17'h256a:	data_out=16'h66f;
17'h256b:	data_out=16'ha00;
17'h256c:	data_out=16'ha00;
17'h256d:	data_out=16'h934;
17'h256e:	data_out=16'h671;
17'h256f:	data_out=16'ha00;
17'h2570:	data_out=16'h683;
17'h2571:	data_out=16'h793;
17'h2572:	data_out=16'ha00;
17'h2573:	data_out=16'ha00;
17'h2574:	data_out=16'ha00;
17'h2575:	data_out=16'ha00;
17'h2576:	data_out=16'h8a00;
17'h2577:	data_out=16'ha00;
17'h2578:	data_out=16'ha00;
17'h2579:	data_out=16'ha00;
17'h257a:	data_out=16'ha00;
17'h257b:	data_out=16'h745;
17'h257c:	data_out=16'h8382;
17'h257d:	data_out=16'h888;
17'h257e:	data_out=16'h9fe;
17'h257f:	data_out=16'ha00;
17'h2580:	data_out=16'h82a7;
17'h2581:	data_out=16'ha00;
17'h2582:	data_out=16'ha00;
17'h2583:	data_out=16'ha00;
17'h2584:	data_out=16'ha00;
17'h2585:	data_out=16'ha00;
17'h2586:	data_out=16'ha00;
17'h2587:	data_out=16'h9ff;
17'h2588:	data_out=16'h9ff;
17'h2589:	data_out=16'h356;
17'h258a:	data_out=16'ha00;
17'h258b:	data_out=16'h9fc;
17'h258c:	data_out=16'ha00;
17'h258d:	data_out=16'ha00;
17'h258e:	data_out=16'h51b;
17'h258f:	data_out=16'ha00;
17'h2590:	data_out=16'h9fa;
17'h2591:	data_out=16'h9f8;
17'h2592:	data_out=16'h9a2;
17'h2593:	data_out=16'ha00;
17'h2594:	data_out=16'ha00;
17'h2595:	data_out=16'ha00;
17'h2596:	data_out=16'ha00;
17'h2597:	data_out=16'ha00;
17'h2598:	data_out=16'h8149;
17'h2599:	data_out=16'h5a8;
17'h259a:	data_out=16'ha00;
17'h259b:	data_out=16'ha00;
17'h259c:	data_out=16'ha00;
17'h259d:	data_out=16'ha00;
17'h259e:	data_out=16'ha00;
17'h259f:	data_out=16'h9fe;
17'h25a0:	data_out=16'h9fb;
17'h25a1:	data_out=16'h53e;
17'h25a2:	data_out=16'h9fc;
17'h25a3:	data_out=16'h8002;
17'h25a4:	data_out=16'h8006;
17'h25a5:	data_out=16'h9fa;
17'h25a6:	data_out=16'ha00;
17'h25a7:	data_out=16'ha00;
17'h25a8:	data_out=16'h5a8;
17'h25a9:	data_out=16'h9fd;
17'h25aa:	data_out=16'ha00;
17'h25ab:	data_out=16'h8a00;
17'h25ac:	data_out=16'ha00;
17'h25ad:	data_out=16'h955;
17'h25ae:	data_out=16'ha00;
17'h25af:	data_out=16'ha00;
17'h25b0:	data_out=16'ha00;
17'h25b1:	data_out=16'h3f1;
17'h25b2:	data_out=16'ha00;
17'h25b3:	data_out=16'ha00;
17'h25b4:	data_out=16'h42;
17'h25b5:	data_out=16'ha00;
17'h25b6:	data_out=16'ha00;
17'h25b7:	data_out=16'ha00;
17'h25b8:	data_out=16'h9da;
17'h25b9:	data_out=16'h974;
17'h25ba:	data_out=16'h411;
17'h25bb:	data_out=16'ha00;
17'h25bc:	data_out=16'ha00;
17'h25bd:	data_out=16'h9fe;
17'h25be:	data_out=16'h5af;
17'h25bf:	data_out=16'ha00;
17'h25c0:	data_out=16'ha00;
17'h25c1:	data_out=16'ha00;
17'h25c2:	data_out=16'ha00;
17'h25c3:	data_out=16'ha00;
17'h25c4:	data_out=16'ha00;
17'h25c5:	data_out=16'ha00;
17'h25c6:	data_out=16'h9fd;
17'h25c7:	data_out=16'h7d7;
17'h25c8:	data_out=16'h9ff;
17'h25c9:	data_out=16'h9fa;
17'h25ca:	data_out=16'h9fd;
17'h25cb:	data_out=16'h9ff;
17'h25cc:	data_out=16'h9fb;
17'h25cd:	data_out=16'h9fb;
17'h25ce:	data_out=16'h9fd;
17'h25cf:	data_out=16'h9fa;
17'h25d0:	data_out=16'ha00;
17'h25d1:	data_out=16'ha00;
17'h25d2:	data_out=16'h197;
17'h25d3:	data_out=16'ha00;
17'h25d4:	data_out=16'h9ff;
17'h25d5:	data_out=16'ha00;
17'h25d6:	data_out=16'h9ff;
17'h25d7:	data_out=16'h812;
17'h25d8:	data_out=16'ha00;
17'h25d9:	data_out=16'ha00;
17'h25da:	data_out=16'ha00;
17'h25db:	data_out=16'h9fa;
17'h25dc:	data_out=16'ha00;
17'h25dd:	data_out=16'ha00;
17'h25de:	data_out=16'ha00;
17'h25df:	data_out=16'h301;
17'h25e0:	data_out=16'ha00;
17'h25e1:	data_out=16'ha00;
17'h25e2:	data_out=16'ha00;
17'h25e3:	data_out=16'ha00;
17'h25e4:	data_out=16'h8703;
17'h25e5:	data_out=16'ha00;
17'h25e6:	data_out=16'h681;
17'h25e7:	data_out=16'h8f2;
17'h25e8:	data_out=16'h558;
17'h25e9:	data_out=16'h880;
17'h25ea:	data_out=16'h502;
17'h25eb:	data_out=16'ha00;
17'h25ec:	data_out=16'ha00;
17'h25ed:	data_out=16'ha00;
17'h25ee:	data_out=16'h503;
17'h25ef:	data_out=16'ha00;
17'h25f0:	data_out=16'h511;
17'h25f1:	data_out=16'ha00;
17'h25f2:	data_out=16'ha00;
17'h25f3:	data_out=16'ha00;
17'h25f4:	data_out=16'ha00;
17'h25f5:	data_out=16'ha00;
17'h25f6:	data_out=16'h8a00;
17'h25f7:	data_out=16'h9ff;
17'h25f8:	data_out=16'ha00;
17'h25f9:	data_out=16'h9fe;
17'h25fa:	data_out=16'ha00;
17'h25fb:	data_out=16'h5b3;
17'h25fc:	data_out=16'h8236;
17'h25fd:	data_out=16'h915;
17'h25fe:	data_out=16'h9fe;
17'h25ff:	data_out=16'ha00;
17'h2600:	data_out=16'h8605;
17'h2601:	data_out=16'h80a;
17'h2602:	data_out=16'h9fd;
17'h2603:	data_out=16'ha00;
17'h2604:	data_out=16'ha00;
17'h2605:	data_out=16'ha00;
17'h2606:	data_out=16'ha00;
17'h2607:	data_out=16'ha00;
17'h2608:	data_out=16'h9e5;
17'h2609:	data_out=16'h4a7;
17'h260a:	data_out=16'h658;
17'h260b:	data_out=16'h9ff;
17'h260c:	data_out=16'ha00;
17'h260d:	data_out=16'ha00;
17'h260e:	data_out=16'h379;
17'h260f:	data_out=16'ha00;
17'h2610:	data_out=16'ha00;
17'h2611:	data_out=16'h9f0;
17'h2612:	data_out=16'h9bd;
17'h2613:	data_out=16'ha00;
17'h2614:	data_out=16'h968;
17'h2615:	data_out=16'h5e7;
17'h2616:	data_out=16'ha00;
17'h2617:	data_out=16'ha00;
17'h2618:	data_out=16'h8142;
17'h2619:	data_out=16'h852;
17'h261a:	data_out=16'ha00;
17'h261b:	data_out=16'ha00;
17'h261c:	data_out=16'ha00;
17'h261d:	data_out=16'h9f7;
17'h261e:	data_out=16'ha00;
17'h261f:	data_out=16'h9fe;
17'h2620:	data_out=16'h993;
17'h2621:	data_out=16'h38b;
17'h2622:	data_out=16'ha00;
17'h2623:	data_out=16'h8019;
17'h2624:	data_out=16'h801c;
17'h2625:	data_out=16'h9ff;
17'h2626:	data_out=16'h80e;
17'h2627:	data_out=16'h9fe;
17'h2628:	data_out=16'h3cb;
17'h2629:	data_out=16'h9ea;
17'h262a:	data_out=16'ha00;
17'h262b:	data_out=16'h8881;
17'h262c:	data_out=16'ha00;
17'h262d:	data_out=16'h96c;
17'h262e:	data_out=16'ha00;
17'h262f:	data_out=16'ha00;
17'h2630:	data_out=16'ha00;
17'h2631:	data_out=16'h818e;
17'h2632:	data_out=16'ha00;
17'h2633:	data_out=16'h6ae;
17'h2634:	data_out=16'h81ca;
17'h2635:	data_out=16'ha00;
17'h2636:	data_out=16'h9fe;
17'h2637:	data_out=16'h9ff;
17'h2638:	data_out=16'h7ba;
17'h2639:	data_out=16'h5da;
17'h263a:	data_out=16'h5e7;
17'h263b:	data_out=16'ha00;
17'h263c:	data_out=16'ha00;
17'h263d:	data_out=16'h9f6;
17'h263e:	data_out=16'h3d0;
17'h263f:	data_out=16'ha00;
17'h2640:	data_out=16'ha00;
17'h2641:	data_out=16'ha00;
17'h2642:	data_out=16'ha00;
17'h2643:	data_out=16'ha00;
17'h2644:	data_out=16'h9f8;
17'h2645:	data_out=16'h68d;
17'h2646:	data_out=16'h901;
17'h2647:	data_out=16'h90c;
17'h2648:	data_out=16'ha00;
17'h2649:	data_out=16'h9ff;
17'h264a:	data_out=16'ha00;
17'h264b:	data_out=16'ha00;
17'h264c:	data_out=16'h9ff;
17'h264d:	data_out=16'ha00;
17'h264e:	data_out=16'h9f0;
17'h264f:	data_out=16'h9ff;
17'h2650:	data_out=16'ha00;
17'h2651:	data_out=16'h9f9;
17'h2652:	data_out=16'h9f;
17'h2653:	data_out=16'ha00;
17'h2654:	data_out=16'h9fd;
17'h2655:	data_out=16'ha00;
17'h2656:	data_out=16'h9f6;
17'h2657:	data_out=16'h8da;
17'h2658:	data_out=16'h9fb;
17'h2659:	data_out=16'ha00;
17'h265a:	data_out=16'ha00;
17'h265b:	data_out=16'h97c;
17'h265c:	data_out=16'ha00;
17'h265d:	data_out=16'ha00;
17'h265e:	data_out=16'ha00;
17'h265f:	data_out=16'h216;
17'h2660:	data_out=16'h7e7;
17'h2661:	data_out=16'ha00;
17'h2662:	data_out=16'ha00;
17'h2663:	data_out=16'h7cc;
17'h2664:	data_out=16'h8511;
17'h2665:	data_out=16'ha00;
17'h2666:	data_out=16'h6fe;
17'h2667:	data_out=16'h9f3;
17'h2668:	data_out=16'h39a;
17'h2669:	data_out=16'h76b;
17'h266a:	data_out=16'h36e;
17'h266b:	data_out=16'ha00;
17'h266c:	data_out=16'h992;
17'h266d:	data_out=16'h7c1;
17'h266e:	data_out=16'h36f;
17'h266f:	data_out=16'ha00;
17'h2670:	data_out=16'h375;
17'h2671:	data_out=16'h5d4;
17'h2672:	data_out=16'ha00;
17'h2673:	data_out=16'ha00;
17'h2674:	data_out=16'ha00;
17'h2675:	data_out=16'ha00;
17'h2676:	data_out=16'h884a;
17'h2677:	data_out=16'ha00;
17'h2678:	data_out=16'ha00;
17'h2679:	data_out=16'h9f4;
17'h267a:	data_out=16'h963;
17'h267b:	data_out=16'h3d2;
17'h267c:	data_out=16'h8197;
17'h267d:	data_out=16'h9de;
17'h267e:	data_out=16'h9ff;
17'h267f:	data_out=16'ha00;
17'h2680:	data_out=16'h8992;
17'h2681:	data_out=16'h8025;
17'h2682:	data_out=16'h7df;
17'h2683:	data_out=16'ha00;
17'h2684:	data_out=16'h9ff;
17'h2685:	data_out=16'ha00;
17'h2686:	data_out=16'h96f;
17'h2687:	data_out=16'h9af;
17'h2688:	data_out=16'h219;
17'h2689:	data_out=16'h27d;
17'h268a:	data_out=16'h8100;
17'h268b:	data_out=16'h9ed;
17'h268c:	data_out=16'ha00;
17'h268d:	data_out=16'h933;
17'h268e:	data_out=16'h1d8;
17'h268f:	data_out=16'h82b;
17'h2690:	data_out=16'ha00;
17'h2691:	data_out=16'h9f4;
17'h2692:	data_out=16'h7f6;
17'h2693:	data_out=16'h9ff;
17'h2694:	data_out=16'h158;
17'h2695:	data_out=16'h223;
17'h2696:	data_out=16'h9b3;
17'h2697:	data_out=16'h5d4;
17'h2698:	data_out=16'h8142;
17'h2699:	data_out=16'h83f;
17'h269a:	data_out=16'ha00;
17'h269b:	data_out=16'h9fb;
17'h269c:	data_out=16'h790;
17'h269d:	data_out=16'h253;
17'h269e:	data_out=16'h428;
17'h269f:	data_out=16'h6ea;
17'h26a0:	data_out=16'h1fd;
17'h26a1:	data_out=16'h1ee;
17'h26a2:	data_out=16'ha00;
17'h26a3:	data_out=16'hb9;
17'h26a4:	data_out=16'hb7;
17'h26a5:	data_out=16'ha00;
17'h26a6:	data_out=16'h8048;
17'h26a7:	data_out=16'h2a7;
17'h26a8:	data_out=16'h220;
17'h26a9:	data_out=16'h6f9;
17'h26aa:	data_out=16'h9fb;
17'h26ab:	data_out=16'h8945;
17'h26ac:	data_out=16'h819;
17'h26ad:	data_out=16'h966;
17'h26ae:	data_out=16'h9fd;
17'h26af:	data_out=16'ha00;
17'h26b0:	data_out=16'ha00;
17'h26b1:	data_out=16'h8641;
17'h26b2:	data_out=16'ha00;
17'h26b3:	data_out=16'h8017;
17'h26b4:	data_out=16'h8569;
17'h26b5:	data_out=16'h9f6;
17'h26b6:	data_out=16'h31b;
17'h26b7:	data_out=16'h881;
17'h26b8:	data_out=16'h80cd;
17'h26b9:	data_out=16'h808c;
17'h26ba:	data_out=16'h35e;
17'h26bb:	data_out=16'h53b;
17'h26bc:	data_out=16'h9fa;
17'h26bd:	data_out=16'h342;
17'h26be:	data_out=16'h222;
17'h26bf:	data_out=16'ha00;
17'h26c0:	data_out=16'ha00;
17'h26c1:	data_out=16'h95f;
17'h26c2:	data_out=16'h9fe;
17'h26c3:	data_out=16'ha00;
17'h26c4:	data_out=16'h263;
17'h26c5:	data_out=16'h274;
17'h26c6:	data_out=16'h5b0;
17'h26c7:	data_out=16'h648;
17'h26c8:	data_out=16'ha00;
17'h26c9:	data_out=16'ha00;
17'h26ca:	data_out=16'ha00;
17'h26cb:	data_out=16'h9fe;
17'h26cc:	data_out=16'ha00;
17'h26cd:	data_out=16'ha00;
17'h26ce:	data_out=16'h9b9;
17'h26cf:	data_out=16'h841;
17'h26d0:	data_out=16'ha00;
17'h26d1:	data_out=16'h90f;
17'h26d2:	data_out=16'h11a;
17'h26d3:	data_out=16'h9fd;
17'h26d4:	data_out=16'h840;
17'h26d5:	data_out=16'h73e;
17'h26d6:	data_out=16'h6e8;
17'h26d7:	data_out=16'h784;
17'h26d8:	data_out=16'h4fa;
17'h26d9:	data_out=16'ha00;
17'h26da:	data_out=16'h9ec;
17'h26db:	data_out=16'h80a9;
17'h26dc:	data_out=16'h5c2;
17'h26dd:	data_out=16'ha00;
17'h26de:	data_out=16'ha00;
17'h26df:	data_out=16'he2;
17'h26e0:	data_out=16'h801e;
17'h26e1:	data_out=16'h4e1;
17'h26e2:	data_out=16'h819;
17'h26e3:	data_out=16'h90;
17'h26e4:	data_out=16'h867b;
17'h26e5:	data_out=16'ha00;
17'h26e6:	data_out=16'h73d;
17'h26e7:	data_out=16'h8dc;
17'h26e8:	data_out=16'h1fd;
17'h26e9:	data_out=16'h264;
17'h26ea:	data_out=16'h1ca;
17'h26eb:	data_out=16'ha00;
17'h26ec:	data_out=16'he6;
17'h26ed:	data_out=16'h89;
17'h26ee:	data_out=16'h1cb;
17'h26ef:	data_out=16'ha00;
17'h26f0:	data_out=16'h1d3;
17'h26f1:	data_out=16'h7f;
17'h26f2:	data_out=16'ha00;
17'h26f3:	data_out=16'ha00;
17'h26f4:	data_out=16'ha00;
17'h26f5:	data_out=16'ha00;
17'h26f6:	data_out=16'h89bc;
17'h26f7:	data_out=16'ha00;
17'h26f8:	data_out=16'ha00;
17'h26f9:	data_out=16'h9be;
17'h26fa:	data_out=16'h16e;
17'h26fb:	data_out=16'h223;
17'h26fc:	data_out=16'h813c;
17'h26fd:	data_out=16'h9dd;
17'h26fe:	data_out=16'h6b1;
17'h26ff:	data_out=16'ha00;
17'h2700:	data_out=16'h8520;
17'h2701:	data_out=16'h800a;
17'h2702:	data_out=16'h4e5;
17'h2703:	data_out=16'h74a;
17'h2704:	data_out=16'h9fd;
17'h2705:	data_out=16'h9ab;
17'h2706:	data_out=16'h4f1;
17'h2707:	data_out=16'h4d8;
17'h2708:	data_out=16'he9;
17'h2709:	data_out=16'h8040;
17'h270a:	data_out=16'h8088;
17'h270b:	data_out=16'h5a3;
17'h270c:	data_out=16'ha00;
17'h270d:	data_out=16'h4d5;
17'h270e:	data_out=16'h167;
17'h270f:	data_out=16'h45a;
17'h2710:	data_out=16'h4b9;
17'h2711:	data_out=16'h7ac;
17'h2712:	data_out=16'h385;
17'h2713:	data_out=16'h96c;
17'h2714:	data_out=16'h41;
17'h2715:	data_out=16'h85;
17'h2716:	data_out=16'h55e;
17'h2717:	data_out=16'h2ab;
17'h2718:	data_out=16'h8062;
17'h2719:	data_out=16'h4c0;
17'h271a:	data_out=16'h9ff;
17'h271b:	data_out=16'h5c2;
17'h271c:	data_out=16'h34f;
17'h271d:	data_out=16'h10f;
17'h271e:	data_out=16'h1b7;
17'h271f:	data_out=16'h3b2;
17'h2720:	data_out=16'hae;
17'h2721:	data_out=16'h170;
17'h2722:	data_out=16'h660;
17'h2723:	data_out=16'h8090;
17'h2724:	data_out=16'h80a8;
17'h2725:	data_out=16'h655;
17'h2726:	data_out=16'h8164;
17'h2727:	data_out=16'h116;
17'h2728:	data_out=16'h184;
17'h2729:	data_out=16'h39e;
17'h272a:	data_out=16'h512;
17'h272b:	data_out=16'h8621;
17'h272c:	data_out=16'h48e;
17'h272d:	data_out=16'h67a;
17'h272e:	data_out=16'h614;
17'h272f:	data_out=16'h849;
17'h2730:	data_out=16'ha00;
17'h2731:	data_out=16'h8327;
17'h2732:	data_out=16'ha00;
17'h2733:	data_out=16'h80a0;
17'h2734:	data_out=16'h82c1;
17'h2735:	data_out=16'h9fc;
17'h2736:	data_out=16'h23f;
17'h2737:	data_out=16'h52e;
17'h2738:	data_out=16'h824c;
17'h2739:	data_out=16'h80d8;
17'h273a:	data_out=16'h11f;
17'h273b:	data_out=16'h2eb;
17'h273c:	data_out=16'h7a8;
17'h273d:	data_out=16'hb2;
17'h273e:	data_out=16'h185;
17'h273f:	data_out=16'h9a6;
17'h2740:	data_out=16'ha00;
17'h2741:	data_out=16'h622;
17'h2742:	data_out=16'h9fd;
17'h2743:	data_out=16'h598;
17'h2744:	data_out=16'h1dd;
17'h2745:	data_out=16'h802c;
17'h2746:	data_out=16'h3a0;
17'h2747:	data_out=16'h3db;
17'h2748:	data_out=16'h65b;
17'h2749:	data_out=16'h641;
17'h274a:	data_out=16'h79a;
17'h274b:	data_out=16'h9fe;
17'h274c:	data_out=16'h65f;
17'h274d:	data_out=16'h647;
17'h274e:	data_out=16'h6df;
17'h274f:	data_out=16'h4fa;
17'h2750:	data_out=16'h91b;
17'h2751:	data_out=16'h394;
17'h2752:	data_out=16'h804f;
17'h2753:	data_out=16'h591;
17'h2754:	data_out=16'h44b;
17'h2755:	data_out=16'h487;
17'h2756:	data_out=16'h44a;
17'h2757:	data_out=16'h418;
17'h2758:	data_out=16'h36d;
17'h2759:	data_out=16'h9ff;
17'h275a:	data_out=16'h4d4;
17'h275b:	data_out=16'h8036;
17'h275c:	data_out=16'h3df;
17'h275d:	data_out=16'h80e;
17'h275e:	data_out=16'h91d;
17'h275f:	data_out=16'hc2;
17'h2760:	data_out=16'h80c5;
17'h2761:	data_out=16'h25d;
17'h2762:	data_out=16'h58b;
17'h2763:	data_out=16'h803f;
17'h2764:	data_out=16'h84b6;
17'h2765:	data_out=16'h8b1;
17'h2766:	data_out=16'h4f0;
17'h2767:	data_out=16'h4e4;
17'h2768:	data_out=16'h175;
17'h2769:	data_out=16'h1f5;
17'h276a:	data_out=16'h161;
17'h276b:	data_out=16'h9fe;
17'h276c:	data_out=16'h122;
17'h276d:	data_out=16'h8046;
17'h276e:	data_out=16'h161;
17'h276f:	data_out=16'ha00;
17'h2770:	data_out=16'h165;
17'h2771:	data_out=16'h78;
17'h2772:	data_out=16'h9da;
17'h2773:	data_out=16'h984;
17'h2774:	data_out=16'ha00;
17'h2775:	data_out=16'h6d1;
17'h2776:	data_out=16'h8729;
17'h2777:	data_out=16'h99c;
17'h2778:	data_out=16'h6dc;
17'h2779:	data_out=16'h5bf;
17'h277a:	data_out=16'h4c;
17'h277b:	data_out=16'h186;
17'h277c:	data_out=16'h8052;
17'h277d:	data_out=16'h5d3;
17'h277e:	data_out=16'h1dd;
17'h277f:	data_out=16'h6c5;
17'h2780:	data_out=16'h841d;
17'h2781:	data_out=16'h82c1;
17'h2782:	data_out=16'h8162;
17'h2783:	data_out=16'h299;
17'h2784:	data_out=16'h6ac;
17'h2785:	data_out=16'h494;
17'h2786:	data_out=16'hc5;
17'h2787:	data_out=16'h1e1;
17'h2788:	data_out=16'h83c9;
17'h2789:	data_out=16'h80ae;
17'h278a:	data_out=16'h81ed;
17'h278b:	data_out=16'h8023;
17'h278c:	data_out=16'h80f;
17'h278d:	data_out=16'hd5;
17'h278e:	data_out=16'h22;
17'h278f:	data_out=16'h8224;
17'h2790:	data_out=16'hb6;
17'h2791:	data_out=16'h514;
17'h2792:	data_out=16'h8136;
17'h2793:	data_out=16'h330;
17'h2794:	data_out=16'h8273;
17'h2795:	data_out=16'h8058;
17'h2796:	data_out=16'h5e;
17'h2797:	data_out=16'h8170;
17'h2798:	data_out=16'h80ee;
17'h2799:	data_out=16'h51c;
17'h279a:	data_out=16'h798;
17'h279b:	data_out=16'h16;
17'h279c:	data_out=16'h8146;
17'h279d:	data_out=16'h81ab;
17'h279e:	data_out=16'h830b;
17'h279f:	data_out=16'h4a;
17'h27a0:	data_out=16'h8018;
17'h27a1:	data_out=16'h40;
17'h27a2:	data_out=16'h3c3;
17'h27a3:	data_out=16'h814b;
17'h27a4:	data_out=16'h814b;
17'h27a5:	data_out=16'h465;
17'h27a6:	data_out=16'h8460;
17'h27a7:	data_out=16'h81e5;
17'h27a8:	data_out=16'h5a;
17'h27a9:	data_out=16'h8037;
17'h27aa:	data_out=16'h8273;
17'h27ab:	data_out=16'h8379;
17'h27ac:	data_out=16'h126;
17'h27ad:	data_out=16'h393;
17'h27ae:	data_out=16'h8096;
17'h27af:	data_out=16'h26a;
17'h27b0:	data_out=16'h74c;
17'h27b1:	data_out=16'h827b;
17'h27b2:	data_out=16'h779;
17'h27b3:	data_out=16'h82ea;
17'h27b4:	data_out=16'h80f2;
17'h27b5:	data_out=16'h663;
17'h27b6:	data_out=16'h82b3;
17'h27b7:	data_out=16'h80c7;
17'h27b8:	data_out=16'h833a;
17'h27b9:	data_out=16'h8490;
17'h27ba:	data_out=16'h808d;
17'h27bb:	data_out=16'hef;
17'h27bc:	data_out=16'h808a;
17'h27bd:	data_out=16'h8151;
17'h27be:	data_out=16'h55;
17'h27bf:	data_out=16'h491;
17'h27c0:	data_out=16'h551;
17'h27c1:	data_out=16'ha4;
17'h27c2:	data_out=16'h6c5;
17'h27c3:	data_out=16'h2b4;
17'h27c4:	data_out=16'h13;
17'h27c5:	data_out=16'h8163;
17'h27c6:	data_out=16'h807f;
17'h27c7:	data_out=16'hdc;
17'h27c8:	data_out=16'hfd;
17'h27c9:	data_out=16'h468;
17'h27ca:	data_out=16'h42f;
17'h27cb:	data_out=16'h973;
17'h27cc:	data_out=16'h3f7;
17'h27cd:	data_out=16'h38a;
17'h27ce:	data_out=16'h8069;
17'h27cf:	data_out=16'h334;
17'h27d0:	data_out=16'h353;
17'h27d1:	data_out=16'h8182;
17'h27d2:	data_out=16'h8131;
17'h27d3:	data_out=16'h3a;
17'h27d4:	data_out=16'h114;
17'h27d5:	data_out=16'h81f9;
17'h27d6:	data_out=16'h7b;
17'h27d7:	data_out=16'h37;
17'h27d8:	data_out=16'h827d;
17'h27d9:	data_out=16'h44b;
17'h27da:	data_out=16'h8146;
17'h27db:	data_out=16'h8376;
17'h27dc:	data_out=16'h192;
17'h27dd:	data_out=16'h28f;
17'h27de:	data_out=16'h3f3;
17'h27df:	data_out=16'h31;
17'h27e0:	data_out=16'h82fc;
17'h27e1:	data_out=16'h8074;
17'h27e2:	data_out=16'h806a;
17'h27e3:	data_out=16'h82ad;
17'h27e4:	data_out=16'h8337;
17'h27e5:	data_out=16'h63b;
17'h27e6:	data_out=16'h532;
17'h27e7:	data_out=16'h50;
17'h27e8:	data_out=16'h4b;
17'h27e9:	data_out=16'h82b6;
17'h27ea:	data_out=16'h1c;
17'h27eb:	data_out=16'h5be;
17'h27ec:	data_out=16'h81f7;
17'h27ed:	data_out=16'h82d7;
17'h27ee:	data_out=16'h12;
17'h27ef:	data_out=16'h7a1;
17'h27f0:	data_out=16'h26;
17'h27f1:	data_out=16'h837e;
17'h27f2:	data_out=16'h3b9;
17'h27f3:	data_out=16'h433;
17'h27f4:	data_out=16'h750;
17'h27f5:	data_out=16'h9;
17'h27f6:	data_out=16'h846c;
17'h27f7:	data_out=16'h4a1;
17'h27f8:	data_out=16'h344;
17'h27f9:	data_out=16'h8265;
17'h27fa:	data_out=16'h827f;
17'h27fb:	data_out=16'h55;
17'h27fc:	data_out=16'h816a;
17'h27fd:	data_out=16'h12c;
17'h27fe:	data_out=16'h808f;
17'h27ff:	data_out=16'h33a;
17'h2800:	data_out=16'h8040;
17'h2801:	data_out=16'h80d1;
17'h2802:	data_out=16'h835a;
17'h2803:	data_out=16'h87;
17'h2804:	data_out=16'h384;
17'h2805:	data_out=16'h1ea;
17'h2806:	data_out=16'h803f;
17'h2807:	data_out=16'h98;
17'h2808:	data_out=16'h8318;
17'h2809:	data_out=16'h1bd;
17'h280a:	data_out=16'h810c;
17'h280b:	data_out=16'h8113;
17'h280c:	data_out=16'h329;
17'h280d:	data_out=16'h8019;
17'h280e:	data_out=16'h8065;
17'h280f:	data_out=16'h823c;
17'h2810:	data_out=16'h8052;
17'h2811:	data_out=16'h369;
17'h2812:	data_out=16'h8293;
17'h2813:	data_out=16'h168;
17'h2814:	data_out=16'h820c;
17'h2815:	data_out=16'hb9;
17'h2816:	data_out=16'h16;
17'h2817:	data_out=16'h8202;
17'h2818:	data_out=16'h80d5;
17'h2819:	data_out=16'h4a4;
17'h281a:	data_out=16'h47c;
17'h281b:	data_out=16'h804f;
17'h281c:	data_out=16'h9d;
17'h281d:	data_out=16'h80dd;
17'h281e:	data_out=16'h81c9;
17'h281f:	data_out=16'h8097;
17'h2820:	data_out=16'h1d6;
17'h2821:	data_out=16'h8057;
17'h2822:	data_out=16'h2fa;
17'h2823:	data_out=16'h81f8;
17'h2824:	data_out=16'h81f8;
17'h2825:	data_out=16'h1f4;
17'h2826:	data_out=16'h8257;
17'h2827:	data_out=16'h80ab;
17'h2828:	data_out=16'h8041;
17'h2829:	data_out=16'h80cb;
17'h282a:	data_out=16'h8377;
17'h282b:	data_out=16'h280;
17'h282c:	data_out=16'h9;
17'h282d:	data_out=16'h1f1;
17'h282e:	data_out=16'h8301;
17'h282f:	data_out=16'h1e2;
17'h2830:	data_out=16'h3ee;
17'h2831:	data_out=16'he1;
17'h2832:	data_out=16'h414;
17'h2833:	data_out=16'h819c;
17'h2834:	data_out=16'h21d;
17'h2835:	data_out=16'h340;
17'h2836:	data_out=16'h83db;
17'h2837:	data_out=16'h8308;
17'h2838:	data_out=16'hff;
17'h2839:	data_out=16'h8147;
17'h283a:	data_out=16'h80ca;
17'h283b:	data_out=16'h91;
17'h283c:	data_out=16'h8323;
17'h283d:	data_out=16'h292;
17'h283e:	data_out=16'h8048;
17'h283f:	data_out=16'h2bb;
17'h2840:	data_out=16'h1c4;
17'h2841:	data_out=16'h81db;
17'h2842:	data_out=16'h1bb;
17'h2843:	data_out=16'h135;
17'h2844:	data_out=16'h105;
17'h2845:	data_out=16'hb5;
17'h2846:	data_out=16'h8185;
17'h2847:	data_out=16'h806d;
17'h2848:	data_out=16'h80ff;
17'h2849:	data_out=16'h20c;
17'h284a:	data_out=16'hcb;
17'h284b:	data_out=16'h254;
17'h284c:	data_out=16'h96;
17'h284d:	data_out=16'h3a7;
17'h284e:	data_out=16'h8227;
17'h284f:	data_out=16'hc2;
17'h2850:	data_out=16'h118;
17'h2851:	data_out=16'h8169;
17'h2852:	data_out=16'h81eb;
17'h2853:	data_out=16'h2e;
17'h2854:	data_out=16'h107;
17'h2855:	data_out=16'h8428;
17'h2856:	data_out=16'h8103;
17'h2857:	data_out=16'h80ec;
17'h2858:	data_out=16'h8491;
17'h2859:	data_out=16'h9c;
17'h285a:	data_out=16'h8260;
17'h285b:	data_out=16'h826a;
17'h285c:	data_out=16'h65;
17'h285d:	data_out=16'h8003;
17'h285e:	data_out=16'h22d;
17'h285f:	data_out=16'h803d;
17'h2860:	data_out=16'h8283;
17'h2861:	data_out=16'h5f;
17'h2862:	data_out=16'h822f;
17'h2863:	data_out=16'h8165;
17'h2864:	data_out=16'h144;
17'h2865:	data_out=16'h3b8;
17'h2866:	data_out=16'h49a;
17'h2867:	data_out=16'h810a;
17'h2868:	data_out=16'h8052;
17'h2869:	data_out=16'h8475;
17'h286a:	data_out=16'h8064;
17'h286b:	data_out=16'h3e9;
17'h286c:	data_out=16'h82ac;
17'h286d:	data_out=16'h8184;
17'h286e:	data_out=16'h8066;
17'h286f:	data_out=16'h36a;
17'h2870:	data_out=16'h8064;
17'h2871:	data_out=16'h8415;
17'h2872:	data_out=16'h11f;
17'h2873:	data_out=16'h256;
17'h2874:	data_out=16'h3eb;
17'h2875:	data_out=16'h81a0;
17'h2876:	data_out=16'h125;
17'h2877:	data_out=16'h24e;
17'h2878:	data_out=16'h27b;
17'h2879:	data_out=16'h84a2;
17'h287a:	data_out=16'h8204;
17'h287b:	data_out=16'h8047;
17'h287c:	data_out=16'h814b;
17'h287d:	data_out=16'h26;
17'h287e:	data_out=16'h1bb;
17'h287f:	data_out=16'hde;
17'h2880:	data_out=16'h11b;
17'h2881:	data_out=16'h69;
17'h2882:	data_out=16'h81c6;
17'h2883:	data_out=16'h8002;
17'h2884:	data_out=16'h121;
17'h2885:	data_out=16'h9d;
17'h2886:	data_out=16'h8065;
17'h2887:	data_out=16'h800c;
17'h2888:	data_out=16'h80d0;
17'h2889:	data_out=16'h139;
17'h288a:	data_out=16'he;
17'h288b:	data_out=16'h80b2;
17'h288c:	data_out=16'h90;
17'h288d:	data_out=16'h8040;
17'h288e:	data_out=16'h8033;
17'h288f:	data_out=16'h8108;
17'h2890:	data_out=16'h804d;
17'h2891:	data_out=16'h170;
17'h2892:	data_out=16'h81a2;
17'h2893:	data_out=16'h83;
17'h2894:	data_out=16'h80da;
17'h2895:	data_out=16'hd1;
17'h2896:	data_out=16'h88;
17'h2897:	data_out=16'h80fc;
17'h2898:	data_out=16'h806f;
17'h2899:	data_out=16'h25f;
17'h289a:	data_out=16'h155;
17'h289b:	data_out=16'h8017;
17'h289c:	data_out=16'h103;
17'h289d:	data_out=16'h2c;
17'h289e:	data_out=16'h808f;
17'h289f:	data_out=16'h8072;
17'h28a0:	data_out=16'h18d;
17'h28a1:	data_out=16'h8039;
17'h28a2:	data_out=16'h11b;
17'h28a3:	data_out=16'h810e;
17'h28a4:	data_out=16'h810c;
17'h28a5:	data_out=16'h3c;
17'h28a6:	data_out=16'h8073;
17'h28a7:	data_out=16'h4a;
17'h28a8:	data_out=16'h8031;
17'h28a9:	data_out=16'h80ac;
17'h28aa:	data_out=16'h81cf;
17'h28ab:	data_out=16'h294;
17'h28ac:	data_out=16'h801d;
17'h28ad:	data_out=16'h4f;
17'h28ae:	data_out=16'h81b7;
17'h28af:	data_out=16'h122;
17'h28b0:	data_out=16'h12e;
17'h28b1:	data_out=16'h171;
17'h28b2:	data_out=16'h138;
17'h28b3:	data_out=16'h8073;
17'h28b4:	data_out=16'h19a;
17'h28b5:	data_out=16'hd8;
17'h28b6:	data_out=16'h81a9;
17'h28b7:	data_out=16'h81a9;
17'h28b8:	data_out=16'h1de;
17'h28b9:	data_out=16'h11;
17'h28ba:	data_out=16'h8082;
17'h28bb:	data_out=16'ha6;
17'h28bc:	data_out=16'h8190;
17'h28bd:	data_out=16'h25f;
17'h28be:	data_out=16'h803d;
17'h28bf:	data_out=16'hda;
17'h28c0:	data_out=16'h9;
17'h28c1:	data_out=16'h80f4;
17'h28c2:	data_out=16'h8090;
17'h28c3:	data_out=16'h17;
17'h28c4:	data_out=16'h84;
17'h28c5:	data_out=16'hf8;
17'h28c6:	data_out=16'h8099;
17'h28c7:	data_out=16'h80a0;
17'h28c8:	data_out=16'h80ef;
17'h28c9:	data_out=16'h54;
17'h28ca:	data_out=16'h8087;
17'h28cb:	data_out=16'h80ca;
17'h28cc:	data_out=16'h80c8;
17'h28cd:	data_out=16'h1a0;
17'h28ce:	data_out=16'h8127;
17'h28cf:	data_out=16'h80ad;
17'h28d0:	data_out=16'h8001;
17'h28d1:	data_out=16'h803d;
17'h28d2:	data_out=16'h80d5;
17'h28d3:	data_out=16'h71;
17'h28d4:	data_out=16'hdd;
17'h28d5:	data_out=16'h81fc;
17'h28d6:	data_out=16'h80c4;
17'h28d7:	data_out=16'h8091;
17'h28d8:	data_out=16'h822e;
17'h28d9:	data_out=16'h805d;
17'h28da:	data_out=16'h8122;
17'h28db:	data_out=16'h8064;
17'h28dc:	data_out=16'h48;
17'h28dd:	data_out=16'h8039;
17'h28de:	data_out=16'hd8;
17'h28df:	data_out=16'h8035;
17'h28e0:	data_out=16'h8110;
17'h28e1:	data_out=16'h9c;
17'h28e2:	data_out=16'h8154;
17'h28e3:	data_out=16'h808b;
17'h28e4:	data_out=16'h172;
17'h28e5:	data_out=16'h130;
17'h28e6:	data_out=16'h1d0;
17'h28e7:	data_out=16'h80c4;
17'h28e8:	data_out=16'h8034;
17'h28e9:	data_out=16'h8202;
17'h28ea:	data_out=16'h8041;
17'h28eb:	data_out=16'h1d1;
17'h28ec:	data_out=16'h80f0;
17'h28ed:	data_out=16'h8074;
17'h28ee:	data_out=16'h803f;
17'h28ef:	data_out=16'hf7;
17'h28f0:	data_out=16'h8041;
17'h28f1:	data_out=16'h8219;
17'h28f2:	data_out=16'h3e;
17'h28f3:	data_out=16'hff;
17'h28f4:	data_out=16'h131;
17'h28f5:	data_out=16'h80ca;
17'h28f6:	data_out=16'h1a2;
17'h28f7:	data_out=16'h21;
17'h28f8:	data_out=16'hf3;
17'h28f9:	data_out=16'h826f;
17'h28fa:	data_out=16'h80d7;
17'h28fb:	data_out=16'h803b;
17'h28fc:	data_out=16'h8096;
17'h28fd:	data_out=16'h8033;
17'h28fe:	data_out=16'h15c;
17'h28ff:	data_out=16'h8021;
17'h2900:	data_out=16'h8001;
17'h2901:	data_out=16'h0;
17'h2902:	data_out=16'h8004;
17'h2903:	data_out=16'h2;
17'h2904:	data_out=16'h8005;
17'h2905:	data_out=16'h4;
17'h2906:	data_out=16'h5;
17'h2907:	data_out=16'h8009;
17'h2908:	data_out=16'h7;
17'h2909:	data_out=16'h8007;
17'h290a:	data_out=16'h8006;
17'h290b:	data_out=16'h6;
17'h290c:	data_out=16'h8001;
17'h290d:	data_out=16'h3;
17'h290e:	data_out=16'h7;
17'h290f:	data_out=16'h5;
17'h2910:	data_out=16'h8003;
17'h2911:	data_out=16'h8002;
17'h2912:	data_out=16'h7;
17'h2913:	data_out=16'h7;
17'h2914:	data_out=16'h8008;
17'h2915:	data_out=16'h8;
17'h2916:	data_out=16'h8005;
17'h2917:	data_out=16'h8005;
17'h2918:	data_out=16'h8005;
17'h2919:	data_out=16'h3;
17'h291a:	data_out=16'h0;
17'h291b:	data_out=16'h7;
17'h291c:	data_out=16'h8001;
17'h291d:	data_out=16'h8008;
17'h291e:	data_out=16'h5;
17'h291f:	data_out=16'h8;
17'h2920:	data_out=16'h1;
17'h2921:	data_out=16'h8008;
17'h2922:	data_out=16'h1;
17'h2923:	data_out=16'h6;
17'h2924:	data_out=16'h4;
17'h2925:	data_out=16'h8003;
17'h2926:	data_out=16'h6;
17'h2927:	data_out=16'h3;
17'h2928:	data_out=16'h8001;
17'h2929:	data_out=16'h9;
17'h292a:	data_out=16'h8000;
17'h292b:	data_out=16'h7;
17'h292c:	data_out=16'h3;
17'h292d:	data_out=16'h8002;
17'h292e:	data_out=16'h3;
17'h292f:	data_out=16'h9;
17'h2930:	data_out=16'h5;
17'h2931:	data_out=16'h1;
17'h2932:	data_out=16'h7;
17'h2933:	data_out=16'h7;
17'h2934:	data_out=16'h8000;
17'h2935:	data_out=16'h8008;
17'h2936:	data_out=16'h8007;
17'h2937:	data_out=16'h3;
17'h2938:	data_out=16'h5;
17'h2939:	data_out=16'h2;
17'h293a:	data_out=16'h1;
17'h293b:	data_out=16'h8005;
17'h293c:	data_out=16'h3;
17'h293d:	data_out=16'h8003;
17'h293e:	data_out=16'h8006;
17'h293f:	data_out=16'h8004;
17'h2940:	data_out=16'h8003;
17'h2941:	data_out=16'h4;
17'h2942:	data_out=16'h8008;
17'h2943:	data_out=16'h8007;
17'h2944:	data_out=16'h8008;
17'h2945:	data_out=16'h8;
17'h2946:	data_out=16'h5;
17'h2947:	data_out=16'h8000;
17'h2948:	data_out=16'h8;
17'h2949:	data_out=16'h8005;
17'h294a:	data_out=16'h8002;
17'h294b:	data_out=16'h1;
17'h294c:	data_out=16'h2;
17'h294d:	data_out=16'h8008;
17'h294e:	data_out=16'h1;
17'h294f:	data_out=16'h8002;
17'h2950:	data_out=16'h3;
17'h2951:	data_out=16'h8002;
17'h2952:	data_out=16'h8004;
17'h2953:	data_out=16'h8007;
17'h2954:	data_out=16'h8000;
17'h2955:	data_out=16'h8002;
17'h2956:	data_out=16'h6;
17'h2957:	data_out=16'h8005;
17'h2958:	data_out=16'h9;
17'h2959:	data_out=16'h8002;
17'h295a:	data_out=16'h8001;
17'h295b:	data_out=16'h3;
17'h295c:	data_out=16'h3;
17'h295d:	data_out=16'h2;
17'h295e:	data_out=16'h8;
17'h295f:	data_out=16'h8008;
17'h2960:	data_out=16'h8002;
17'h2961:	data_out=16'h8009;
17'h2962:	data_out=16'h8006;
17'h2963:	data_out=16'h8001;
17'h2964:	data_out=16'h8;
17'h2965:	data_out=16'h7;
17'h2966:	data_out=16'h8;
17'h2967:	data_out=16'h7;
17'h2968:	data_out=16'h8006;
17'h2969:	data_out=16'h8003;
17'h296a:	data_out=16'h8001;
17'h296b:	data_out=16'h5;
17'h296c:	data_out=16'h8002;
17'h296d:	data_out=16'h9;
17'h296e:	data_out=16'h8006;
17'h296f:	data_out=16'h8008;
17'h2970:	data_out=16'h8002;
17'h2971:	data_out=16'h8001;
17'h2972:	data_out=16'h8006;
17'h2973:	data_out=16'h7;
17'h2974:	data_out=16'h6;
17'h2975:	data_out=16'h9;
17'h2976:	data_out=16'h8007;
17'h2977:	data_out=16'h6;
17'h2978:	data_out=16'h8002;
17'h2979:	data_out=16'h2;
17'h297a:	data_out=16'h0;
17'h297b:	data_out=16'h8008;
17'h297c:	data_out=16'h8005;
17'h297d:	data_out=16'h8001;
17'h297e:	data_out=16'h8007;
17'h297f:	data_out=16'h2;
17'h2980:	data_out=16'h8000;
17'h2981:	data_out=16'h8005;
17'h2982:	data_out=16'h8009;
17'h2983:	data_out=16'h8001;
17'h2984:	data_out=16'h8006;
17'h2985:	data_out=16'h8;
17'h2986:	data_out=16'h8004;
17'h2987:	data_out=16'h8004;
17'h2988:	data_out=16'h8004;
17'h2989:	data_out=16'h5;
17'h298a:	data_out=16'h8008;
17'h298b:	data_out=16'h3;
17'h298c:	data_out=16'h5;
17'h298d:	data_out=16'h8004;
17'h298e:	data_out=16'h4;
17'h298f:	data_out=16'h8006;
17'h2990:	data_out=16'h4;
17'h2991:	data_out=16'h8;
17'h2992:	data_out=16'h8009;
17'h2993:	data_out=16'h1;
17'h2994:	data_out=16'h7;
17'h2995:	data_out=16'h8006;
17'h2996:	data_out=16'h8002;
17'h2997:	data_out=16'h8004;
17'h2998:	data_out=16'h5;
17'h2999:	data_out=16'h8;
17'h299a:	data_out=16'h8003;
17'h299b:	data_out=16'h9;
17'h299c:	data_out=16'h8002;
17'h299d:	data_out=16'h8002;
17'h299e:	data_out=16'h1;
17'h299f:	data_out=16'h6;
17'h29a0:	data_out=16'h3;
17'h29a1:	data_out=16'h2;
17'h29a2:	data_out=16'h8004;
17'h29a3:	data_out=16'h6;
17'h29a4:	data_out=16'h1;
17'h29a5:	data_out=16'h1;
17'h29a6:	data_out=16'h8007;
17'h29a7:	data_out=16'h5;
17'h29a8:	data_out=16'h8003;
17'h29a9:	data_out=16'h8006;
17'h29aa:	data_out=16'h8001;
17'h29ab:	data_out=16'h8008;
17'h29ac:	data_out=16'h8001;
17'h29ad:	data_out=16'h8006;
17'h29ae:	data_out=16'h8005;
17'h29af:	data_out=16'h8006;
17'h29b0:	data_out=16'h8008;
17'h29b1:	data_out=16'h8004;
17'h29b2:	data_out=16'h4;
17'h29b3:	data_out=16'h9;
17'h29b4:	data_out=16'h8001;
17'h29b5:	data_out=16'h8007;
17'h29b6:	data_out=16'h8004;
17'h29b7:	data_out=16'h8006;
17'h29b8:	data_out=16'h8008;
17'h29b9:	data_out=16'h2;
17'h29ba:	data_out=16'h8006;
17'h29bb:	data_out=16'h8001;
17'h29bc:	data_out=16'h8009;
17'h29bd:	data_out=16'h5;
17'h29be:	data_out=16'h8004;
17'h29bf:	data_out=16'h3;
17'h29c0:	data_out=16'h8003;
17'h29c1:	data_out=16'h1;
17'h29c2:	data_out=16'h8000;
17'h29c3:	data_out=16'h7;
17'h29c4:	data_out=16'h8007;
17'h29c5:	data_out=16'h2;
17'h29c6:	data_out=16'h3;
17'h29c7:	data_out=16'h8001;
17'h29c8:	data_out=16'h5;
17'h29c9:	data_out=16'h8007;
17'h29ca:	data_out=16'h1;
17'h29cb:	data_out=16'h8005;
17'h29cc:	data_out=16'h8004;
17'h29cd:	data_out=16'h5;
17'h29ce:	data_out=16'h8002;
17'h29cf:	data_out=16'h8002;
17'h29d0:	data_out=16'h8008;
17'h29d1:	data_out=16'h8007;
17'h29d2:	data_out=16'h8002;
17'h29d3:	data_out=16'h8001;
17'h29d4:	data_out=16'h8004;
17'h29d5:	data_out=16'h3;
17'h29d6:	data_out=16'h3;
17'h29d7:	data_out=16'h8003;
17'h29d8:	data_out=16'h8005;
17'h29d9:	data_out=16'h6;
17'h29da:	data_out=16'h4;
17'h29db:	data_out=16'h8004;
17'h29dc:	data_out=16'h1;
17'h29dd:	data_out=16'h8009;
17'h29de:	data_out=16'h8;
17'h29df:	data_out=16'h8;
17'h29e0:	data_out=16'h1;
17'h29e1:	data_out=16'h8001;
17'h29e2:	data_out=16'h5;
17'h29e3:	data_out=16'h3;
17'h29e4:	data_out=16'h8008;
17'h29e5:	data_out=16'h8001;
17'h29e6:	data_out=16'h8006;
17'h29e7:	data_out=16'h6;
17'h29e8:	data_out=16'h1;
17'h29e9:	data_out=16'h3;
17'h29ea:	data_out=16'h8008;
17'h29eb:	data_out=16'h7;
17'h29ec:	data_out=16'h8001;
17'h29ed:	data_out=16'h8000;
17'h29ee:	data_out=16'h8005;
17'h29ef:	data_out=16'h8000;
17'h29f0:	data_out=16'h2;
17'h29f1:	data_out=16'h2;
17'h29f2:	data_out=16'h8;
17'h29f3:	data_out=16'h7;
17'h29f4:	data_out=16'h8004;
17'h29f5:	data_out=16'h2;
17'h29f6:	data_out=16'h8006;
17'h29f7:	data_out=16'h0;
17'h29f8:	data_out=16'h8001;
17'h29f9:	data_out=16'h8;
17'h29fa:	data_out=16'h5;
17'h29fb:	data_out=16'h9;
17'h29fc:	data_out=16'h8;
17'h29fd:	data_out=16'h4;
17'h29fe:	data_out=16'h8;
17'h29ff:	data_out=16'h0;
17'h2a00:	data_out=16'h8007;
17'h2a01:	data_out=16'h4;
17'h2a02:	data_out=16'h8005;
17'h2a03:	data_out=16'h8006;
17'h2a04:	data_out=16'h8006;
17'h2a05:	data_out=16'h8003;
17'h2a06:	data_out=16'h8009;
17'h2a07:	data_out=16'h4;
17'h2a08:	data_out=16'h8009;
17'h2a09:	data_out=16'h8007;
17'h2a0a:	data_out=16'h2;
17'h2a0b:	data_out=16'h8000;
17'h2a0c:	data_out=16'h1;
17'h2a0d:	data_out=16'h6;
17'h2a0e:	data_out=16'h9;
17'h2a0f:	data_out=16'h8006;
17'h2a10:	data_out=16'h8000;
17'h2a11:	data_out=16'h8;
17'h2a12:	data_out=16'h8008;
17'h2a13:	data_out=16'h5;
17'h2a14:	data_out=16'h1;
17'h2a15:	data_out=16'h8004;
17'h2a16:	data_out=16'h8004;
17'h2a17:	data_out=16'h9;
17'h2a18:	data_out=16'h8006;
17'h2a19:	data_out=16'h8008;
17'h2a1a:	data_out=16'h9;
17'h2a1b:	data_out=16'h8006;
17'h2a1c:	data_out=16'h5;
17'h2a1d:	data_out=16'h7;
17'h2a1e:	data_out=16'h3;
17'h2a1f:	data_out=16'h7;
17'h2a20:	data_out=16'h2;
17'h2a21:	data_out=16'h7;
17'h2a22:	data_out=16'h8008;
17'h2a23:	data_out=16'h5;
17'h2a24:	data_out=16'h8005;
17'h2a25:	data_out=16'h8007;
17'h2a26:	data_out=16'h0;
17'h2a27:	data_out=16'h8005;
17'h2a28:	data_out=16'h8006;
17'h2a29:	data_out=16'h8007;
17'h2a2a:	data_out=16'h4;
17'h2a2b:	data_out=16'h5;
17'h2a2c:	data_out=16'h9;
17'h2a2d:	data_out=16'h4;
17'h2a2e:	data_out=16'h8;
17'h2a2f:	data_out=16'h8001;
17'h2a30:	data_out=16'h3;
17'h2a31:	data_out=16'h8009;
17'h2a32:	data_out=16'h8005;
17'h2a33:	data_out=16'h8005;
17'h2a34:	data_out=16'h8004;
17'h2a35:	data_out=16'h8001;
17'h2a36:	data_out=16'h8005;
17'h2a37:	data_out=16'h8001;
17'h2a38:	data_out=16'h0;
17'h2a39:	data_out=16'h8005;
17'h2a3a:	data_out=16'h2;
17'h2a3b:	data_out=16'h8004;
17'h2a3c:	data_out=16'h8007;
17'h2a3d:	data_out=16'h8004;
17'h2a3e:	data_out=16'h8006;
17'h2a3f:	data_out=16'h4;
17'h2a40:	data_out=16'h8006;
17'h2a41:	data_out=16'h8005;
17'h2a42:	data_out=16'h0;
17'h2a43:	data_out=16'h8003;
17'h2a44:	data_out=16'h8003;
17'h2a45:	data_out=16'h8008;
17'h2a46:	data_out=16'h2;
17'h2a47:	data_out=16'h0;
17'h2a48:	data_out=16'h8006;
17'h2a49:	data_out=16'h8003;
17'h2a4a:	data_out=16'h8004;
17'h2a4b:	data_out=16'h8006;
17'h2a4c:	data_out=16'h8009;
17'h2a4d:	data_out=16'h8005;
17'h2a4e:	data_out=16'h2;
17'h2a4f:	data_out=16'h4;
17'h2a50:	data_out=16'h8004;
17'h2a51:	data_out=16'h6;
17'h2a52:	data_out=16'h8;
17'h2a53:	data_out=16'h0;
17'h2a54:	data_out=16'h8004;
17'h2a55:	data_out=16'h8006;
17'h2a56:	data_out=16'h9;
17'h2a57:	data_out=16'h5;
17'h2a58:	data_out=16'h8002;
17'h2a59:	data_out=16'h2;
17'h2a5a:	data_out=16'h8008;
17'h2a5b:	data_out=16'h0;
17'h2a5c:	data_out=16'h7;
17'h2a5d:	data_out=16'h8005;
17'h2a5e:	data_out=16'h8005;
17'h2a5f:	data_out=16'h8008;
17'h2a60:	data_out=16'h8000;
17'h2a61:	data_out=16'h5;
17'h2a62:	data_out=16'h8002;
17'h2a63:	data_out=16'h6;
17'h2a64:	data_out=16'h6;
17'h2a65:	data_out=16'h9;
17'h2a66:	data_out=16'h8003;
17'h2a67:	data_out=16'h8009;
17'h2a68:	data_out=16'h8004;
17'h2a69:	data_out=16'h3;
17'h2a6a:	data_out=16'h8006;
17'h2a6b:	data_out=16'h8003;
17'h2a6c:	data_out=16'h7;
17'h2a6d:	data_out=16'h5;
17'h2a6e:	data_out=16'h8008;
17'h2a6f:	data_out=16'h8007;
17'h2a70:	data_out=16'h1;
17'h2a71:	data_out=16'h9;
17'h2a72:	data_out=16'h3;
17'h2a73:	data_out=16'h6;
17'h2a74:	data_out=16'h8007;
17'h2a75:	data_out=16'h3;
17'h2a76:	data_out=16'h3;
17'h2a77:	data_out=16'h8000;
17'h2a78:	data_out=16'h8004;
17'h2a79:	data_out=16'h4;
17'h2a7a:	data_out=16'h9;
17'h2a7b:	data_out=16'h8006;
17'h2a7c:	data_out=16'h8;
17'h2a7d:	data_out=16'h8005;
17'h2a7e:	data_out=16'h8006;
17'h2a7f:	data_out=16'h8001;
17'h2a80:	data_out=16'h8009;
17'h2a81:	data_out=16'h2;
17'h2a82:	data_out=16'h8004;
17'h2a83:	data_out=16'h6;
17'h2a84:	data_out=16'h1;
17'h2a85:	data_out=16'h2;
17'h2a86:	data_out=16'h6;
17'h2a87:	data_out=16'h7;
17'h2a88:	data_out=16'h8005;
17'h2a89:	data_out=16'h8009;
17'h2a8a:	data_out=16'h8005;
17'h2a8b:	data_out=16'h8007;
17'h2a8c:	data_out=16'h5;
17'h2a8d:	data_out=16'h8004;
17'h2a8e:	data_out=16'h8004;
17'h2a8f:	data_out=16'h8003;
17'h2a90:	data_out=16'h8005;
17'h2a91:	data_out=16'h8;
17'h2a92:	data_out=16'h8006;
17'h2a93:	data_out=16'h8003;
17'h2a94:	data_out=16'h1;
17'h2a95:	data_out=16'h6;
17'h2a96:	data_out=16'h6;
17'h2a97:	data_out=16'h6;
17'h2a98:	data_out=16'h1;
17'h2a99:	data_out=16'h6;
17'h2a9a:	data_out=16'h9;
17'h2a9b:	data_out=16'h8000;
17'h2a9c:	data_out=16'h8008;
17'h2a9d:	data_out=16'h8006;
17'h2a9e:	data_out=16'h8;
17'h2a9f:	data_out=16'h8007;
17'h2aa0:	data_out=16'h5;
17'h2aa1:	data_out=16'h8006;
17'h2aa2:	data_out=16'h8;
17'h2aa3:	data_out=16'h8003;
17'h2aa4:	data_out=16'h5;
17'h2aa5:	data_out=16'h6;
17'h2aa6:	data_out=16'h8005;
17'h2aa7:	data_out=16'h8008;
17'h2aa8:	data_out=16'h6;
17'h2aa9:	data_out=16'h8001;
17'h2aaa:	data_out=16'h8006;
17'h2aab:	data_out=16'h1;
17'h2aac:	data_out=16'h3;
17'h2aad:	data_out=16'h8001;
17'h2aae:	data_out=16'h7;
17'h2aaf:	data_out=16'h8;
17'h2ab0:	data_out=16'h8003;
17'h2ab1:	data_out=16'h8008;
17'h2ab2:	data_out=16'h8004;
17'h2ab3:	data_out=16'h8;
17'h2ab4:	data_out=16'h7;
17'h2ab5:	data_out=16'h8007;
17'h2ab6:	data_out=16'h5;
17'h2ab7:	data_out=16'h8001;
17'h2ab8:	data_out=16'h8;
17'h2ab9:	data_out=16'h5;
17'h2aba:	data_out=16'h7;
17'h2abb:	data_out=16'h8009;
17'h2abc:	data_out=16'h8;
17'h2abd:	data_out=16'h6;
17'h2abe:	data_out=16'h8007;
17'h2abf:	data_out=16'h4;
17'h2ac0:	data_out=16'h8009;
17'h2ac1:	data_out=16'h8008;
17'h2ac2:	data_out=16'h8008;
17'h2ac3:	data_out=16'h6;
17'h2ac4:	data_out=16'h7;
17'h2ac5:	data_out=16'h8004;
17'h2ac6:	data_out=16'h6;
17'h2ac7:	data_out=16'h4;
17'h2ac8:	data_out=16'h3;
17'h2ac9:	data_out=16'h8009;
17'h2aca:	data_out=16'h8004;
17'h2acb:	data_out=16'h8002;
17'h2acc:	data_out=16'h8001;
17'h2acd:	data_out=16'h8006;
17'h2ace:	data_out=16'h8004;
17'h2acf:	data_out=16'h5;
17'h2ad0:	data_out=16'h8004;
17'h2ad1:	data_out=16'h1;
17'h2ad2:	data_out=16'h4;
17'h2ad3:	data_out=16'h8006;
17'h2ad4:	data_out=16'h2;
17'h2ad5:	data_out=16'h8001;
17'h2ad6:	data_out=16'h2;
17'h2ad7:	data_out=16'h1;
17'h2ad8:	data_out=16'h8005;
17'h2ad9:	data_out=16'h0;
17'h2ada:	data_out=16'h1;
17'h2adb:	data_out=16'h8006;
17'h2adc:	data_out=16'h8003;
17'h2add:	data_out=16'h3;
17'h2ade:	data_out=16'h6;
17'h2adf:	data_out=16'h8003;
17'h2ae0:	data_out=16'h5;
17'h2ae1:	data_out=16'h7;
17'h2ae2:	data_out=16'h8006;
17'h2ae3:	data_out=16'h2;
17'h2ae4:	data_out=16'h8006;
17'h2ae5:	data_out=16'h8009;
17'h2ae6:	data_out=16'h8003;
17'h2ae7:	data_out=16'h6;
17'h2ae8:	data_out=16'h8008;
17'h2ae9:	data_out=16'h2;
17'h2aea:	data_out=16'h8005;
17'h2aeb:	data_out=16'h8000;
17'h2aec:	data_out=16'h5;
17'h2aed:	data_out=16'h0;
17'h2aee:	data_out=16'h8004;
17'h2aef:	data_out=16'h8008;
17'h2af0:	data_out=16'h8008;
17'h2af1:	data_out=16'h9;
17'h2af2:	data_out=16'h8005;
17'h2af3:	data_out=16'h3;
17'h2af4:	data_out=16'h8001;
17'h2af5:	data_out=16'h6;
17'h2af6:	data_out=16'h8005;
17'h2af7:	data_out=16'h3;
17'h2af8:	data_out=16'h8003;
17'h2af9:	data_out=16'h6;
17'h2afa:	data_out=16'h6;
17'h2afb:	data_out=16'h3;
17'h2afc:	data_out=16'h8000;
17'h2afd:	data_out=16'h3;
17'h2afe:	data_out=16'h9;
17'h2aff:	data_out=16'h8005;
17'h2b00:	data_out=16'h6;
17'h2b01:	data_out=16'h21;
17'h2b02:	data_out=16'h28;
17'h2b03:	data_out=16'h2c;
17'h2b04:	data_out=16'h8;
17'h2b05:	data_out=16'h1d;
17'h2b06:	data_out=16'h1d;
17'h2b07:	data_out=16'h8;
17'h2b08:	data_out=16'h10;
17'h2b09:	data_out=16'h8007;
17'h2b0a:	data_out=16'h1d;
17'h2b0b:	data_out=16'h30;
17'h2b0c:	data_out=16'h8004;
17'h2b0d:	data_out=16'h35;
17'h2b0e:	data_out=16'hc;
17'h2b0f:	data_out=16'h2b;
17'h2b10:	data_out=16'h16;
17'h2b11:	data_out=16'h13;
17'h2b12:	data_out=16'h21;
17'h2b13:	data_out=16'h30;
17'h2b14:	data_out=16'h57;
17'h2b15:	data_out=16'h1a;
17'h2b16:	data_out=16'h24;
17'h2b17:	data_out=16'h63;
17'h2b18:	data_out=16'h8004;
17'h2b19:	data_out=16'h800f;
17'h2b1a:	data_out=16'h10;
17'h2b1b:	data_out=16'h31;
17'h2b1c:	data_out=16'h2f;
17'h2b1d:	data_out=16'h25;
17'h2b1e:	data_out=16'h3b;
17'h2b1f:	data_out=16'h1f;
17'h2b20:	data_out=16'h2d;
17'h2b21:	data_out=16'hd;
17'h2b22:	data_out=16'h1d;
17'h2b23:	data_out=16'h3;
17'h2b24:	data_out=16'h2;
17'h2b25:	data_out=16'h9;
17'h2b26:	data_out=16'h8001;
17'h2b27:	data_out=16'h25;
17'h2b28:	data_out=16'h7;
17'h2b29:	data_out=16'h2a;
17'h2b2a:	data_out=16'h18;
17'h2b2b:	data_out=16'h8002;
17'h2b2c:	data_out=16'h33;
17'h2b2d:	data_out=16'h13;
17'h2b2e:	data_out=16'h2f;
17'h2b2f:	data_out=16'h36;
17'h2b30:	data_out=16'h3b;
17'h2b31:	data_out=16'h15;
17'h2b32:	data_out=16'h31;
17'h2b33:	data_out=16'h4b;
17'h2b34:	data_out=16'h2;
17'h2b35:	data_out=16'hb;
17'h2b36:	data_out=16'h27;
17'h2b37:	data_out=16'h27;
17'h2b38:	data_out=16'h8001;
17'h2b39:	data_out=16'h28;
17'h2b3a:	data_out=16'h16;
17'h2b3b:	data_out=16'h8003;
17'h2b3c:	data_out=16'h31;
17'h2b3d:	data_out=16'hc;
17'h2b3e:	data_out=16'h6;
17'h2b3f:	data_out=16'h16;
17'h2b40:	data_out=16'h14;
17'h2b41:	data_out=16'h28;
17'h2b42:	data_out=16'h8000;
17'h2b43:	data_out=16'h11;
17'h2b44:	data_out=16'h19;
17'h2b45:	data_out=16'h17;
17'h2b46:	data_out=16'h2b;
17'h2b47:	data_out=16'h7;
17'h2b48:	data_out=16'h1a;
17'h2b49:	data_out=16'h3;
17'h2b4a:	data_out=16'h9;
17'h2b4b:	data_out=16'h8001;
17'h2b4c:	data_out=16'h8005;
17'h2b4d:	data_out=16'h1c;
17'h2b4e:	data_out=16'h10;
17'h2b4f:	data_out=16'h8;
17'h2b50:	data_out=16'he;
17'h2b51:	data_out=16'h2e;
17'h2b52:	data_out=16'h6;
17'h2b53:	data_out=16'h3a;
17'h2b54:	data_out=16'h41;
17'h2b55:	data_out=16'h38;
17'h2b56:	data_out=16'h33;
17'h2b57:	data_out=16'h15;
17'h2b58:	data_out=16'h2a;
17'h2b59:	data_out=16'h1e;
17'h2b5a:	data_out=16'h21;
17'h2b5b:	data_out=16'h37;
17'h2b5c:	data_out=16'h1a;
17'h2b5d:	data_out=16'h25;
17'h2b5e:	data_out=16'h2b;
17'h2b5f:	data_out=16'h13;
17'h2b60:	data_out=16'h15;
17'h2b61:	data_out=16'h2e;
17'h2b62:	data_out=16'h32;
17'h2b63:	data_out=16'h4b;
17'h2b64:	data_out=16'h3;
17'h2b65:	data_out=16'h13;
17'h2b66:	data_out=16'h800c;
17'h2b67:	data_out=16'h1d;
17'h2b68:	data_out=16'h4;
17'h2b69:	data_out=16'h15;
17'h2b6a:	data_out=16'h13;
17'h2b6b:	data_out=16'hb;
17'h2b6c:	data_out=16'h2c;
17'h2b6d:	data_out=16'h46;
17'h2b6e:	data_out=16'h5;
17'h2b6f:	data_out=16'h25;
17'h2b70:	data_out=16'hd;
17'h2b71:	data_out=16'h21;
17'h2b72:	data_out=16'h1a;
17'h2b73:	data_out=16'h24;
17'h2b74:	data_out=16'h34;
17'h2b75:	data_out=16'h1b;
17'h2b76:	data_out=16'hc;
17'h2b77:	data_out=16'h7;
17'h2b78:	data_out=16'h3;
17'h2b79:	data_out=16'h24;
17'h2b7a:	data_out=16'h4a;
17'h2b7b:	data_out=16'hc;
17'h2b7c:	data_out=16'h19;
17'h2b7d:	data_out=16'h1d;
17'h2b7e:	data_out=16'h8003;
17'h2b7f:	data_out=16'hb;
17'h2b80:	data_out=16'h46;
17'h2b81:	data_out=16'h804d;
17'h2b82:	data_out=16'h814a;
17'h2b83:	data_out=16'h814a;
17'h2b84:	data_out=16'h9b;
17'h2b85:	data_out=16'h80e4;
17'h2b86:	data_out=16'h8101;
17'h2b87:	data_out=16'h8020;
17'h2b88:	data_out=16'h2;
17'h2b89:	data_out=16'h8034;
17'h2b8a:	data_out=16'hd9;
17'h2b8b:	data_out=16'h8053;
17'h2b8c:	data_out=16'h206;
17'h2b8d:	data_out=16'h8171;
17'h2b8e:	data_out=16'h805b;
17'h2b8f:	data_out=16'h81d4;
17'h2b90:	data_out=16'h8055;
17'h2b91:	data_out=16'hcc;
17'h2b92:	data_out=16'h8117;
17'h2b93:	data_out=16'h8129;
17'h2b94:	data_out=16'h820b;
17'h2b95:	data_out=16'h80a6;
17'h2b96:	data_out=16'h80c0;
17'h2b97:	data_out=16'h81fe;
17'h2b98:	data_out=16'h8087;
17'h2b99:	data_out=16'h113;
17'h2b9a:	data_out=16'hb8;
17'h2b9b:	data_out=16'h8196;
17'h2b9c:	data_out=16'h819f;
17'h2b9d:	data_out=16'h800c;
17'h2b9e:	data_out=16'h821b;
17'h2b9f:	data_out=16'h81b4;
17'h2ba0:	data_out=16'h8132;
17'h2ba1:	data_out=16'h8064;
17'h2ba2:	data_out=16'h8074;
17'h2ba3:	data_out=16'h58;
17'h2ba4:	data_out=16'h51;
17'h2ba5:	data_out=16'hd;
17'h2ba6:	data_out=16'h806d;
17'h2ba7:	data_out=16'h8021;
17'h2ba8:	data_out=16'h8058;
17'h2ba9:	data_out=16'h8174;
17'h2baa:	data_out=16'h80e3;
17'h2bab:	data_out=16'h2e;
17'h2bac:	data_out=16'h807a;
17'h2bad:	data_out=16'h9a;
17'h2bae:	data_out=16'h8196;
17'h2baf:	data_out=16'h8124;
17'h2bb0:	data_out=16'h101;
17'h2bb1:	data_out=16'hd8;
17'h2bb2:	data_out=16'h105;
17'h2bb3:	data_out=16'h8224;
17'h2bb4:	data_out=16'h8b;
17'h2bb5:	data_out=16'h12c;
17'h2bb6:	data_out=16'h8104;
17'h2bb7:	data_out=16'h817b;
17'h2bb8:	data_out=16'h815b;
17'h2bb9:	data_out=16'h81fa;
17'h2bba:	data_out=16'h80b3;
17'h2bbb:	data_out=16'h12a;
17'h2bbc:	data_out=16'h8100;
17'h2bbd:	data_out=16'h80b8;
17'h2bbe:	data_out=16'h8065;
17'h2bbf:	data_out=16'h8067;
17'h2bc0:	data_out=16'h80af;
17'h2bc1:	data_out=16'h812f;
17'h2bc2:	data_out=16'h105;
17'h2bc3:	data_out=16'h814f;
17'h2bc4:	data_out=16'h45;
17'h2bc5:	data_out=16'h80bd;
17'h2bc6:	data_out=16'h80f2;
17'h2bc7:	data_out=16'h80ae;
17'h2bc8:	data_out=16'h810e;
17'h2bc9:	data_out=16'h800a;
17'h2bca:	data_out=16'h21;
17'h2bcb:	data_out=16'h149;
17'h2bcc:	data_out=16'h8000;
17'h2bcd:	data_out=16'h808b;
17'h2bce:	data_out=16'h809f;
17'h2bcf:	data_out=16'h27;
17'h2bd0:	data_out=16'h8128;
17'h2bd1:	data_out=16'h8194;
17'h2bd2:	data_out=16'h15;
17'h2bd3:	data_out=16'h8113;
17'h2bd4:	data_out=16'h8114;
17'h2bd5:	data_out=16'h8156;
17'h2bd6:	data_out=16'h8135;
17'h2bd7:	data_out=16'h8107;
17'h2bd8:	data_out=16'h8137;
17'h2bd9:	data_out=16'h809a;
17'h2bda:	data_out=16'h818d;
17'h2bdb:	data_out=16'h8123;
17'h2bdc:	data_out=16'h804d;
17'h2bdd:	data_out=16'h80ca;
17'h2bde:	data_out=16'h80e0;
17'h2bdf:	data_out=16'h80a7;
17'h2be0:	data_out=16'h8055;
17'h2be1:	data_out=16'h80a1;
17'h2be2:	data_out=16'h81e7;
17'h2be3:	data_out=16'h8208;
17'h2be4:	data_out=16'h39;
17'h2be5:	data_out=16'hb7;
17'h2be6:	data_out=16'hda;
17'h2be7:	data_out=16'h8107;
17'h2be8:	data_out=16'h8055;
17'h2be9:	data_out=16'h803d;
17'h2bea:	data_out=16'h8067;
17'h2beb:	data_out=16'h8015;
17'h2bec:	data_out=16'h22;
17'h2bed:	data_out=16'h8218;
17'h2bee:	data_out=16'h805a;
17'h2bef:	data_out=16'h8087;
17'h2bf0:	data_out=16'h8057;
17'h2bf1:	data_out=16'h81a9;
17'h2bf2:	data_out=16'h80da;
17'h2bf3:	data_out=16'h80d7;
17'h2bf4:	data_out=16'h109;
17'h2bf5:	data_out=16'h80f8;
17'h2bf6:	data_out=16'h30;
17'h2bf7:	data_out=16'h804b;
17'h2bf8:	data_out=16'h80c4;
17'h2bf9:	data_out=16'h81cf;
17'h2bfa:	data_out=16'h8213;
17'h2bfb:	data_out=16'h8057;
17'h2bfc:	data_out=16'h80c4;
17'h2bfd:	data_out=16'h819b;
17'h2bfe:	data_out=16'h8028;
17'h2bff:	data_out=16'h809c;
17'h2c00:	data_out=16'h81aa;
17'h2c01:	data_out=16'h81c4;
17'h2c02:	data_out=16'h8139;
17'h2c03:	data_out=16'h80fc;
17'h2c04:	data_out=16'h1e4;
17'h2c05:	data_out=16'hf;
17'h2c06:	data_out=16'h58;
17'h2c07:	data_out=16'h33;
17'h2c08:	data_out=16'h8108;
17'h2c09:	data_out=16'h8041;
17'h2c0a:	data_out=16'h816b;
17'h2c0b:	data_out=16'h8092;
17'h2c0c:	data_out=16'h163;
17'h2c0d:	data_out=16'h80a8;
17'h2c0e:	data_out=16'h801a;
17'h2c0f:	data_out=16'h81a1;
17'h2c10:	data_out=16'h8093;
17'h2c11:	data_out=16'h1e;
17'h2c12:	data_out=16'h812a;
17'h2c13:	data_out=16'h80cc;
17'h2c14:	data_out=16'h826d;
17'h2c15:	data_out=16'h808a;
17'h2c16:	data_out=16'h80a3;
17'h2c17:	data_out=16'h828d;
17'h2c18:	data_out=16'h8017;
17'h2c19:	data_out=16'h65;
17'h2c1a:	data_out=16'h239;
17'h2c1b:	data_out=16'h8232;
17'h2c1c:	data_out=16'h820b;
17'h2c1d:	data_out=16'h81f7;
17'h2c1e:	data_out=16'h8257;
17'h2c1f:	data_out=16'h8066;
17'h2c20:	data_out=16'h815c;
17'h2c21:	data_out=16'h8020;
17'h2c22:	data_out=16'h8034;
17'h2c23:	data_out=16'h58;
17'h2c24:	data_out=16'h52;
17'h2c25:	data_out=16'h92;
17'h2c26:	data_out=16'h8220;
17'h2c27:	data_out=16'h81ee;
17'h2c28:	data_out=16'h8018;
17'h2c29:	data_out=16'h8208;
17'h2c2a:	data_out=16'h81a6;
17'h2c2b:	data_out=16'h80ba;
17'h2c2c:	data_out=16'h804a;
17'h2c2d:	data_out=16'h80f6;
17'h2c2e:	data_out=16'h8184;
17'h2c2f:	data_out=16'h812a;
17'h2c30:	data_out=16'h23c;
17'h2c31:	data_out=16'h80fe;
17'h2c32:	data_out=16'h22f;
17'h2c33:	data_out=16'h8261;
17'h2c34:	data_out=16'h8182;
17'h2c35:	data_out=16'h16e;
17'h2c36:	data_out=16'h811f;
17'h2c37:	data_out=16'h8143;
17'h2c38:	data_out=16'h81d7;
17'h2c39:	data_out=16'h824d;
17'h2c3a:	data_out=16'h806d;
17'h2c3b:	data_out=16'h2b;
17'h2c3c:	data_out=16'h81ce;
17'h2c3d:	data_out=16'h815d;
17'h2c3e:	data_out=16'h8015;
17'h2c3f:	data_out=16'ha7;
17'h2c40:	data_out=16'h1aa;
17'h2c41:	data_out=16'h80d1;
17'h2c42:	data_out=16'h154;
17'h2c43:	data_out=16'h32;
17'h2c44:	data_out=16'h807b;
17'h2c45:	data_out=16'h8093;
17'h2c46:	data_out=16'h81b7;
17'h2c47:	data_out=16'h8033;
17'h2c48:	data_out=16'h80d0;
17'h2c49:	data_out=16'h98;
17'h2c4a:	data_out=16'h152;
17'h2c4b:	data_out=16'h149;
17'h2c4c:	data_out=16'h131;
17'h2c4d:	data_out=16'h8048;
17'h2c4e:	data_out=16'h80c6;
17'h2c4f:	data_out=16'h13a;
17'h2c50:	data_out=16'h10a;
17'h2c51:	data_out=16'h8166;
17'h2c52:	data_out=16'h35;
17'h2c53:	data_out=16'h826e;
17'h2c54:	data_out=16'h816b;
17'h2c55:	data_out=16'h8140;
17'h2c56:	data_out=16'h8103;
17'h2c57:	data_out=16'h80b1;
17'h2c58:	data_out=16'h812e;
17'h2c59:	data_out=16'h113;
17'h2c5a:	data_out=16'h827f;
17'h2c5b:	data_out=16'h8133;
17'h2c5c:	data_out=16'h8101;
17'h2c5d:	data_out=16'h80a8;
17'h2c5e:	data_out=16'h80c1;
17'h2c5f:	data_out=16'h8044;
17'h2c60:	data_out=16'h8227;
17'h2c61:	data_out=16'h80b1;
17'h2c62:	data_out=16'h8209;
17'h2c63:	data_out=16'h824e;
17'h2c64:	data_out=16'h8127;
17'h2c65:	data_out=16'hb4;
17'h2c66:	data_out=16'h65;
17'h2c67:	data_out=16'h816b;
17'h2c68:	data_out=16'h801c;
17'h2c69:	data_out=16'h80f4;
17'h2c6a:	data_out=16'h801a;
17'h2c6b:	data_out=16'hde;
17'h2c6c:	data_out=16'h8197;
17'h2c6d:	data_out=16'h8267;
17'h2c6e:	data_out=16'h801d;
17'h2c6f:	data_out=16'he6;
17'h2c70:	data_out=16'h8019;
17'h2c71:	data_out=16'h815e;
17'h2c72:	data_out=16'h807b;
17'h2c73:	data_out=16'h8086;
17'h2c74:	data_out=16'h23b;
17'h2c75:	data_out=16'h8159;
17'h2c76:	data_out=16'h8149;
17'h2c77:	data_out=16'h126;
17'h2c78:	data_out=16'haf;
17'h2c79:	data_out=16'h8190;
17'h2c7a:	data_out=16'h8256;
17'h2c7b:	data_out=16'h8017;
17'h2c7c:	data_out=16'h804b;
17'h2c7d:	data_out=16'h8018;
17'h2c7e:	data_out=16'h80cd;
17'h2c7f:	data_out=16'h13d;
17'h2c80:	data_out=16'h86f8;
17'h2c81:	data_out=16'h843b;
17'h2c82:	data_out=16'h81f5;
17'h2c83:	data_out=16'h82df;
17'h2c84:	data_out=16'h2ce;
17'h2c85:	data_out=16'h2e1;
17'h2c86:	data_out=16'h19a;
17'h2c87:	data_out=16'h813b;
17'h2c88:	data_out=16'h8360;
17'h2c89:	data_out=16'h8458;
17'h2c8a:	data_out=16'h8578;
17'h2c8b:	data_out=16'h3ed;
17'h2c8c:	data_out=16'h3f0;
17'h2c8d:	data_out=16'h8029;
17'h2c8e:	data_out=16'h8080;
17'h2c8f:	data_out=16'h82a3;
17'h2c90:	data_out=16'h8449;
17'h2c91:	data_out=16'h46;
17'h2c92:	data_out=16'h822e;
17'h2c93:	data_out=16'h81af;
17'h2c94:	data_out=16'h81ec;
17'h2c95:	data_out=16'h8301;
17'h2c96:	data_out=16'h83be;
17'h2c97:	data_out=16'h80c3;
17'h2c98:	data_out=16'h823b;
17'h2c99:	data_out=16'h325;
17'h2c9a:	data_out=16'h463;
17'h2c9b:	data_out=16'h359;
17'h2c9c:	data_out=16'h80d6;
17'h2c9d:	data_out=16'h832a;
17'h2c9e:	data_out=16'h8149;
17'h2c9f:	data_out=16'h8103;
17'h2ca0:	data_out=16'h8212;
17'h2ca1:	data_out=16'h8071;
17'h2ca2:	data_out=16'h8280;
17'h2ca3:	data_out=16'h832d;
17'h2ca4:	data_out=16'h832e;
17'h2ca5:	data_out=16'h80c5;
17'h2ca6:	data_out=16'h868d;
17'h2ca7:	data_out=16'h81ec;
17'h2ca8:	data_out=16'h8055;
17'h2ca9:	data_out=16'h83b3;
17'h2caa:	data_out=16'h8601;
17'h2cab:	data_out=16'h14e;
17'h2cac:	data_out=16'h824c;
17'h2cad:	data_out=16'h8369;
17'h2cae:	data_out=16'h838c;
17'h2caf:	data_out=16'h809d;
17'h2cb0:	data_out=16'h4a4;
17'h2cb1:	data_out=16'h80ef;
17'h2cb2:	data_out=16'h490;
17'h2cb3:	data_out=16'h82b3;
17'h2cb4:	data_out=16'h83b6;
17'h2cb5:	data_out=16'h338;
17'h2cb6:	data_out=16'h836c;
17'h2cb7:	data_out=16'h81b9;
17'h2cb8:	data_out=16'h828b;
17'h2cb9:	data_out=16'h820b;
17'h2cba:	data_out=16'h864a;
17'h2cbb:	data_out=16'h8;
17'h2cbc:	data_out=16'h810c;
17'h2cbd:	data_out=16'h866d;
17'h2cbe:	data_out=16'h804f;
17'h2cbf:	data_out=16'h2f0;
17'h2cc0:	data_out=16'h80c1;
17'h2cc1:	data_out=16'h16b;
17'h2cc2:	data_out=16'h2c;
17'h2cc3:	data_out=16'h328;
17'h2cc4:	data_out=16'h8170;
17'h2cc5:	data_out=16'h8310;
17'h2cc6:	data_out=16'h3a;
17'h2cc7:	data_out=16'h854c;
17'h2cc8:	data_out=16'h80c6;
17'h2cc9:	data_out=16'h8131;
17'h2cca:	data_out=16'h112;
17'h2ccb:	data_out=16'h369;
17'h2ccc:	data_out=16'h8155;
17'h2ccd:	data_out=16'h8288;
17'h2cce:	data_out=16'h81e0;
17'h2ccf:	data_out=16'h81c5;
17'h2cd0:	data_out=16'h81be;
17'h2cd1:	data_out=16'h80c7;
17'h2cd2:	data_out=16'h839b;
17'h2cd3:	data_out=16'h448;
17'h2cd4:	data_out=16'h82d8;
17'h2cd5:	data_out=16'h8130;
17'h2cd6:	data_out=16'h868e;
17'h2cd7:	data_out=16'h863e;
17'h2cd8:	data_out=16'h81d9;
17'h2cd9:	data_out=16'h82a7;
17'h2cda:	data_out=16'h4e4;
17'h2cdb:	data_out=16'h8123;
17'h2cdc:	data_out=16'h802b;
17'h2cdd:	data_out=16'h83c4;
17'h2cde:	data_out=16'h8008;
17'h2cdf:	data_out=16'h821d;
17'h2ce0:	data_out=16'h878d;
17'h2ce1:	data_out=16'h8161;
17'h2ce2:	data_out=16'h439;
17'h2ce3:	data_out=16'h8249;
17'h2ce4:	data_out=16'h8333;
17'h2ce5:	data_out=16'h1aa;
17'h2ce6:	data_out=16'h30d;
17'h2ce7:	data_out=16'h8244;
17'h2ce8:	data_out=16'h8062;
17'h2ce9:	data_out=16'h8506;
17'h2cea:	data_out=16'h8093;
17'h2ceb:	data_out=16'h28b;
17'h2cec:	data_out=16'h89f4;
17'h2ced:	data_out=16'h826f;
17'h2cee:	data_out=16'h80a2;
17'h2cef:	data_out=16'h318;
17'h2cf0:	data_out=16'h8089;
17'h2cf1:	data_out=16'h8376;
17'h2cf2:	data_out=16'h8296;
17'h2cf3:	data_out=16'h80dd;
17'h2cf4:	data_out=16'h4b2;
17'h2cf5:	data_out=16'h65f;
17'h2cf6:	data_out=16'h2;
17'h2cf7:	data_out=16'h8196;
17'h2cf8:	data_out=16'h4cc;
17'h2cf9:	data_out=16'h84a0;
17'h2cfa:	data_out=16'h81fb;
17'h2cfb:	data_out=16'h804e;
17'h2cfc:	data_out=16'h812e;
17'h2cfd:	data_out=16'h36a;
17'h2cfe:	data_out=16'h83c8;
17'h2cff:	data_out=16'h83a1;
17'h2d00:	data_out=16'h8a00;
17'h2d01:	data_out=16'h8910;
17'h2d02:	data_out=16'h8465;
17'h2d03:	data_out=16'h8090;
17'h2d04:	data_out=16'ha00;
17'h2d05:	data_out=16'h5e7;
17'h2d06:	data_out=16'h3e1;
17'h2d07:	data_out=16'h1ad;
17'h2d08:	data_out=16'h89b8;
17'h2d09:	data_out=16'h81d0;
17'h2d0a:	data_out=16'h8941;
17'h2d0b:	data_out=16'h4f;
17'h2d0c:	data_out=16'ha00;
17'h2d0d:	data_out=16'h812c;
17'h2d0e:	data_out=16'h80d8;
17'h2d0f:	data_out=16'h8539;
17'h2d10:	data_out=16'h80d6;
17'h2d11:	data_out=16'h3b1;
17'h2d12:	data_out=16'h81bd;
17'h2d13:	data_out=16'h80d7;
17'h2d14:	data_out=16'h86fc;
17'h2d15:	data_out=16'h8353;
17'h2d16:	data_out=16'h83a0;
17'h2d17:	data_out=16'h853d;
17'h2d18:	data_out=16'h83dd;
17'h2d19:	data_out=16'h4d6;
17'h2d1a:	data_out=16'ha00;
17'h2d1b:	data_out=16'h810a;
17'h2d1c:	data_out=16'h851a;
17'h2d1d:	data_out=16'h885d;
17'h2d1e:	data_out=16'h8787;
17'h2d1f:	data_out=16'h817f;
17'h2d20:	data_out=16'h84d1;
17'h2d21:	data_out=16'h80c0;
17'h2d22:	data_out=16'h802e;
17'h2d23:	data_out=16'h8376;
17'h2d24:	data_out=16'h8377;
17'h2d25:	data_out=16'h402;
17'h2d26:	data_out=16'h89d9;
17'h2d27:	data_out=16'h87ef;
17'h2d28:	data_out=16'h807c;
17'h2d29:	data_out=16'h85e3;
17'h2d2a:	data_out=16'h87f0;
17'h2d2b:	data_out=16'h813f;
17'h2d2c:	data_out=16'h820e;
17'h2d2d:	data_out=16'h54;
17'h2d2e:	data_out=16'h8574;
17'h2d2f:	data_out=16'h80cf;
17'h2d30:	data_out=16'ha00;
17'h2d31:	data_out=16'h8811;
17'h2d32:	data_out=16'ha00;
17'h2d33:	data_out=16'h8885;
17'h2d34:	data_out=16'h8933;
17'h2d35:	data_out=16'h828;
17'h2d36:	data_out=16'h87fa;
17'h2d37:	data_out=16'h8426;
17'h2d38:	data_out=16'h87d9;
17'h2d39:	data_out=16'h88a6;
17'h2d3a:	data_out=16'h8377;
17'h2d3b:	data_out=16'h11b;
17'h2d3c:	data_out=16'h8447;
17'h2d3d:	data_out=16'h8721;
17'h2d3e:	data_out=16'h807e;
17'h2d3f:	data_out=16'h5e1;
17'h2d40:	data_out=16'ha00;
17'h2d41:	data_out=16'h81dd;
17'h2d42:	data_out=16'h5d6;
17'h2d43:	data_out=16'h3f9;
17'h2d44:	data_out=16'h8425;
17'h2d45:	data_out=16'h835a;
17'h2d46:	data_out=16'h836d;
17'h2d47:	data_out=16'h820b;
17'h2d48:	data_out=16'h157;
17'h2d49:	data_out=16'h422;
17'h2d4a:	data_out=16'h626;
17'h2d4b:	data_out=16'h6fd;
17'h2d4c:	data_out=16'h3b4;
17'h2d4d:	data_out=16'h804b;
17'h2d4e:	data_out=16'h8413;
17'h2d4f:	data_out=16'h250;
17'h2d50:	data_out=16'h52a;
17'h2d51:	data_out=16'h8394;
17'h2d52:	data_out=16'h8363;
17'h2d53:	data_out=16'h824a;
17'h2d54:	data_out=16'h85a9;
17'h2d55:	data_out=16'h85cb;
17'h2d56:	data_out=16'h85a1;
17'h2d57:	data_out=16'h84ec;
17'h2d58:	data_out=16'h8693;
17'h2d59:	data_out=16'h4bd;
17'h2d5a:	data_out=16'h80f1;
17'h2d5b:	data_out=16'h884b;
17'h2d5c:	data_out=16'h80ad;
17'h2d5d:	data_out=16'h8250;
17'h2d5e:	data_out=16'h9b;
17'h2d5f:	data_out=16'h82fc;
17'h2d60:	data_out=16'h8a00;
17'h2d61:	data_out=16'h84a0;
17'h2d62:	data_out=16'h831f;
17'h2d63:	data_out=16'h87f9;
17'h2d64:	data_out=16'h896c;
17'h2d65:	data_out=16'h7af;
17'h2d66:	data_out=16'h4ea;
17'h2d67:	data_out=16'h810c;
17'h2d68:	data_out=16'h80a6;
17'h2d69:	data_out=16'h8997;
17'h2d6a:	data_out=16'h8111;
17'h2d6b:	data_out=16'h861;
17'h2d6c:	data_out=16'h8a00;
17'h2d6d:	data_out=16'h8820;
17'h2d6e:	data_out=16'h80fe;
17'h2d6f:	data_out=16'ha00;
17'h2d70:	data_out=16'h80e6;
17'h2d71:	data_out=16'h880a;
17'h2d72:	data_out=16'h188;
17'h2d73:	data_out=16'h1bf;
17'h2d74:	data_out=16'ha00;
17'h2d75:	data_out=16'hcc;
17'h2d76:	data_out=16'h82ae;
17'h2d77:	data_out=16'h5be;
17'h2d78:	data_out=16'h72c;
17'h2d79:	data_out=16'h87dc;
17'h2d7a:	data_out=16'h8719;
17'h2d7b:	data_out=16'h807c;
17'h2d7c:	data_out=16'h8314;
17'h2d7d:	data_out=16'h311;
17'h2d7e:	data_out=16'h81d3;
17'h2d7f:	data_out=16'h276;
17'h2d80:	data_out=16'h8a00;
17'h2d81:	data_out=16'h8a00;
17'h2d82:	data_out=16'h8921;
17'h2d83:	data_out=16'h8046;
17'h2d84:	data_out=16'ha00;
17'h2d85:	data_out=16'ha00;
17'h2d86:	data_out=16'h7fd;
17'h2d87:	data_out=16'h541;
17'h2d88:	data_out=16'h8a00;
17'h2d89:	data_out=16'h381;
17'h2d8a:	data_out=16'h89a6;
17'h2d8b:	data_out=16'h40;
17'h2d8c:	data_out=16'ha00;
17'h2d8d:	data_out=16'h85a0;
17'h2d8e:	data_out=16'h81e9;
17'h2d8f:	data_out=16'h899e;
17'h2d90:	data_out=16'h252;
17'h2d91:	data_out=16'h6ae;
17'h2d92:	data_out=16'h8096;
17'h2d93:	data_out=16'h81c9;
17'h2d94:	data_out=16'h8950;
17'h2d95:	data_out=16'h83db;
17'h2d96:	data_out=16'h8604;
17'h2d97:	data_out=16'h87e5;
17'h2d98:	data_out=16'h859c;
17'h2d99:	data_out=16'h98d;
17'h2d9a:	data_out=16'ha00;
17'h2d9b:	data_out=16'h8084;
17'h2d9c:	data_out=16'h84f3;
17'h2d9d:	data_out=16'h8792;
17'h2d9e:	data_out=16'h89ff;
17'h2d9f:	data_out=16'h99;
17'h2da0:	data_out=16'h8038;
17'h2da1:	data_out=16'h81ac;
17'h2da2:	data_out=16'h58e;
17'h2da3:	data_out=16'h85a4;
17'h2da4:	data_out=16'h85a3;
17'h2da5:	data_out=16'h7ef;
17'h2da6:	data_out=16'h89db;
17'h2da7:	data_out=16'h873f;
17'h2da8:	data_out=16'h8129;
17'h2da9:	data_out=16'h89d4;
17'h2daa:	data_out=16'h8994;
17'h2dab:	data_out=16'h3a6;
17'h2dac:	data_out=16'h8481;
17'h2dad:	data_out=16'h110;
17'h2dae:	data_out=16'h88f1;
17'h2daf:	data_out=16'h33b;
17'h2db0:	data_out=16'ha00;
17'h2db1:	data_out=16'h88a7;
17'h2db2:	data_out=16'ha00;
17'h2db3:	data_out=16'h8a00;
17'h2db4:	data_out=16'h8a00;
17'h2db5:	data_out=16'h947;
17'h2db6:	data_out=16'h8a00;
17'h2db7:	data_out=16'h888e;
17'h2db8:	data_out=16'h8397;
17'h2db9:	data_out=16'h8a00;
17'h2dba:	data_out=16'h27;
17'h2dbb:	data_out=16'h573;
17'h2dbc:	data_out=16'h89a0;
17'h2dbd:	data_out=16'h8395;
17'h2dbe:	data_out=16'h8112;
17'h2dbf:	data_out=16'ha00;
17'h2dc0:	data_out=16'ha00;
17'h2dc1:	data_out=16'h8611;
17'h2dc2:	data_out=16'h650;
17'h2dc3:	data_out=16'h78e;
17'h2dc4:	data_out=16'h83dc;
17'h2dc5:	data_out=16'h83ea;
17'h2dc6:	data_out=16'h85ac;
17'h2dc7:	data_out=16'h80c3;
17'h2dc8:	data_out=16'h52e;
17'h2dc9:	data_out=16'h8f6;
17'h2dca:	data_out=16'h981;
17'h2dcb:	data_out=16'h307;
17'h2dcc:	data_out=16'h271;
17'h2dcd:	data_out=16'h5e6;
17'h2dce:	data_out=16'h8642;
17'h2dcf:	data_out=16'h2a7;
17'h2dd0:	data_out=16'ha00;
17'h2dd1:	data_out=16'h8867;
17'h2dd2:	data_out=16'h8507;
17'h2dd3:	data_out=16'h104;
17'h2dd4:	data_out=16'h8285;
17'h2dd5:	data_out=16'h89ac;
17'h2dd6:	data_out=16'h864e;
17'h2dd7:	data_out=16'h845b;
17'h2dd8:	data_out=16'h8a00;
17'h2dd9:	data_out=16'ha00;
17'h2dda:	data_out=16'h835b;
17'h2ddb:	data_out=16'h8880;
17'h2ddc:	data_out=16'h4b;
17'h2ddd:	data_out=16'h8308;
17'h2dde:	data_out=16'h456;
17'h2ddf:	data_out=16'h8372;
17'h2de0:	data_out=16'h8992;
17'h2de1:	data_out=16'h84d0;
17'h2de2:	data_out=16'h87d9;
17'h2de3:	data_out=16'h89e8;
17'h2de4:	data_out=16'h8990;
17'h2de5:	data_out=16'ha00;
17'h2de6:	data_out=16'h984;
17'h2de7:	data_out=16'h197;
17'h2de8:	data_out=16'h8177;
17'h2de9:	data_out=16'h8a00;
17'h2dea:	data_out=16'h8213;
17'h2deb:	data_out=16'h9e8;
17'h2dec:	data_out=16'h8a00;
17'h2ded:	data_out=16'h8a00;
17'h2dee:	data_out=16'h8212;
17'h2def:	data_out=16'ha00;
17'h2df0:	data_out=16'h8203;
17'h2df1:	data_out=16'h89ce;
17'h2df2:	data_out=16'h3de;
17'h2df3:	data_out=16'h560;
17'h2df4:	data_out=16'ha00;
17'h2df5:	data_out=16'h834f;
17'h2df6:	data_out=16'h34e;
17'h2df7:	data_out=16'ha00;
17'h2df8:	data_out=16'ha00;
17'h2df9:	data_out=16'h8a00;
17'h2dfa:	data_out=16'h8923;
17'h2dfb:	data_out=16'h8111;
17'h2dfc:	data_out=16'h8407;
17'h2dfd:	data_out=16'h7c0;
17'h2dfe:	data_out=16'h3d7;
17'h2dff:	data_out=16'h619;
17'h2e00:	data_out=16'h8a00;
17'h2e01:	data_out=16'h89bd;
17'h2e02:	data_out=16'h8a00;
17'h2e03:	data_out=16'h80fa;
17'h2e04:	data_out=16'ha00;
17'h2e05:	data_out=16'h9fd;
17'h2e06:	data_out=16'h950;
17'h2e07:	data_out=16'ha00;
17'h2e08:	data_out=16'h8a00;
17'h2e09:	data_out=16'h8b1;
17'h2e0a:	data_out=16'h88f2;
17'h2e0b:	data_out=16'h87c7;
17'h2e0c:	data_out=16'ha00;
17'h2e0d:	data_out=16'h8a00;
17'h2e0e:	data_out=16'h81d3;
17'h2e0f:	data_out=16'h89cc;
17'h2e10:	data_out=16'h66e;
17'h2e11:	data_out=16'h6a5;
17'h2e12:	data_out=16'h898d;
17'h2e13:	data_out=16'h861e;
17'h2e14:	data_out=16'h89fe;
17'h2e15:	data_out=16'h8404;
17'h2e16:	data_out=16'h89af;
17'h2e17:	data_out=16'h89ff;
17'h2e18:	data_out=16'h89f8;
17'h2e19:	data_out=16'ha00;
17'h2e1a:	data_out=16'ha00;
17'h2e1b:	data_out=16'h84c7;
17'h2e1c:	data_out=16'h810f;
17'h2e1d:	data_out=16'h83ea;
17'h2e1e:	data_out=16'h89fd;
17'h2e1f:	data_out=16'he9;
17'h2e20:	data_out=16'h9ab;
17'h2e21:	data_out=16'h8199;
17'h2e22:	data_out=16'ha00;
17'h2e23:	data_out=16'h8614;
17'h2e24:	data_out=16'h860f;
17'h2e25:	data_out=16'ha00;
17'h2e26:	data_out=16'h89ff;
17'h2e27:	data_out=16'h82bc;
17'h2e28:	data_out=16'h809f;
17'h2e29:	data_out=16'h89ff;
17'h2e2a:	data_out=16'h8968;
17'h2e2b:	data_out=16'h9fc;
17'h2e2c:	data_out=16'h885c;
17'h2e2d:	data_out=16'h2a4;
17'h2e2e:	data_out=16'h88ff;
17'h2e2f:	data_out=16'h9f0;
17'h2e30:	data_out=16'ha00;
17'h2e31:	data_out=16'h85ae;
17'h2e32:	data_out=16'ha00;
17'h2e33:	data_out=16'h8a00;
17'h2e34:	data_out=16'h868a;
17'h2e35:	data_out=16'h9c1;
17'h2e36:	data_out=16'h89fe;
17'h2e37:	data_out=16'h8a00;
17'h2e38:	data_out=16'h9d9;
17'h2e39:	data_out=16'h8a00;
17'h2e3a:	data_out=16'h4b6;
17'h2e3b:	data_out=16'ha00;
17'h2e3c:	data_out=16'h8a00;
17'h2e3d:	data_out=16'h439;
17'h2e3e:	data_out=16'h8099;
17'h2e3f:	data_out=16'h9fd;
17'h2e40:	data_out=16'ha00;
17'h2e41:	data_out=16'h8a00;
17'h2e42:	data_out=16'h8b9;
17'h2e43:	data_out=16'ha00;
17'h2e44:	data_out=16'h8228;
17'h2e45:	data_out=16'h842d;
17'h2e46:	data_out=16'h875d;
17'h2e47:	data_out=16'h80cd;
17'h2e48:	data_out=16'h6f2;
17'h2e49:	data_out=16'ha00;
17'h2e4a:	data_out=16'ha00;
17'h2e4b:	data_out=16'h69f;
17'h2e4c:	data_out=16'h2b;
17'h2e4d:	data_out=16'ha00;
17'h2e4e:	data_out=16'h878e;
17'h2e4f:	data_out=16'h2f0;
17'h2e50:	data_out=16'ha00;
17'h2e51:	data_out=16'h8a00;
17'h2e52:	data_out=16'h84cb;
17'h2e53:	data_out=16'h60c;
17'h2e54:	data_out=16'h6c9;
17'h2e55:	data_out=16'h89fc;
17'h2e56:	data_out=16'h8a00;
17'h2e57:	data_out=16'h8703;
17'h2e58:	data_out=16'h8a00;
17'h2e59:	data_out=16'ha00;
17'h2e5a:	data_out=16'h8a00;
17'h2e5b:	data_out=16'h8504;
17'h2e5c:	data_out=16'h342;
17'h2e5d:	data_out=16'h839f;
17'h2e5e:	data_out=16'h9f5;
17'h2e5f:	data_out=16'h84a8;
17'h2e60:	data_out=16'h89dc;
17'h2e61:	data_out=16'hfc;
17'h2e62:	data_out=16'h88d3;
17'h2e63:	data_out=16'h8a00;
17'h2e64:	data_out=16'h877a;
17'h2e65:	data_out=16'ha00;
17'h2e66:	data_out=16'ha00;
17'h2e67:	data_out=16'h2d6;
17'h2e68:	data_out=16'h814c;
17'h2e69:	data_out=16'h8a00;
17'h2e6a:	data_out=16'h81f9;
17'h2e6b:	data_out=16'h9fe;
17'h2e6c:	data_out=16'h89ff;
17'h2e6d:	data_out=16'h89ff;
17'h2e6e:	data_out=16'h81f8;
17'h2e6f:	data_out=16'ha00;
17'h2e70:	data_out=16'h81e5;
17'h2e71:	data_out=16'h89fe;
17'h2e72:	data_out=16'ha00;
17'h2e73:	data_out=16'h9fd;
17'h2e74:	data_out=16'ha00;
17'h2e75:	data_out=16'h89f8;
17'h2e76:	data_out=16'h9ff;
17'h2e77:	data_out=16'ha00;
17'h2e78:	data_out=16'ha00;
17'h2e79:	data_out=16'h8a00;
17'h2e7a:	data_out=16'h89fb;
17'h2e7b:	data_out=16'h807e;
17'h2e7c:	data_out=16'h8680;
17'h2e7d:	data_out=16'h9fe;
17'h2e7e:	data_out=16'h77e;
17'h2e7f:	data_out=16'ha00;
17'h2e80:	data_out=16'h89f0;
17'h2e81:	data_out=16'h84b7;
17'h2e82:	data_out=16'h8991;
17'h2e83:	data_out=16'h9fd;
17'h2e84:	data_out=16'ha00;
17'h2e85:	data_out=16'ha00;
17'h2e86:	data_out=16'h9fe;
17'h2e87:	data_out=16'h9f1;
17'h2e88:	data_out=16'h89fd;
17'h2e89:	data_out=16'ha00;
17'h2e8a:	data_out=16'h8514;
17'h2e8b:	data_out=16'h859c;
17'h2e8c:	data_out=16'h9fc;
17'h2e8d:	data_out=16'h8a00;
17'h2e8e:	data_out=16'h804e;
17'h2e8f:	data_out=16'h882b;
17'h2e90:	data_out=16'ha00;
17'h2e91:	data_out=16'h765;
17'h2e92:	data_out=16'h8a00;
17'h2e93:	data_out=16'h9ff;
17'h2e94:	data_out=16'h8835;
17'h2e95:	data_out=16'h400;
17'h2e96:	data_out=16'h859c;
17'h2e97:	data_out=16'h88b4;
17'h2e98:	data_out=16'h8a00;
17'h2e99:	data_out=16'ha00;
17'h2e9a:	data_out=16'ha00;
17'h2e9b:	data_out=16'h3be;
17'h2e9c:	data_out=16'h99d;
17'h2e9d:	data_out=16'h51b;
17'h2e9e:	data_out=16'h8737;
17'h2e9f:	data_out=16'h6b5;
17'h2ea0:	data_out=16'h9ff;
17'h2ea1:	data_out=16'ha;
17'h2ea2:	data_out=16'ha00;
17'h2ea3:	data_out=16'h89c5;
17'h2ea4:	data_out=16'h89c4;
17'h2ea5:	data_out=16'ha00;
17'h2ea6:	data_out=16'h89fb;
17'h2ea7:	data_out=16'h6e2;
17'h2ea8:	data_out=16'h1b3;
17'h2ea9:	data_out=16'h89b8;
17'h2eaa:	data_out=16'h8686;
17'h2eab:	data_out=16'ha00;
17'h2eac:	data_out=16'h80dc;
17'h2ead:	data_out=16'h6a7;
17'h2eae:	data_out=16'h86d8;
17'h2eaf:	data_out=16'ha00;
17'h2eb0:	data_out=16'ha00;
17'h2eb1:	data_out=16'hfe;
17'h2eb2:	data_out=16'ha00;
17'h2eb3:	data_out=16'h883c;
17'h2eb4:	data_out=16'h8388;
17'h2eb5:	data_out=16'h9df;
17'h2eb6:	data_out=16'h8833;
17'h2eb7:	data_out=16'h891f;
17'h2eb8:	data_out=16'h9fe;
17'h2eb9:	data_out=16'h8877;
17'h2eba:	data_out=16'ha00;
17'h2ebb:	data_out=16'ha00;
17'h2ebc:	data_out=16'h865d;
17'h2ebd:	data_out=16'h9ff;
17'h2ebe:	data_out=16'h1d2;
17'h2ebf:	data_out=16'ha00;
17'h2ec0:	data_out=16'ha00;
17'h2ec1:	data_out=16'h8507;
17'h2ec2:	data_out=16'h9fc;
17'h2ec3:	data_out=16'ha00;
17'h2ec4:	data_out=16'h776;
17'h2ec5:	data_out=16'h3f1;
17'h2ec6:	data_out=16'h8389;
17'h2ec7:	data_out=16'h7ac;
17'h2ec8:	data_out=16'ha00;
17'h2ec9:	data_out=16'ha00;
17'h2eca:	data_out=16'h9fc;
17'h2ecb:	data_out=16'ha00;
17'h2ecc:	data_out=16'h582;
17'h2ecd:	data_out=16'ha00;
17'h2ece:	data_out=16'h837b;
17'h2ecf:	data_out=16'ha00;
17'h2ed0:	data_out=16'ha00;
17'h2ed1:	data_out=16'h8a00;
17'h2ed2:	data_out=16'h8711;
17'h2ed3:	data_out=16'h9fa;
17'h2ed4:	data_out=16'h9ff;
17'h2ed5:	data_out=16'h88b0;
17'h2ed6:	data_out=16'h2a6;
17'h2ed7:	data_out=16'h79e;
17'h2ed8:	data_out=16'h8a00;
17'h2ed9:	data_out=16'ha00;
17'h2eda:	data_out=16'h8914;
17'h2edb:	data_out=16'h90f;
17'h2edc:	data_out=16'h97e;
17'h2edd:	data_out=16'h90a;
17'h2ede:	data_out=16'ha00;
17'h2edf:	data_out=16'h82c1;
17'h2ee0:	data_out=16'h89fa;
17'h2ee1:	data_out=16'ha00;
17'h2ee2:	data_out=16'h8594;
17'h2ee3:	data_out=16'h87f1;
17'h2ee4:	data_out=16'h83d0;
17'h2ee5:	data_out=16'ha00;
17'h2ee6:	data_out=16'ha00;
17'h2ee7:	data_out=16'h9ff;
17'h2ee8:	data_out=16'haa;
17'h2ee9:	data_out=16'h8a00;
17'h2eea:	data_out=16'h806f;
17'h2eeb:	data_out=16'ha00;
17'h2eec:	data_out=16'h89f0;
17'h2eed:	data_out=16'h87d9;
17'h2eee:	data_out=16'h806f;
17'h2eef:	data_out=16'ha00;
17'h2ef0:	data_out=16'h8060;
17'h2ef1:	data_out=16'h8988;
17'h2ef2:	data_out=16'ha00;
17'h2ef3:	data_out=16'ha00;
17'h2ef4:	data_out=16'h9fc;
17'h2ef5:	data_out=16'h89ee;
17'h2ef6:	data_out=16'ha00;
17'h2ef7:	data_out=16'ha00;
17'h2ef8:	data_out=16'ha00;
17'h2ef9:	data_out=16'h86ce;
17'h2efa:	data_out=16'h87e2;
17'h2efb:	data_out=16'h208;
17'h2efc:	data_out=16'h87f4;
17'h2efd:	data_out=16'ha00;
17'h2efe:	data_out=16'h9f9;
17'h2eff:	data_out=16'ha00;
17'h2f00:	data_out=16'h89f3;
17'h2f01:	data_out=16'h18d;
17'h2f02:	data_out=16'h89fb;
17'h2f03:	data_out=16'h9fc;
17'h2f04:	data_out=16'ha00;
17'h2f05:	data_out=16'ha00;
17'h2f06:	data_out=16'h9fd;
17'h2f07:	data_out=16'h9ff;
17'h2f08:	data_out=16'h89f8;
17'h2f09:	data_out=16'ha00;
17'h2f0a:	data_out=16'h81e8;
17'h2f0b:	data_out=16'h8537;
17'h2f0c:	data_out=16'ha00;
17'h2f0d:	data_out=16'h8a00;
17'h2f0e:	data_out=16'h81df;
17'h2f0f:	data_out=16'h88c3;
17'h2f10:	data_out=16'ha00;
17'h2f11:	data_out=16'h7b8;
17'h2f12:	data_out=16'h8a00;
17'h2f13:	data_out=16'h59a;
17'h2f14:	data_out=16'h88bb;
17'h2f15:	data_out=16'h3c2;
17'h2f16:	data_out=16'h859f;
17'h2f17:	data_out=16'h89a8;
17'h2f18:	data_out=16'h8a00;
17'h2f19:	data_out=16'ha00;
17'h2f1a:	data_out=16'ha00;
17'h2f1b:	data_out=16'h4a;
17'h2f1c:	data_out=16'h958;
17'h2f1d:	data_out=16'h9e0;
17'h2f1e:	data_out=16'h86bf;
17'h2f1f:	data_out=16'h2b1;
17'h2f20:	data_out=16'ha00;
17'h2f21:	data_out=16'h80d4;
17'h2f22:	data_out=16'ha00;
17'h2f23:	data_out=16'h88b4;
17'h2f24:	data_out=16'h88ad;
17'h2f25:	data_out=16'ha00;
17'h2f26:	data_out=16'h89f6;
17'h2f27:	data_out=16'h9ec;
17'h2f28:	data_out=16'hec;
17'h2f29:	data_out=16'h89fa;
17'h2f2a:	data_out=16'h861d;
17'h2f2b:	data_out=16'h9fd;
17'h2f2c:	data_out=16'h8492;
17'h2f2d:	data_out=16'h8141;
17'h2f2e:	data_out=16'h87a0;
17'h2f2f:	data_out=16'ha00;
17'h2f30:	data_out=16'ha00;
17'h2f31:	data_out=16'h8b6;
17'h2f32:	data_out=16'ha00;
17'h2f33:	data_out=16'h884d;
17'h2f34:	data_out=16'h82f1;
17'h2f35:	data_out=16'h9f3;
17'h2f36:	data_out=16'h8730;
17'h2f37:	data_out=16'h8992;
17'h2f38:	data_out=16'h9f8;
17'h2f39:	data_out=16'h888a;
17'h2f3a:	data_out=16'h874;
17'h2f3b:	data_out=16'ha00;
17'h2f3c:	data_out=16'h85e8;
17'h2f3d:	data_out=16'ha00;
17'h2f3e:	data_out=16'hef;
17'h2f3f:	data_out=16'ha00;
17'h2f40:	data_out=16'ha00;
17'h2f41:	data_out=16'h825a;
17'h2f42:	data_out=16'ha00;
17'h2f43:	data_out=16'ha00;
17'h2f44:	data_out=16'h9d4;
17'h2f45:	data_out=16'h39a;
17'h2f46:	data_out=16'h87ba;
17'h2f47:	data_out=16'h191;
17'h2f48:	data_out=16'ha00;
17'h2f49:	data_out=16'ha00;
17'h2f4a:	data_out=16'ha00;
17'h2f4b:	data_out=16'ha00;
17'h2f4c:	data_out=16'h6a2;
17'h2f4d:	data_out=16'ha00;
17'h2f4e:	data_out=16'h82dc;
17'h2f4f:	data_out=16'ha00;
17'h2f50:	data_out=16'ha00;
17'h2f51:	data_out=16'h8a00;
17'h2f52:	data_out=16'h85b5;
17'h2f53:	data_out=16'h9f4;
17'h2f54:	data_out=16'ha00;
17'h2f55:	data_out=16'h8991;
17'h2f56:	data_out=16'h85ec;
17'h2f57:	data_out=16'h813a;
17'h2f58:	data_out=16'h89ff;
17'h2f59:	data_out=16'ha00;
17'h2f5a:	data_out=16'h87db;
17'h2f5b:	data_out=16'ha00;
17'h2f5c:	data_out=16'h946;
17'h2f5d:	data_out=16'ha00;
17'h2f5e:	data_out=16'ha00;
17'h2f5f:	data_out=16'h84f7;
17'h2f60:	data_out=16'h89f3;
17'h2f61:	data_out=16'ha00;
17'h2f62:	data_out=16'h8569;
17'h2f63:	data_out=16'h87c2;
17'h2f64:	data_out=16'h809a;
17'h2f65:	data_out=16'ha00;
17'h2f66:	data_out=16'ha00;
17'h2f67:	data_out=16'ha00;
17'h2f68:	data_out=16'h16;
17'h2f69:	data_out=16'h89fe;
17'h2f6a:	data_out=16'h8254;
17'h2f6b:	data_out=16'ha00;
17'h2f6c:	data_out=16'h89ee;
17'h2f6d:	data_out=16'h87a0;
17'h2f6e:	data_out=16'h8253;
17'h2f6f:	data_out=16'ha00;
17'h2f70:	data_out=16'h8231;
17'h2f71:	data_out=16'h89fa;
17'h2f72:	data_out=16'ha00;
17'h2f73:	data_out=16'ha00;
17'h2f74:	data_out=16'ha00;
17'h2f75:	data_out=16'h88bf;
17'h2f76:	data_out=16'ha00;
17'h2f77:	data_out=16'ha00;
17'h2f78:	data_out=16'ha00;
17'h2f79:	data_out=16'h87a0;
17'h2f7a:	data_out=16'h87be;
17'h2f7b:	data_out=16'hed;
17'h2f7c:	data_out=16'h8a00;
17'h2f7d:	data_out=16'ha00;
17'h2f7e:	data_out=16'h995;
17'h2f7f:	data_out=16'ha00;
17'h2f80:	data_out=16'h8a00;
17'h2f81:	data_out=16'h34e;
17'h2f82:	data_out=16'h89ff;
17'h2f83:	data_out=16'h720;
17'h2f84:	data_out=16'ha00;
17'h2f85:	data_out=16'ha00;
17'h2f86:	data_out=16'ha00;
17'h2f87:	data_out=16'ha00;
17'h2f88:	data_out=16'h89fe;
17'h2f89:	data_out=16'h986;
17'h2f8a:	data_out=16'h8037;
17'h2f8b:	data_out=16'h8017;
17'h2f8c:	data_out=16'ha00;
17'h2f8d:	data_out=16'h8a00;
17'h2f8e:	data_out=16'h864c;
17'h2f8f:	data_out=16'h89ff;
17'h2f90:	data_out=16'ha00;
17'h2f91:	data_out=16'h54c;
17'h2f92:	data_out=16'h8a00;
17'h2f93:	data_out=16'h11;
17'h2f94:	data_out=16'h89f7;
17'h2f95:	data_out=16'h85c3;
17'h2f96:	data_out=16'h87f1;
17'h2f97:	data_out=16'h89fa;
17'h2f98:	data_out=16'h8a00;
17'h2f99:	data_out=16'ha00;
17'h2f9a:	data_out=16'ha00;
17'h2f9b:	data_out=16'h29a;
17'h2f9c:	data_out=16'h774;
17'h2f9d:	data_out=16'h8f6;
17'h2f9e:	data_out=16'h89b8;
17'h2f9f:	data_out=16'h8863;
17'h2fa0:	data_out=16'h9fd;
17'h2fa1:	data_out=16'h84a6;
17'h2fa2:	data_out=16'ha00;
17'h2fa3:	data_out=16'h8790;
17'h2fa4:	data_out=16'h8787;
17'h2fa5:	data_out=16'h9ff;
17'h2fa6:	data_out=16'h8a00;
17'h2fa7:	data_out=16'h9df;
17'h2fa8:	data_out=16'h82cf;
17'h2fa9:	data_out=16'h89ff;
17'h2faa:	data_out=16'h887e;
17'h2fab:	data_out=16'ha00;
17'h2fac:	data_out=16'h87c3;
17'h2fad:	data_out=16'h8866;
17'h2fae:	data_out=16'h8907;
17'h2faf:	data_out=16'ha00;
17'h2fb0:	data_out=16'ha00;
17'h2fb1:	data_out=16'h687;
17'h2fb2:	data_out=16'ha00;
17'h2fb3:	data_out=16'h89fa;
17'h2fb4:	data_out=16'h88a3;
17'h2fb5:	data_out=16'h9e2;
17'h2fb6:	data_out=16'h8924;
17'h2fb7:	data_out=16'h89ff;
17'h2fb8:	data_out=16'h9e1;
17'h2fb9:	data_out=16'h89fc;
17'h2fba:	data_out=16'h686;
17'h2fbb:	data_out=16'ha00;
17'h2fbc:	data_out=16'h84f6;
17'h2fbd:	data_out=16'h9f2;
17'h2fbe:	data_out=16'h82c6;
17'h2fbf:	data_out=16'ha00;
17'h2fc0:	data_out=16'ha00;
17'h2fc1:	data_out=16'h23;
17'h2fc2:	data_out=16'h9ff;
17'h2fc3:	data_out=16'ha00;
17'h2fc4:	data_out=16'h914;
17'h2fc5:	data_out=16'h8612;
17'h2fc6:	data_out=16'h84d3;
17'h2fc7:	data_out=16'h894a;
17'h2fc8:	data_out=16'ha00;
17'h2fc9:	data_out=16'ha00;
17'h2fca:	data_out=16'ha00;
17'h2fcb:	data_out=16'h9ff;
17'h2fcc:	data_out=16'h106;
17'h2fcd:	data_out=16'ha00;
17'h2fce:	data_out=16'h81e7;
17'h2fcf:	data_out=16'h4f2;
17'h2fd0:	data_out=16'ha00;
17'h2fd1:	data_out=16'h8a00;
17'h2fd2:	data_out=16'h8577;
17'h2fd3:	data_out=16'h9f9;
17'h2fd4:	data_out=16'h9fc;
17'h2fd5:	data_out=16'h8a00;
17'h2fd6:	data_out=16'h89ff;
17'h2fd7:	data_out=16'h89ff;
17'h2fd8:	data_out=16'h8a00;
17'h2fd9:	data_out=16'ha00;
17'h2fda:	data_out=16'h803a;
17'h2fdb:	data_out=16'h9ec;
17'h2fdc:	data_out=16'h8e8;
17'h2fdd:	data_out=16'h8de;
17'h2fde:	data_out=16'ha00;
17'h2fdf:	data_out=16'h88df;
17'h2fe0:	data_out=16'h89ff;
17'h2fe1:	data_out=16'ha00;
17'h2fe2:	data_out=16'h86a7;
17'h2fe3:	data_out=16'h897c;
17'h2fe4:	data_out=16'h82ab;
17'h2fe5:	data_out=16'ha00;
17'h2fe6:	data_out=16'ha00;
17'h2fe7:	data_out=16'h9ff;
17'h2fe8:	data_out=16'h83c4;
17'h2fe9:	data_out=16'h8a00;
17'h2fea:	data_out=16'h8753;
17'h2feb:	data_out=16'ha00;
17'h2fec:	data_out=16'h8a00;
17'h2fed:	data_out=16'h897f;
17'h2fee:	data_out=16'h8751;
17'h2fef:	data_out=16'ha00;
17'h2ff0:	data_out=16'h86c3;
17'h2ff1:	data_out=16'h89ff;
17'h2ff2:	data_out=16'ha00;
17'h2ff3:	data_out=16'ha00;
17'h2ff4:	data_out=16'ha00;
17'h2ff5:	data_out=16'h154;
17'h2ff6:	data_out=16'ha00;
17'h2ff7:	data_out=16'h9ff;
17'h2ff8:	data_out=16'ha00;
17'h2ff9:	data_out=16'h8a00;
17'h2ffa:	data_out=16'h8980;
17'h2ffb:	data_out=16'h82c3;
17'h2ffc:	data_out=16'h8a00;
17'h2ffd:	data_out=16'ha00;
17'h2ffe:	data_out=16'h91a;
17'h2fff:	data_out=16'ha00;
17'h3000:	data_out=16'h8a00;
17'h3001:	data_out=16'h963;
17'h3002:	data_out=16'h8a00;
17'h3003:	data_out=16'h95f;
17'h3004:	data_out=16'ha00;
17'h3005:	data_out=16'ha00;
17'h3006:	data_out=16'h9ff;
17'h3007:	data_out=16'h9ff;
17'h3008:	data_out=16'h89ff;
17'h3009:	data_out=16'h36;
17'h300a:	data_out=16'h9ea;
17'h300b:	data_out=16'h21c;
17'h300c:	data_out=16'ha00;
17'h300d:	data_out=16'h8a00;
17'h300e:	data_out=16'h8654;
17'h300f:	data_out=16'h8a00;
17'h3010:	data_out=16'ha00;
17'h3011:	data_out=16'h4c8;
17'h3012:	data_out=16'h8a00;
17'h3013:	data_out=16'h977;
17'h3014:	data_out=16'h8952;
17'h3015:	data_out=16'h4d7;
17'h3016:	data_out=16'h8426;
17'h3017:	data_out=16'h8975;
17'h3018:	data_out=16'h8a00;
17'h3019:	data_out=16'ha00;
17'h301a:	data_out=16'ha00;
17'h301b:	data_out=16'h254;
17'h301c:	data_out=16'h8c2;
17'h301d:	data_out=16'h918;
17'h301e:	data_out=16'h8971;
17'h301f:	data_out=16'h87a4;
17'h3020:	data_out=16'h9fd;
17'h3021:	data_out=16'h855c;
17'h3022:	data_out=16'h5c6;
17'h3023:	data_out=16'h89a5;
17'h3024:	data_out=16'h8995;
17'h3025:	data_out=16'h9fe;
17'h3026:	data_out=16'h8a00;
17'h3027:	data_out=16'h9d9;
17'h3028:	data_out=16'h8391;
17'h3029:	data_out=16'h8a00;
17'h302a:	data_out=16'h89fc;
17'h302b:	data_out=16'h9ff;
17'h302c:	data_out=16'h17a;
17'h302d:	data_out=16'h8a00;
17'h302e:	data_out=16'h89f0;
17'h302f:	data_out=16'ha00;
17'h3030:	data_out=16'ha00;
17'h3031:	data_out=16'h87e;
17'h3032:	data_out=16'ha00;
17'h3033:	data_out=16'h88d5;
17'h3034:	data_out=16'h8336;
17'h3035:	data_out=16'h9e0;
17'h3036:	data_out=16'h89ce;
17'h3037:	data_out=16'h8a00;
17'h3038:	data_out=16'h9d2;
17'h3039:	data_out=16'h894f;
17'h303a:	data_out=16'h8116;
17'h303b:	data_out=16'ha00;
17'h303c:	data_out=16'h211;
17'h303d:	data_out=16'h9e9;
17'h303e:	data_out=16'h8385;
17'h303f:	data_out=16'ha00;
17'h3040:	data_out=16'ha00;
17'h3041:	data_out=16'h442;
17'h3042:	data_out=16'h9bf;
17'h3043:	data_out=16'ha00;
17'h3044:	data_out=16'h9c9;
17'h3045:	data_out=16'h4e0;
17'h3046:	data_out=16'h8a00;
17'h3047:	data_out=16'h89fc;
17'h3048:	data_out=16'h9ff;
17'h3049:	data_out=16'h9fd;
17'h304a:	data_out=16'ha00;
17'h304b:	data_out=16'h9fc;
17'h304c:	data_out=16'h89c6;
17'h304d:	data_out=16'ha00;
17'h304e:	data_out=16'h83f7;
17'h304f:	data_out=16'h88c7;
17'h3050:	data_out=16'ha00;
17'h3051:	data_out=16'h8a00;
17'h3052:	data_out=16'h8843;
17'h3053:	data_out=16'ha00;
17'h3054:	data_out=16'h9fe;
17'h3055:	data_out=16'h8a00;
17'h3056:	data_out=16'h8a00;
17'h3057:	data_out=16'h89ff;
17'h3058:	data_out=16'h8a00;
17'h3059:	data_out=16'ha00;
17'h305a:	data_out=16'h8069;
17'h305b:	data_out=16'h9f2;
17'h305c:	data_out=16'h9db;
17'h305d:	data_out=16'ha00;
17'h305e:	data_out=16'ha00;
17'h305f:	data_out=16'h8909;
17'h3060:	data_out=16'h8a00;
17'h3061:	data_out=16'ha00;
17'h3062:	data_out=16'h879c;
17'h3063:	data_out=16'h87e5;
17'h3064:	data_out=16'h8096;
17'h3065:	data_out=16'ha00;
17'h3066:	data_out=16'ha00;
17'h3067:	data_out=16'ha00;
17'h3068:	data_out=16'h84b3;
17'h3069:	data_out=16'h8a00;
17'h306a:	data_out=16'h88ad;
17'h306b:	data_out=16'ha00;
17'h306c:	data_out=16'h8a00;
17'h306d:	data_out=16'h87fa;
17'h306e:	data_out=16'h88aa;
17'h306f:	data_out=16'ha00;
17'h3070:	data_out=16'h86b8;
17'h3071:	data_out=16'h8a00;
17'h3072:	data_out=16'ha00;
17'h3073:	data_out=16'ha00;
17'h3074:	data_out=16'ha00;
17'h3075:	data_out=16'h9f6;
17'h3076:	data_out=16'ha00;
17'h3077:	data_out=16'h9fd;
17'h3078:	data_out=16'ha00;
17'h3079:	data_out=16'h8a00;
17'h307a:	data_out=16'h884e;
17'h307b:	data_out=16'h8382;
17'h307c:	data_out=16'h8a00;
17'h307d:	data_out=16'ha00;
17'h307e:	data_out=16'h81f7;
17'h307f:	data_out=16'ha00;
17'h3080:	data_out=16'h89ff;
17'h3081:	data_out=16'h943;
17'h3082:	data_out=16'h8a00;
17'h3083:	data_out=16'h94c;
17'h3084:	data_out=16'ha00;
17'h3085:	data_out=16'ha00;
17'h3086:	data_out=16'h9ff;
17'h3087:	data_out=16'h9fe;
17'h3088:	data_out=16'h8a00;
17'h3089:	data_out=16'hbf;
17'h308a:	data_out=16'h9fb;
17'h308b:	data_out=16'h77;
17'h308c:	data_out=16'h9fe;
17'h308d:	data_out=16'h8a00;
17'h308e:	data_out=16'h88a5;
17'h308f:	data_out=16'h8a00;
17'h3090:	data_out=16'ha00;
17'h3091:	data_out=16'h468;
17'h3092:	data_out=16'h8a00;
17'h3093:	data_out=16'h95c;
17'h3094:	data_out=16'h8912;
17'h3095:	data_out=16'h9f6;
17'h3096:	data_out=16'h9e9;
17'h3097:	data_out=16'h86d4;
17'h3098:	data_out=16'h8a00;
17'h3099:	data_out=16'ha00;
17'h309a:	data_out=16'ha00;
17'h309b:	data_out=16'h84b2;
17'h309c:	data_out=16'h802;
17'h309d:	data_out=16'h926;
17'h309e:	data_out=16'h896f;
17'h309f:	data_out=16'h859a;
17'h30a0:	data_out=16'ha00;
17'h30a1:	data_out=16'h8784;
17'h30a2:	data_out=16'h7cf;
17'h30a3:	data_out=16'h89ce;
17'h30a4:	data_out=16'h89ce;
17'h30a5:	data_out=16'h93f;
17'h30a6:	data_out=16'h8a00;
17'h30a7:	data_out=16'h9f2;
17'h30a8:	data_out=16'h85a3;
17'h30a9:	data_out=16'h8a00;
17'h30aa:	data_out=16'h89fc;
17'h30ab:	data_out=16'h9fb;
17'h30ac:	data_out=16'h9f4;
17'h30ad:	data_out=16'h8a00;
17'h30ae:	data_out=16'h89ee;
17'h30af:	data_out=16'ha00;
17'h30b0:	data_out=16'ha00;
17'h30b1:	data_out=16'h872;
17'h30b2:	data_out=16'ha00;
17'h30b3:	data_out=16'h88bd;
17'h30b4:	data_out=16'h354;
17'h30b5:	data_out=16'h9eb;
17'h30b6:	data_out=16'h89fe;
17'h30b7:	data_out=16'h8a00;
17'h30b8:	data_out=16'h950;
17'h30b9:	data_out=16'h8994;
17'h30ba:	data_out=16'h807d;
17'h30bb:	data_out=16'ha00;
17'h30bc:	data_out=16'h314;
17'h30bd:	data_out=16'h9f0;
17'h30be:	data_out=16'h8597;
17'h30bf:	data_out=16'ha00;
17'h30c0:	data_out=16'ha00;
17'h30c1:	data_out=16'h603;
17'h30c2:	data_out=16'h8d7;
17'h30c3:	data_out=16'ha00;
17'h30c4:	data_out=16'h9d2;
17'h30c5:	data_out=16'h9f5;
17'h30c6:	data_out=16'h8a00;
17'h30c7:	data_out=16'h89e7;
17'h30c8:	data_out=16'h9ff;
17'h30c9:	data_out=16'h9fe;
17'h30ca:	data_out=16'ha00;
17'h30cb:	data_out=16'h9fb;
17'h30cc:	data_out=16'h89d6;
17'h30cd:	data_out=16'ha00;
17'h30ce:	data_out=16'h8529;
17'h30cf:	data_out=16'h8893;
17'h30d0:	data_out=16'ha00;
17'h30d1:	data_out=16'h8a00;
17'h30d2:	data_out=16'h882c;
17'h30d3:	data_out=16'ha00;
17'h30d4:	data_out=16'ha00;
17'h30d5:	data_out=16'h8a00;
17'h30d6:	data_out=16'h8a00;
17'h30d7:	data_out=16'h89fe;
17'h30d8:	data_out=16'h8a00;
17'h30d9:	data_out=16'ha00;
17'h30da:	data_out=16'h8a00;
17'h30db:	data_out=16'ha00;
17'h30dc:	data_out=16'h9b0;
17'h30dd:	data_out=16'ha00;
17'h30de:	data_out=16'ha00;
17'h30df:	data_out=16'h88c7;
17'h30e0:	data_out=16'h8a00;
17'h30e1:	data_out=16'ha00;
17'h30e2:	data_out=16'h8620;
17'h30e3:	data_out=16'h86c6;
17'h30e4:	data_out=16'h866d;
17'h30e5:	data_out=16'ha00;
17'h30e6:	data_out=16'ha00;
17'h30e7:	data_out=16'ha00;
17'h30e8:	data_out=16'h86c1;
17'h30e9:	data_out=16'h8a00;
17'h30ea:	data_out=16'h8971;
17'h30eb:	data_out=16'ha00;
17'h30ec:	data_out=16'h89ff;
17'h30ed:	data_out=16'h8711;
17'h30ee:	data_out=16'h896e;
17'h30ef:	data_out=16'ha00;
17'h30f0:	data_out=16'h890a;
17'h30f1:	data_out=16'h8a00;
17'h30f2:	data_out=16'ha00;
17'h30f3:	data_out=16'ha00;
17'h30f4:	data_out=16'ha00;
17'h30f5:	data_out=16'h9cc;
17'h30f6:	data_out=16'ha00;
17'h30f7:	data_out=16'h9fd;
17'h30f8:	data_out=16'ha00;
17'h30f9:	data_out=16'h8a00;
17'h30fa:	data_out=16'h8767;
17'h30fb:	data_out=16'h8593;
17'h30fc:	data_out=16'h8a00;
17'h30fd:	data_out=16'ha00;
17'h30fe:	data_out=16'hc3;
17'h30ff:	data_out=16'ha00;
17'h3100:	data_out=16'h8a00;
17'h3101:	data_out=16'h729;
17'h3102:	data_out=16'h8a00;
17'h3103:	data_out=16'h8e7;
17'h3104:	data_out=16'ha00;
17'h3105:	data_out=16'ha00;
17'h3106:	data_out=16'h9ff;
17'h3107:	data_out=16'h9ff;
17'h3108:	data_out=16'h8a00;
17'h3109:	data_out=16'h82ff;
17'h310a:	data_out=16'h9fb;
17'h310b:	data_out=16'h16d;
17'h310c:	data_out=16'h9fe;
17'h310d:	data_out=16'h88c4;
17'h310e:	data_out=16'h8a00;
17'h310f:	data_out=16'h8a00;
17'h3110:	data_out=16'ha00;
17'h3111:	data_out=16'h275;
17'h3112:	data_out=16'h8a00;
17'h3113:	data_out=16'h9b7;
17'h3114:	data_out=16'h87bc;
17'h3115:	data_out=16'h9f6;
17'h3116:	data_out=16'h9e9;
17'h3117:	data_out=16'h456;
17'h3118:	data_out=16'h8a00;
17'h3119:	data_out=16'ha00;
17'h311a:	data_out=16'ha00;
17'h311b:	data_out=16'h2d3;
17'h311c:	data_out=16'h82f;
17'h311d:	data_out=16'h7ad;
17'h311e:	data_out=16'h8a00;
17'h311f:	data_out=16'h80df;
17'h3120:	data_out=16'ha00;
17'h3121:	data_out=16'h8999;
17'h3122:	data_out=16'h8458;
17'h3123:	data_out=16'h89c6;
17'h3124:	data_out=16'h89c5;
17'h3125:	data_out=16'h873c;
17'h3126:	data_out=16'h8a00;
17'h3127:	data_out=16'ha00;
17'h3128:	data_out=16'h875e;
17'h3129:	data_out=16'h8a00;
17'h312a:	data_out=16'h8a00;
17'h312b:	data_out=16'h9fb;
17'h312c:	data_out=16'h9f3;
17'h312d:	data_out=16'h8a00;
17'h312e:	data_out=16'h89f3;
17'h312f:	data_out=16'ha00;
17'h3130:	data_out=16'ha00;
17'h3131:	data_out=16'h982;
17'h3132:	data_out=16'ha00;
17'h3133:	data_out=16'h8801;
17'h3134:	data_out=16'h8495;
17'h3135:	data_out=16'h9fe;
17'h3136:	data_out=16'h89ff;
17'h3137:	data_out=16'h8a00;
17'h3138:	data_out=16'h8322;
17'h3139:	data_out=16'h89c8;
17'h313a:	data_out=16'h8452;
17'h313b:	data_out=16'ha00;
17'h313c:	data_out=16'h467;
17'h313d:	data_out=16'h9e7;
17'h313e:	data_out=16'h8750;
17'h313f:	data_out=16'ha00;
17'h3140:	data_out=16'ha00;
17'h3141:	data_out=16'h784;
17'h3142:	data_out=16'hce;
17'h3143:	data_out=16'ha00;
17'h3144:	data_out=16'h9f8;
17'h3145:	data_out=16'h9f5;
17'h3146:	data_out=16'h8a00;
17'h3147:	data_out=16'h89ec;
17'h3148:	data_out=16'h9ff;
17'h3149:	data_out=16'h8113;
17'h314a:	data_out=16'ha00;
17'h314b:	data_out=16'h866;
17'h314c:	data_out=16'h89f6;
17'h314d:	data_out=16'h177;
17'h314e:	data_out=16'h8381;
17'h314f:	data_out=16'h89e2;
17'h3150:	data_out=16'ha00;
17'h3151:	data_out=16'h885e;
17'h3152:	data_out=16'h89a8;
17'h3153:	data_out=16'ha00;
17'h3154:	data_out=16'ha00;
17'h3155:	data_out=16'h8a00;
17'h3156:	data_out=16'h8a00;
17'h3157:	data_out=16'h8a00;
17'h3158:	data_out=16'h8a00;
17'h3159:	data_out=16'ha00;
17'h315a:	data_out=16'h13;
17'h315b:	data_out=16'ha00;
17'h315c:	data_out=16'h9bd;
17'h315d:	data_out=16'h9ff;
17'h315e:	data_out=16'ha00;
17'h315f:	data_out=16'h899a;
17'h3160:	data_out=16'h8a00;
17'h3161:	data_out=16'ha00;
17'h3162:	data_out=16'h8691;
17'h3163:	data_out=16'h8352;
17'h3164:	data_out=16'h89fb;
17'h3165:	data_out=16'ha00;
17'h3166:	data_out=16'ha00;
17'h3167:	data_out=16'h809f;
17'h3168:	data_out=16'h88b0;
17'h3169:	data_out=16'h8a00;
17'h316a:	data_out=16'h8a00;
17'h316b:	data_out=16'ha00;
17'h316c:	data_out=16'h8a00;
17'h316d:	data_out=16'h842a;
17'h316e:	data_out=16'h8a00;
17'h316f:	data_out=16'ha00;
17'h3170:	data_out=16'h8a00;
17'h3171:	data_out=16'h8a00;
17'h3172:	data_out=16'ha00;
17'h3173:	data_out=16'ha00;
17'h3174:	data_out=16'ha00;
17'h3175:	data_out=16'h9ed;
17'h3176:	data_out=16'h383;
17'h3177:	data_out=16'h96e;
17'h3178:	data_out=16'ha00;
17'h3179:	data_out=16'h8a00;
17'h317a:	data_out=16'h83fd;
17'h317b:	data_out=16'h874a;
17'h317c:	data_out=16'h8a00;
17'h317d:	data_out=16'ha00;
17'h317e:	data_out=16'h84a3;
17'h317f:	data_out=16'ha00;
17'h3180:	data_out=16'h8a00;
17'h3181:	data_out=16'h8a5;
17'h3182:	data_out=16'h8a00;
17'h3183:	data_out=16'h9bc;
17'h3184:	data_out=16'ha00;
17'h3185:	data_out=16'ha00;
17'h3186:	data_out=16'h9ff;
17'h3187:	data_out=16'h9ff;
17'h3188:	data_out=16'h89fc;
17'h3189:	data_out=16'h8747;
17'h318a:	data_out=16'ha00;
17'h318b:	data_out=16'h8701;
17'h318c:	data_out=16'h9f3;
17'h318d:	data_out=16'h74d;
17'h318e:	data_out=16'h8a00;
17'h318f:	data_out=16'h8a00;
17'h3190:	data_out=16'h948;
17'h3191:	data_out=16'h361;
17'h3192:	data_out=16'h8a00;
17'h3193:	data_out=16'h9f4;
17'h3194:	data_out=16'h8341;
17'h3195:	data_out=16'h9fd;
17'h3196:	data_out=16'h9fe;
17'h3197:	data_out=16'h9d2;
17'h3198:	data_out=16'h8a00;
17'h3199:	data_out=16'ha00;
17'h319a:	data_out=16'ha00;
17'h319b:	data_out=16'h68e;
17'h319c:	data_out=16'h9c7;
17'h319d:	data_out=16'h902;
17'h319e:	data_out=16'h897c;
17'h319f:	data_out=16'h16a;
17'h31a0:	data_out=16'ha00;
17'h31a1:	data_out=16'h89b0;
17'h31a2:	data_out=16'h8894;
17'h31a3:	data_out=16'h89ed;
17'h31a4:	data_out=16'h89ed;
17'h31a5:	data_out=16'h89f6;
17'h31a6:	data_out=16'h8a00;
17'h31a7:	data_out=16'h9fe;
17'h31a8:	data_out=16'h87b2;
17'h31a9:	data_out=16'h8a00;
17'h31aa:	data_out=16'h89fd;
17'h31ab:	data_out=16'ha00;
17'h31ac:	data_out=16'ha00;
17'h31ad:	data_out=16'h8a00;
17'h31ae:	data_out=16'h89f1;
17'h31af:	data_out=16'ha00;
17'h31b0:	data_out=16'ha00;
17'h31b1:	data_out=16'ha00;
17'h31b2:	data_out=16'ha00;
17'h31b3:	data_out=16'h871e;
17'h31b4:	data_out=16'h87d1;
17'h31b5:	data_out=16'ha00;
17'h31b6:	data_out=16'h89ef;
17'h31b7:	data_out=16'h8a00;
17'h31b8:	data_out=16'h87b7;
17'h31b9:	data_out=16'h88f9;
17'h31ba:	data_out=16'h894e;
17'h31bb:	data_out=16'ha00;
17'h31bc:	data_out=16'h9c1;
17'h31bd:	data_out=16'h9e6;
17'h31be:	data_out=16'h87a6;
17'h31bf:	data_out=16'ha00;
17'h31c0:	data_out=16'ha00;
17'h31c1:	data_out=16'h87b;
17'h31c2:	data_out=16'h8a00;
17'h31c3:	data_out=16'ha00;
17'h31c4:	data_out=16'ha00;
17'h31c5:	data_out=16'h9fd;
17'h31c6:	data_out=16'h8a00;
17'h31c7:	data_out=16'h8a00;
17'h31c8:	data_out=16'h9ff;
17'h31c9:	data_out=16'h89f3;
17'h31ca:	data_out=16'ha00;
17'h31cb:	data_out=16'h158;
17'h31cc:	data_out=16'h89fe;
17'h31cd:	data_out=16'h83e6;
17'h31ce:	data_out=16'h80db;
17'h31cf:	data_out=16'h89f2;
17'h31d0:	data_out=16'ha00;
17'h31d1:	data_out=16'h8081;
17'h31d2:	data_out=16'h89ea;
17'h31d3:	data_out=16'ha00;
17'h31d4:	data_out=16'ha00;
17'h31d5:	data_out=16'h8a00;
17'h31d6:	data_out=16'h8a00;
17'h31d7:	data_out=16'h8a00;
17'h31d8:	data_out=16'h8a00;
17'h31d9:	data_out=16'ha00;
17'h31da:	data_out=16'h5ee;
17'h31db:	data_out=16'h9f9;
17'h31dc:	data_out=16'h9ff;
17'h31dd:	data_out=16'ha00;
17'h31de:	data_out=16'ha00;
17'h31df:	data_out=16'h89f4;
17'h31e0:	data_out=16'h8a00;
17'h31e1:	data_out=16'ha00;
17'h31e2:	data_out=16'h832f;
17'h31e3:	data_out=16'h80da;
17'h31e4:	data_out=16'h89e8;
17'h31e5:	data_out=16'ha00;
17'h31e6:	data_out=16'ha00;
17'h31e7:	data_out=16'h85c5;
17'h31e8:	data_out=16'h88d8;
17'h31e9:	data_out=16'h8a00;
17'h31ea:	data_out=16'h8a00;
17'h31eb:	data_out=16'ha00;
17'h31ec:	data_out=16'h8a00;
17'h31ed:	data_out=16'h8277;
17'h31ee:	data_out=16'h8a00;
17'h31ef:	data_out=16'ha00;
17'h31f0:	data_out=16'h8a00;
17'h31f1:	data_out=16'h8a00;
17'h31f2:	data_out=16'ha00;
17'h31f3:	data_out=16'ha00;
17'h31f4:	data_out=16'ha00;
17'h31f5:	data_out=16'ha00;
17'h31f6:	data_out=16'h88f2;
17'h31f7:	data_out=16'h83fc;
17'h31f8:	data_out=16'ha00;
17'h31f9:	data_out=16'h8a00;
17'h31fa:	data_out=16'hd6;
17'h31fb:	data_out=16'h87a0;
17'h31fc:	data_out=16'h8a00;
17'h31fd:	data_out=16'ha00;
17'h31fe:	data_out=16'h87c8;
17'h31ff:	data_out=16'ha00;
17'h3200:	data_out=16'h8a00;
17'h3201:	data_out=16'h9fe;
17'h3202:	data_out=16'h8a00;
17'h3203:	data_out=16'h9d1;
17'h3204:	data_out=16'ha00;
17'h3205:	data_out=16'ha00;
17'h3206:	data_out=16'ha00;
17'h3207:	data_out=16'h9fb;
17'h3208:	data_out=16'h8a00;
17'h3209:	data_out=16'h8258;
17'h320a:	data_out=16'h9fe;
17'h320b:	data_out=16'h78f;
17'h320c:	data_out=16'h9f5;
17'h320d:	data_out=16'h387;
17'h320e:	data_out=16'h8a00;
17'h320f:	data_out=16'h8a00;
17'h3210:	data_out=16'h9ef;
17'h3211:	data_out=16'h6ed;
17'h3212:	data_out=16'h8a00;
17'h3213:	data_out=16'h9fd;
17'h3214:	data_out=16'h3f;
17'h3215:	data_out=16'h4a6;
17'h3216:	data_out=16'h9fd;
17'h3217:	data_out=16'h9f9;
17'h3218:	data_out=16'h8a00;
17'h3219:	data_out=16'ha00;
17'h321a:	data_out=16'ha00;
17'h321b:	data_out=16'h9c3;
17'h321c:	data_out=16'h9da;
17'h321d:	data_out=16'h9ea;
17'h321e:	data_out=16'h8589;
17'h321f:	data_out=16'h3ad;
17'h3220:	data_out=16'h9fd;
17'h3221:	data_out=16'h8a00;
17'h3222:	data_out=16'h835d;
17'h3223:	data_out=16'h89f6;
17'h3224:	data_out=16'h89f6;
17'h3225:	data_out=16'h846b;
17'h3226:	data_out=16'h8a00;
17'h3227:	data_out=16'h9fc;
17'h3228:	data_out=16'h87da;
17'h3229:	data_out=16'h8a00;
17'h322a:	data_out=16'h8a00;
17'h322b:	data_out=16'h9f7;
17'h322c:	data_out=16'h9ff;
17'h322d:	data_out=16'h8a00;
17'h322e:	data_out=16'h88ed;
17'h322f:	data_out=16'ha00;
17'h3230:	data_out=16'ha00;
17'h3231:	data_out=16'ha00;
17'h3232:	data_out=16'ha00;
17'h3233:	data_out=16'h83db;
17'h3234:	data_out=16'h880b;
17'h3235:	data_out=16'ha00;
17'h3236:	data_out=16'h89e0;
17'h3237:	data_out=16'h8a00;
17'h3238:	data_out=16'h341;
17'h3239:	data_out=16'h88c2;
17'h323a:	data_out=16'h891a;
17'h323b:	data_out=16'ha00;
17'h323c:	data_out=16'h9ed;
17'h323d:	data_out=16'h980;
17'h323e:	data_out=16'h87ca;
17'h323f:	data_out=16'ha00;
17'h3240:	data_out=16'ha00;
17'h3241:	data_out=16'h9d9;
17'h3242:	data_out=16'h89fc;
17'h3243:	data_out=16'ha00;
17'h3244:	data_out=16'h9fe;
17'h3245:	data_out=16'h5d5;
17'h3246:	data_out=16'h8a00;
17'h3247:	data_out=16'h8a00;
17'h3248:	data_out=16'ha00;
17'h3249:	data_out=16'h81a0;
17'h324a:	data_out=16'ha00;
17'h324b:	data_out=16'h254;
17'h324c:	data_out=16'h8a00;
17'h324d:	data_out=16'h22e;
17'h324e:	data_out=16'h2f1;
17'h324f:	data_out=16'h89f8;
17'h3250:	data_out=16'ha00;
17'h3251:	data_out=16'h8072;
17'h3252:	data_out=16'h89f7;
17'h3253:	data_out=16'ha00;
17'h3254:	data_out=16'h9f6;
17'h3255:	data_out=16'h88da;
17'h3256:	data_out=16'h8a00;
17'h3257:	data_out=16'h8a00;
17'h3258:	data_out=16'h8a00;
17'h3259:	data_out=16'ha00;
17'h325a:	data_out=16'h9d5;
17'h325b:	data_out=16'h9f1;
17'h325c:	data_out=16'ha00;
17'h325d:	data_out=16'ha00;
17'h325e:	data_out=16'ha00;
17'h325f:	data_out=16'h89fc;
17'h3260:	data_out=16'h8a00;
17'h3261:	data_out=16'ha00;
17'h3262:	data_out=16'h15f;
17'h3263:	data_out=16'h46d;
17'h3264:	data_out=16'h89fe;
17'h3265:	data_out=16'ha00;
17'h3266:	data_out=16'ha00;
17'h3267:	data_out=16'h82d2;
17'h3268:	data_out=16'h893e;
17'h3269:	data_out=16'h8a00;
17'h326a:	data_out=16'h8a00;
17'h326b:	data_out=16'ha00;
17'h326c:	data_out=16'h8a00;
17'h326d:	data_out=16'h2d6;
17'h326e:	data_out=16'h8a00;
17'h326f:	data_out=16'ha00;
17'h3270:	data_out=16'h8a00;
17'h3271:	data_out=16'h8a00;
17'h3272:	data_out=16'ha00;
17'h3273:	data_out=16'ha00;
17'h3274:	data_out=16'ha00;
17'h3275:	data_out=16'ha00;
17'h3276:	data_out=16'h8348;
17'h3277:	data_out=16'h466;
17'h3278:	data_out=16'ha00;
17'h3279:	data_out=16'h8a00;
17'h327a:	data_out=16'h51a;
17'h327b:	data_out=16'h87c4;
17'h327c:	data_out=16'h8a00;
17'h327d:	data_out=16'ha00;
17'h327e:	data_out=16'h38b;
17'h327f:	data_out=16'ha00;
17'h3280:	data_out=16'h8a00;
17'h3281:	data_out=16'h9fe;
17'h3282:	data_out=16'h8815;
17'h3283:	data_out=16'h9d1;
17'h3284:	data_out=16'ha00;
17'h3285:	data_out=16'ha00;
17'h3286:	data_out=16'ha00;
17'h3287:	data_out=16'ha00;
17'h3288:	data_out=16'h88e9;
17'h3289:	data_out=16'h2a4;
17'h328a:	data_out=16'ha00;
17'h328b:	data_out=16'h917;
17'h328c:	data_out=16'ha00;
17'h328d:	data_out=16'h82f7;
17'h328e:	data_out=16'h85f6;
17'h328f:	data_out=16'h89fb;
17'h3290:	data_out=16'h997;
17'h3291:	data_out=16'h9e2;
17'h3292:	data_out=16'h8a00;
17'h3293:	data_out=16'ha00;
17'h3294:	data_out=16'h8440;
17'h3295:	data_out=16'h8765;
17'h3296:	data_out=16'h5ef;
17'h3297:	data_out=16'h9ff;
17'h3298:	data_out=16'h8a00;
17'h3299:	data_out=16'ha00;
17'h329a:	data_out=16'ha00;
17'h329b:	data_out=16'h9e8;
17'h329c:	data_out=16'h9e1;
17'h329d:	data_out=16'h9fc;
17'h329e:	data_out=16'h868d;
17'h329f:	data_out=16'h8069;
17'h32a0:	data_out=16'h9eb;
17'h32a1:	data_out=16'h84c7;
17'h32a2:	data_out=16'h909;
17'h32a3:	data_out=16'h741;
17'h32a4:	data_out=16'h733;
17'h32a5:	data_out=16'h801;
17'h32a6:	data_out=16'h8a00;
17'h32a7:	data_out=16'h9fd;
17'h32a8:	data_out=16'h8273;
17'h32a9:	data_out=16'h8a00;
17'h32aa:	data_out=16'h8899;
17'h32ab:	data_out=16'h9f6;
17'h32ac:	data_out=16'h64e;
17'h32ad:	data_out=16'h8a00;
17'h32ae:	data_out=16'h87eb;
17'h32af:	data_out=16'ha00;
17'h32b0:	data_out=16'ha00;
17'h32b1:	data_out=16'ha00;
17'h32b2:	data_out=16'ha00;
17'h32b3:	data_out=16'h86c9;
17'h32b4:	data_out=16'h895c;
17'h32b5:	data_out=16'h9fb;
17'h32b6:	data_out=16'h88af;
17'h32b7:	data_out=16'h8173;
17'h32b8:	data_out=16'h7fb;
17'h32b9:	data_out=16'h89fd;
17'h32ba:	data_out=16'h85ae;
17'h32bb:	data_out=16'ha00;
17'h32bc:	data_out=16'h9fc;
17'h32bd:	data_out=16'h370;
17'h32be:	data_out=16'h825e;
17'h32bf:	data_out=16'ha00;
17'h32c0:	data_out=16'ha00;
17'h32c1:	data_out=16'h9e7;
17'h32c2:	data_out=16'h89f6;
17'h32c3:	data_out=16'ha00;
17'h32c4:	data_out=16'h9f5;
17'h32c5:	data_out=16'h869d;
17'h32c6:	data_out=16'h8a00;
17'h32c7:	data_out=16'h8a00;
17'h32c8:	data_out=16'ha00;
17'h32c9:	data_out=16'h7b7;
17'h32ca:	data_out=16'ha00;
17'h32cb:	data_out=16'h29f;
17'h32cc:	data_out=16'h58f;
17'h32cd:	data_out=16'h9b7;
17'h32ce:	data_out=16'h95a;
17'h32cf:	data_out=16'h8274;
17'h32d0:	data_out=16'ha00;
17'h32d1:	data_out=16'h8215;
17'h32d2:	data_out=16'h515;
17'h32d3:	data_out=16'ha00;
17'h32d4:	data_out=16'h9ec;
17'h32d5:	data_out=16'h8850;
17'h32d6:	data_out=16'h8a00;
17'h32d7:	data_out=16'h8a00;
17'h32d8:	data_out=16'h8893;
17'h32d9:	data_out=16'ha00;
17'h32da:	data_out=16'h9f5;
17'h32db:	data_out=16'h9ed;
17'h32dc:	data_out=16'ha00;
17'h32dd:	data_out=16'h9ff;
17'h32de:	data_out=16'ha00;
17'h32df:	data_out=16'h8a00;
17'h32e0:	data_out=16'h89ea;
17'h32e1:	data_out=16'ha00;
17'h32e2:	data_out=16'h265;
17'h32e3:	data_out=16'h128;
17'h32e4:	data_out=16'h89fe;
17'h32e5:	data_out=16'ha00;
17'h32e6:	data_out=16'ha00;
17'h32e7:	data_out=16'h89f8;
17'h32e8:	data_out=16'h83f6;
17'h32e9:	data_out=16'h8a00;
17'h32ea:	data_out=16'h86d8;
17'h32eb:	data_out=16'ha00;
17'h32ec:	data_out=16'h8a00;
17'h32ed:	data_out=16'h804d;
17'h32ee:	data_out=16'h86d3;
17'h32ef:	data_out=16'ha00;
17'h32f0:	data_out=16'h8654;
17'h32f1:	data_out=16'h8919;
17'h32f2:	data_out=16'ha00;
17'h32f3:	data_out=16'ha00;
17'h32f4:	data_out=16'ha00;
17'h32f5:	data_out=16'ha00;
17'h32f6:	data_out=16'h80bd;
17'h32f7:	data_out=16'h938;
17'h32f8:	data_out=16'ha00;
17'h32f9:	data_out=16'h8694;
17'h32fa:	data_out=16'h1f6;
17'h32fb:	data_out=16'h8255;
17'h32fc:	data_out=16'h8a00;
17'h32fd:	data_out=16'h9f7;
17'h32fe:	data_out=16'h804;
17'h32ff:	data_out=16'h9fe;
17'h3300:	data_out=16'h89fe;
17'h3301:	data_out=16'h276;
17'h3302:	data_out=16'h5b8;
17'h3303:	data_out=16'h9d1;
17'h3304:	data_out=16'ha00;
17'h3305:	data_out=16'ha00;
17'h3306:	data_out=16'ha00;
17'h3307:	data_out=16'ha00;
17'h3308:	data_out=16'h8813;
17'h3309:	data_out=16'h181;
17'h330a:	data_out=16'h530;
17'h330b:	data_out=16'h5c7;
17'h330c:	data_out=16'h9fe;
17'h330d:	data_out=16'h9de;
17'h330e:	data_out=16'h167;
17'h330f:	data_out=16'h856a;
17'h3310:	data_out=16'h79b;
17'h3311:	data_out=16'h9fd;
17'h3312:	data_out=16'h8a00;
17'h3313:	data_out=16'ha00;
17'h3314:	data_out=16'h860e;
17'h3315:	data_out=16'h8797;
17'h3316:	data_out=16'ha00;
17'h3317:	data_out=16'h9fb;
17'h3318:	data_out=16'h8a00;
17'h3319:	data_out=16'ha00;
17'h331a:	data_out=16'ha00;
17'h331b:	data_out=16'h9f6;
17'h331c:	data_out=16'h9ee;
17'h331d:	data_out=16'h9fe;
17'h331e:	data_out=16'h86ab;
17'h331f:	data_out=16'h157;
17'h3320:	data_out=16'h9dd;
17'h3321:	data_out=16'h25d;
17'h3322:	data_out=16'h941;
17'h3323:	data_out=16'h9ff;
17'h3324:	data_out=16'h9ff;
17'h3325:	data_out=16'h87f;
17'h3326:	data_out=16'h89f6;
17'h3327:	data_out=16'h9fc;
17'h3328:	data_out=16'h452;
17'h3329:	data_out=16'h8a00;
17'h332a:	data_out=16'h844d;
17'h332b:	data_out=16'h503;
17'h332c:	data_out=16'h9fd;
17'h332d:	data_out=16'h8a00;
17'h332e:	data_out=16'h8755;
17'h332f:	data_out=16'ha00;
17'h3330:	data_out=16'ha00;
17'h3331:	data_out=16'h1aa;
17'h3332:	data_out=16'ha00;
17'h3333:	data_out=16'h89fc;
17'h3334:	data_out=16'h89d8;
17'h3335:	data_out=16'h9fc;
17'h3336:	data_out=16'h8867;
17'h3337:	data_out=16'h9e8;
17'h3338:	data_out=16'h88a;
17'h3339:	data_out=16'h89fd;
17'h333a:	data_out=16'h880d;
17'h333b:	data_out=16'ha00;
17'h333c:	data_out=16'ha00;
17'h333d:	data_out=16'h89fb;
17'h333e:	data_out=16'h465;
17'h333f:	data_out=16'ha00;
17'h3340:	data_out=16'ha00;
17'h3341:	data_out=16'h9f4;
17'h3342:	data_out=16'h80b8;
17'h3343:	data_out=16'h9fe;
17'h3344:	data_out=16'h9f3;
17'h3345:	data_out=16'h86a5;
17'h3346:	data_out=16'h82ea;
17'h3347:	data_out=16'h8a00;
17'h3348:	data_out=16'ha00;
17'h3349:	data_out=16'h844;
17'h334a:	data_out=16'ha00;
17'h334b:	data_out=16'h3d3;
17'h334c:	data_out=16'h83d;
17'h334d:	data_out=16'h9c5;
17'h334e:	data_out=16'h9e6;
17'h334f:	data_out=16'h63c;
17'h3350:	data_out=16'ha00;
17'h3351:	data_out=16'h2cf;
17'h3352:	data_out=16'h7aa;
17'h3353:	data_out=16'ha00;
17'h3354:	data_out=16'h9e2;
17'h3355:	data_out=16'h822e;
17'h3356:	data_out=16'h89c3;
17'h3357:	data_out=16'h8a00;
17'h3358:	data_out=16'h8772;
17'h3359:	data_out=16'ha00;
17'h335a:	data_out=16'h9f3;
17'h335b:	data_out=16'h9f0;
17'h335c:	data_out=16'ha00;
17'h335d:	data_out=16'h9f7;
17'h335e:	data_out=16'ha00;
17'h335f:	data_out=16'h8a00;
17'h3360:	data_out=16'h89e1;
17'h3361:	data_out=16'ha00;
17'h3362:	data_out=16'h63f;
17'h3363:	data_out=16'h8394;
17'h3364:	data_out=16'h89fe;
17'h3365:	data_out=16'ha00;
17'h3366:	data_out=16'ha00;
17'h3367:	data_out=16'h89ff;
17'h3368:	data_out=16'h301;
17'h3369:	data_out=16'h89ff;
17'h336a:	data_out=16'hb8;
17'h336b:	data_out=16'ha00;
17'h336c:	data_out=16'h89fd;
17'h336d:	data_out=16'h8500;
17'h336e:	data_out=16'hbd;
17'h336f:	data_out=16'ha00;
17'h3370:	data_out=16'h121;
17'h3371:	data_out=16'h892c;
17'h3372:	data_out=16'ha00;
17'h3373:	data_out=16'ha00;
17'h3374:	data_out=16'ha00;
17'h3375:	data_out=16'ha00;
17'h3376:	data_out=16'h89e6;
17'h3377:	data_out=16'h9a1;
17'h3378:	data_out=16'ha00;
17'h3379:	data_out=16'h30e;
17'h337a:	data_out=16'h80ee;
17'h337b:	data_out=16'h46e;
17'h337c:	data_out=16'h8a00;
17'h337d:	data_out=16'h9e1;
17'h337e:	data_out=16'h779;
17'h337f:	data_out=16'h9f3;
17'h3380:	data_out=16'h89ff;
17'h3381:	data_out=16'h84cb;
17'h3382:	data_out=16'h9e0;
17'h3383:	data_out=16'h9eb;
17'h3384:	data_out=16'h9fb;
17'h3385:	data_out=16'ha00;
17'h3386:	data_out=16'h9fe;
17'h3387:	data_out=16'ha00;
17'h3388:	data_out=16'h8875;
17'h3389:	data_out=16'h539;
17'h338a:	data_out=16'h8374;
17'h338b:	data_out=16'h566;
17'h338c:	data_out=16'h9f7;
17'h338d:	data_out=16'h9ea;
17'h338e:	data_out=16'h2e0;
17'h338f:	data_out=16'h45d;
17'h3390:	data_out=16'h85b;
17'h3391:	data_out=16'h9f6;
17'h3392:	data_out=16'h89fe;
17'h3393:	data_out=16'h9fd;
17'h3394:	data_out=16'h814a;
17'h3395:	data_out=16'h825a;
17'h3396:	data_out=16'h9ff;
17'h3397:	data_out=16'h9f6;
17'h3398:	data_out=16'h89fb;
17'h3399:	data_out=16'ha00;
17'h339a:	data_out=16'ha00;
17'h339b:	data_out=16'h9ed;
17'h339c:	data_out=16'h9ef;
17'h339d:	data_out=16'h8fd;
17'h339e:	data_out=16'ha0;
17'h339f:	data_out=16'h9ec;
17'h33a0:	data_out=16'h9ea;
17'h33a1:	data_out=16'h388;
17'h33a2:	data_out=16'h9af;
17'h33a3:	data_out=16'h6ba;
17'h33a4:	data_out=16'h6b8;
17'h33a5:	data_out=16'h95e;
17'h33a6:	data_out=16'h89ff;
17'h33a7:	data_out=16'ha00;
17'h33a8:	data_out=16'h4f3;
17'h33a9:	data_out=16'h8a00;
17'h33aa:	data_out=16'h8207;
17'h33ab:	data_out=16'h83de;
17'h33ac:	data_out=16'h9ff;
17'h33ad:	data_out=16'h8a00;
17'h33ae:	data_out=16'h8271;
17'h33af:	data_out=16'ha00;
17'h33b0:	data_out=16'ha00;
17'h33b1:	data_out=16'h80bc;
17'h33b2:	data_out=16'ha00;
17'h33b3:	data_out=16'h84e7;
17'h33b4:	data_out=16'h89ea;
17'h33b5:	data_out=16'h9f9;
17'h33b6:	data_out=16'h8860;
17'h33b7:	data_out=16'h9e3;
17'h33b8:	data_out=16'h948;
17'h33b9:	data_out=16'h88f3;
17'h33ba:	data_out=16'h8219;
17'h33bb:	data_out=16'ha00;
17'h33bc:	data_out=16'h9fb;
17'h33bd:	data_out=16'h87b9;
17'h33be:	data_out=16'h502;
17'h33bf:	data_out=16'ha00;
17'h33c0:	data_out=16'ha00;
17'h33c1:	data_out=16'h9ea;
17'h33c2:	data_out=16'h8410;
17'h33c3:	data_out=16'ha00;
17'h33c4:	data_out=16'h9fa;
17'h33c5:	data_out=16'h817f;
17'h33c6:	data_out=16'h8a00;
17'h33c7:	data_out=16'h8a00;
17'h33c8:	data_out=16'h9fe;
17'h33c9:	data_out=16'h94f;
17'h33ca:	data_out=16'ha00;
17'h33cb:	data_out=16'h54b;
17'h33cc:	data_out=16'h92b;
17'h33cd:	data_out=16'h9e8;
17'h33ce:	data_out=16'h979;
17'h33cf:	data_out=16'h860;
17'h33d0:	data_out=16'ha00;
17'h33d1:	data_out=16'h7db;
17'h33d2:	data_out=16'h400;
17'h33d3:	data_out=16'h9fd;
17'h33d4:	data_out=16'h9ee;
17'h33d5:	data_out=16'h49a;
17'h33d6:	data_out=16'h89aa;
17'h33d7:	data_out=16'h89ff;
17'h33d8:	data_out=16'h8448;
17'h33d9:	data_out=16'ha00;
17'h33da:	data_out=16'h9f1;
17'h33db:	data_out=16'h9ee;
17'h33dc:	data_out=16'h9ff;
17'h33dd:	data_out=16'h9f2;
17'h33de:	data_out=16'ha00;
17'h33df:	data_out=16'h89ff;
17'h33e0:	data_out=16'h89fb;
17'h33e1:	data_out=16'ha00;
17'h33e2:	data_out=16'h9f2;
17'h33e3:	data_out=16'h67;
17'h33e4:	data_out=16'h89ff;
17'h33e5:	data_out=16'ha00;
17'h33e6:	data_out=16'ha00;
17'h33e7:	data_out=16'h89fe;
17'h33e8:	data_out=16'h3f1;
17'h33e9:	data_out=16'h89f9;
17'h33ea:	data_out=16'h265;
17'h33eb:	data_out=16'ha00;
17'h33ec:	data_out=16'h89fe;
17'h33ed:	data_out=16'h8097;
17'h33ee:	data_out=16'h268;
17'h33ef:	data_out=16'ha00;
17'h33f0:	data_out=16'h2af;
17'h33f1:	data_out=16'h81bb;
17'h33f2:	data_out=16'h9ff;
17'h33f3:	data_out=16'ha00;
17'h33f4:	data_out=16'ha00;
17'h33f5:	data_out=16'ha00;
17'h33f6:	data_out=16'h89d8;
17'h33f7:	data_out=16'h9dd;
17'h33f8:	data_out=16'ha00;
17'h33f9:	data_out=16'h60c;
17'h33fa:	data_out=16'h2ab;
17'h33fb:	data_out=16'h509;
17'h33fc:	data_out=16'h89ef;
17'h33fd:	data_out=16'h9f8;
17'h33fe:	data_out=16'h825;
17'h33ff:	data_out=16'h9f9;
17'h3400:	data_out=16'h89fe;
17'h3401:	data_out=16'h8814;
17'h3402:	data_out=16'h9e8;
17'h3403:	data_out=16'h9de;
17'h3404:	data_out=16'h9fe;
17'h3405:	data_out=16'ha00;
17'h3406:	data_out=16'h9fe;
17'h3407:	data_out=16'ha00;
17'h3408:	data_out=16'h86de;
17'h3409:	data_out=16'h809a;
17'h340a:	data_out=16'h8872;
17'h340b:	data_out=16'h814c;
17'h340c:	data_out=16'h9fa;
17'h340d:	data_out=16'h9f4;
17'h340e:	data_out=16'h374;
17'h340f:	data_out=16'h9ea;
17'h3410:	data_out=16'h90;
17'h3411:	data_out=16'h9c0;
17'h3412:	data_out=16'h89c9;
17'h3413:	data_out=16'h9fc;
17'h3414:	data_out=16'h9;
17'h3415:	data_out=16'h176;
17'h3416:	data_out=16'ha00;
17'h3417:	data_out=16'h7da;
17'h3418:	data_out=16'h84ec;
17'h3419:	data_out=16'ha00;
17'h341a:	data_out=16'ha00;
17'h341b:	data_out=16'h9f1;
17'h341c:	data_out=16'h9de;
17'h341d:	data_out=16'h8826;
17'h341e:	data_out=16'h2d5;
17'h341f:	data_out=16'h979;
17'h3420:	data_out=16'h890;
17'h3421:	data_out=16'h3e2;
17'h3422:	data_out=16'h726;
17'h3423:	data_out=16'h6b1;
17'h3424:	data_out=16'h6bf;
17'h3425:	data_out=16'h9ee;
17'h3426:	data_out=16'h89ff;
17'h3427:	data_out=16'h8059;
17'h3428:	data_out=16'h4c7;
17'h3429:	data_out=16'h8a00;
17'h342a:	data_out=16'h14f;
17'h342b:	data_out=16'h89ea;
17'h342c:	data_out=16'h9ff;
17'h342d:	data_out=16'h8a00;
17'h342e:	data_out=16'h276;
17'h342f:	data_out=16'ha00;
17'h3430:	data_out=16'ha00;
17'h3431:	data_out=16'h8691;
17'h3432:	data_out=16'ha00;
17'h3433:	data_out=16'h8292;
17'h3434:	data_out=16'h89fe;
17'h3435:	data_out=16'h9ee;
17'h3436:	data_out=16'h8222;
17'h3437:	data_out=16'h9ec;
17'h3438:	data_out=16'h238;
17'h3439:	data_out=16'h843b;
17'h343a:	data_out=16'h857c;
17'h343b:	data_out=16'ha00;
17'h343c:	data_out=16'h9bb;
17'h343d:	data_out=16'h824a;
17'h343e:	data_out=16'h4d0;
17'h343f:	data_out=16'ha00;
17'h3440:	data_out=16'ha00;
17'h3441:	data_out=16'h9e0;
17'h3442:	data_out=16'h8400;
17'h3443:	data_out=16'h9fe;
17'h3444:	data_out=16'h9f8;
17'h3445:	data_out=16'h205;
17'h3446:	data_out=16'h8a00;
17'h3447:	data_out=16'h869c;
17'h3448:	data_out=16'ha00;
17'h3449:	data_out=16'h9ed;
17'h344a:	data_out=16'ha00;
17'h344b:	data_out=16'h6bb;
17'h344c:	data_out=16'h9ec;
17'h344d:	data_out=16'h7d2;
17'h344e:	data_out=16'h979;
17'h344f:	data_out=16'h92d;
17'h3450:	data_out=16'h9fc;
17'h3451:	data_out=16'h9d9;
17'h3452:	data_out=16'h3b5;
17'h3453:	data_out=16'h9ff;
17'h3454:	data_out=16'h992;
17'h3455:	data_out=16'h9e8;
17'h3456:	data_out=16'h85c8;
17'h3457:	data_out=16'h89ed;
17'h3458:	data_out=16'h808;
17'h3459:	data_out=16'ha00;
17'h345a:	data_out=16'h9c6;
17'h345b:	data_out=16'h811;
17'h345c:	data_out=16'h9f8;
17'h345d:	data_out=16'h9fa;
17'h345e:	data_out=16'ha00;
17'h345f:	data_out=16'h8391;
17'h3460:	data_out=16'h89ff;
17'h3461:	data_out=16'ha00;
17'h3462:	data_out=16'h99a;
17'h3463:	data_out=16'h56;
17'h3464:	data_out=16'h8a00;
17'h3465:	data_out=16'ha00;
17'h3466:	data_out=16'ha00;
17'h3467:	data_out=16'h8a00;
17'h3468:	data_out=16'h429;
17'h3469:	data_out=16'h89e5;
17'h346a:	data_out=16'h329;
17'h346b:	data_out=16'ha00;
17'h346c:	data_out=16'h89fe;
17'h346d:	data_out=16'h803b;
17'h346e:	data_out=16'h32b;
17'h346f:	data_out=16'ha00;
17'h3470:	data_out=16'h356;
17'h3471:	data_out=16'h748;
17'h3472:	data_out=16'ha00;
17'h3473:	data_out=16'ha00;
17'h3474:	data_out=16'ha00;
17'h3475:	data_out=16'ha00;
17'h3476:	data_out=16'h89f8;
17'h3477:	data_out=16'h9f6;
17'h3478:	data_out=16'ha00;
17'h3479:	data_out=16'h9d7;
17'h347a:	data_out=16'h265;
17'h347b:	data_out=16'h4d5;
17'h347c:	data_out=16'h827b;
17'h347d:	data_out=16'h9fa;
17'h347e:	data_out=16'h80f8;
17'h347f:	data_out=16'h9fe;
17'h3480:	data_out=16'h83fc;
17'h3481:	data_out=16'h87be;
17'h3482:	data_out=16'h91e;
17'h3483:	data_out=16'h897;
17'h3484:	data_out=16'h9fb;
17'h3485:	data_out=16'h9ff;
17'h3486:	data_out=16'h8e1;
17'h3487:	data_out=16'h9ff;
17'h3488:	data_out=16'h8404;
17'h3489:	data_out=16'h8792;
17'h348a:	data_out=16'h88c4;
17'h348b:	data_out=16'h8a00;
17'h348c:	data_out=16'h9f7;
17'h348d:	data_out=16'h9f8;
17'h348e:	data_out=16'h262;
17'h348f:	data_out=16'h897;
17'h3490:	data_out=16'h8745;
17'h3491:	data_out=16'h835;
17'h3492:	data_out=16'h89d3;
17'h3493:	data_out=16'h9fc;
17'h3494:	data_out=16'h8632;
17'h3495:	data_out=16'h39a;
17'h3496:	data_out=16'h9fb;
17'h3497:	data_out=16'h84d6;
17'h3498:	data_out=16'h377;
17'h3499:	data_out=16'h9fc;
17'h349a:	data_out=16'h9fd;
17'h349b:	data_out=16'h1e8;
17'h349c:	data_out=16'h22b;
17'h349d:	data_out=16'h8a00;
17'h349e:	data_out=16'h81ee;
17'h349f:	data_out=16'h777;
17'h34a0:	data_out=16'h8205;
17'h34a1:	data_out=16'h298;
17'h34a2:	data_out=16'h838c;
17'h34a3:	data_out=16'h66e;
17'h34a4:	data_out=16'h678;
17'h34a5:	data_out=16'h9fe;
17'h34a6:	data_out=16'h89fa;
17'h34a7:	data_out=16'h89f8;
17'h34a8:	data_out=16'h3d8;
17'h34a9:	data_out=16'h8a00;
17'h34aa:	data_out=16'h80c5;
17'h34ab:	data_out=16'h8a00;
17'h34ac:	data_out=16'h9fb;
17'h34ad:	data_out=16'h8a00;
17'h34ae:	data_out=16'h845e;
17'h34af:	data_out=16'h1c1;
17'h34b0:	data_out=16'ha00;
17'h34b1:	data_out=16'h89fe;
17'h34b2:	data_out=16'h9ff;
17'h34b3:	data_out=16'h8819;
17'h34b4:	data_out=16'h8a00;
17'h34b5:	data_out=16'h9c8;
17'h34b6:	data_out=16'h8269;
17'h34b7:	data_out=16'h6c4;
17'h34b8:	data_out=16'h839c;
17'h34b9:	data_out=16'h87be;
17'h34ba:	data_out=16'h8900;
17'h34bb:	data_out=16'h8218;
17'h34bc:	data_out=16'h80db;
17'h34bd:	data_out=16'haa;
17'h34be:	data_out=16'h3f6;
17'h34bf:	data_out=16'h9fe;
17'h34c0:	data_out=16'ha00;
17'h34c1:	data_out=16'h9de;
17'h34c2:	data_out=16'h82c2;
17'h34c3:	data_out=16'h9fc;
17'h34c4:	data_out=16'h80b6;
17'h34c5:	data_out=16'h3e9;
17'h34c6:	data_out=16'h89fa;
17'h34c7:	data_out=16'h8546;
17'h34c8:	data_out=16'hf5;
17'h34c9:	data_out=16'h9fe;
17'h34ca:	data_out=16'h9fd;
17'h34cb:	data_out=16'h9c;
17'h34cc:	data_out=16'ha00;
17'h34cd:	data_out=16'h8375;
17'h34ce:	data_out=16'h8193;
17'h34cf:	data_out=16'h9dd;
17'h34d0:	data_out=16'h9f3;
17'h34d1:	data_out=16'h9ee;
17'h34d2:	data_out=16'h6ae;
17'h34d3:	data_out=16'h833b;
17'h34d4:	data_out=16'h8286;
17'h34d5:	data_out=16'h370;
17'h34d6:	data_out=16'h75c;
17'h34d7:	data_out=16'h822b;
17'h34d8:	data_out=16'h959;
17'h34d9:	data_out=16'h9ff;
17'h34da:	data_out=16'h84dd;
17'h34db:	data_out=16'h844e;
17'h34dc:	data_out=16'h8204;
17'h34dd:	data_out=16'h9f7;
17'h34de:	data_out=16'h25b;
17'h34df:	data_out=16'h50;
17'h34e0:	data_out=16'h89ff;
17'h34e1:	data_out=16'h1a8;
17'h34e2:	data_out=16'h7a6;
17'h34e3:	data_out=16'h8796;
17'h34e4:	data_out=16'h8a00;
17'h34e5:	data_out=16'ha00;
17'h34e6:	data_out=16'h9fe;
17'h34e7:	data_out=16'h8a00;
17'h34e8:	data_out=16'h301;
17'h34e9:	data_out=16'h892a;
17'h34ea:	data_out=16'h253;
17'h34eb:	data_out=16'h9ff;
17'h34ec:	data_out=16'hb3;
17'h34ed:	data_out=16'h879c;
17'h34ee:	data_out=16'h254;
17'h34ef:	data_out=16'h9ff;
17'h34f0:	data_out=16'h25d;
17'h34f1:	data_out=16'h9f5;
17'h34f2:	data_out=16'h9fc;
17'h34f3:	data_out=16'h9fc;
17'h34f4:	data_out=16'ha00;
17'h34f5:	data_out=16'h856;
17'h34f6:	data_out=16'h8a00;
17'h34f7:	data_out=16'h9f7;
17'h34f8:	data_out=16'h9f5;
17'h34f9:	data_out=16'h5b2;
17'h34fa:	data_out=16'h85c8;
17'h34fb:	data_out=16'h411;
17'h34fc:	data_out=16'h2ce;
17'h34fd:	data_out=16'h9f4;
17'h34fe:	data_out=16'h8992;
17'h34ff:	data_out=16'h9ff;
17'h3500:	data_out=16'h825d;
17'h3501:	data_out=16'h89e2;
17'h3502:	data_out=16'ha00;
17'h3503:	data_out=16'h29e;
17'h3504:	data_out=16'h9fa;
17'h3505:	data_out=16'ha00;
17'h3506:	data_out=16'h444;
17'h3507:	data_out=16'h91f;
17'h3508:	data_out=16'h804f;
17'h3509:	data_out=16'h869d;
17'h350a:	data_out=16'h89ff;
17'h350b:	data_out=16'h8a00;
17'h350c:	data_out=16'h9f5;
17'h350d:	data_out=16'ha00;
17'h350e:	data_out=16'h2cd;
17'h350f:	data_out=16'h9ff;
17'h3510:	data_out=16'h884d;
17'h3511:	data_out=16'h4fd;
17'h3512:	data_out=16'h8936;
17'h3513:	data_out=16'h6c5;
17'h3514:	data_out=16'h89a1;
17'h3515:	data_out=16'h314;
17'h3516:	data_out=16'h7d2;
17'h3517:	data_out=16'h89f8;
17'h3518:	data_out=16'h653;
17'h3519:	data_out=16'h823;
17'h351a:	data_out=16'h9ff;
17'h351b:	data_out=16'h8379;
17'h351c:	data_out=16'h84a0;
17'h351d:	data_out=16'h8a00;
17'h351e:	data_out=16'h8553;
17'h351f:	data_out=16'h78a;
17'h3520:	data_out=16'h868b;
17'h3521:	data_out=16'h2cd;
17'h3522:	data_out=16'h8264;
17'h3523:	data_out=16'h813;
17'h3524:	data_out=16'h81a;
17'h3525:	data_out=16'h9ff;
17'h3526:	data_out=16'h85b2;
17'h3527:	data_out=16'h89ff;
17'h3528:	data_out=16'h2c3;
17'h3529:	data_out=16'h89ff;
17'h352a:	data_out=16'h8019;
17'h352b:	data_out=16'h8a00;
17'h352c:	data_out=16'h664;
17'h352d:	data_out=16'h8a00;
17'h352e:	data_out=16'h116;
17'h352f:	data_out=16'h84f4;
17'h3530:	data_out=16'ha00;
17'h3531:	data_out=16'h89ff;
17'h3532:	data_out=16'ha00;
17'h3533:	data_out=16'h8a00;
17'h3534:	data_out=16'h8a00;
17'h3535:	data_out=16'h9f3;
17'h3536:	data_out=16'h80de;
17'h3537:	data_out=16'h8f9;
17'h3538:	data_out=16'h8851;
17'h3539:	data_out=16'h89b1;
17'h353a:	data_out=16'h8961;
17'h353b:	data_out=16'h853e;
17'h353c:	data_out=16'h85a7;
17'h353d:	data_out=16'h824e;
17'h353e:	data_out=16'h2c3;
17'h353f:	data_out=16'ha00;
17'h3540:	data_out=16'ha00;
17'h3541:	data_out=16'h899;
17'h3542:	data_out=16'h789;
17'h3543:	data_out=16'h820;
17'h3544:	data_out=16'h86bc;
17'h3545:	data_out=16'h339;
17'h3546:	data_out=16'h89d1;
17'h3547:	data_out=16'h9;
17'h3548:	data_out=16'h8178;
17'h3549:	data_out=16'ha00;
17'h354a:	data_out=16'h9fb;
17'h354b:	data_out=16'h414;
17'h354c:	data_out=16'ha00;
17'h354d:	data_out=16'h82e3;
17'h354e:	data_out=16'h6b;
17'h354f:	data_out=16'h9fc;
17'h3550:	data_out=16'h9f0;
17'h3551:	data_out=16'ha00;
17'h3552:	data_out=16'h8ea;
17'h3553:	data_out=16'h890f;
17'h3554:	data_out=16'h86bf;
17'h3555:	data_out=16'haa;
17'h3556:	data_out=16'ha00;
17'h3557:	data_out=16'h780;
17'h3558:	data_out=16'h879;
17'h3559:	data_out=16'h9ff;
17'h355a:	data_out=16'h88bf;
17'h355b:	data_out=16'h8697;
17'h355c:	data_out=16'h89a4;
17'h355d:	data_out=16'h99e;
17'h355e:	data_out=16'h84fa;
17'h355f:	data_out=16'h218;
17'h3560:	data_out=16'h89fb;
17'h3561:	data_out=16'h864d;
17'h3562:	data_out=16'h21;
17'h3563:	data_out=16'h8a00;
17'h3564:	data_out=16'h8a00;
17'h3565:	data_out=16'h9fa;
17'h3566:	data_out=16'h6de;
17'h3567:	data_out=16'h8a00;
17'h3568:	data_out=16'h2c5;
17'h3569:	data_out=16'h8318;
17'h356a:	data_out=16'h2d2;
17'h356b:	data_out=16'h9fd;
17'h356c:	data_out=16'h160;
17'h356d:	data_out=16'h8a00;
17'h356e:	data_out=16'h2d3;
17'h356f:	data_out=16'h9ff;
17'h3570:	data_out=16'h2d1;
17'h3571:	data_out=16'h9fd;
17'h3572:	data_out=16'h84c;
17'h3573:	data_out=16'h9ff;
17'h3574:	data_out=16'ha00;
17'h3575:	data_out=16'h82d8;
17'h3576:	data_out=16'h8a00;
17'h3577:	data_out=16'h9fa;
17'h3578:	data_out=16'h8a7;
17'h3579:	data_out=16'h968;
17'h357a:	data_out=16'h8958;
17'h357b:	data_out=16'h2c4;
17'h357c:	data_out=16'h43a;
17'h357d:	data_out=16'h78a;
17'h357e:	data_out=16'h8a00;
17'h357f:	data_out=16'ha00;
17'h3580:	data_out=16'h897d;
17'h3581:	data_out=16'h89fc;
17'h3582:	data_out=16'h74;
17'h3583:	data_out=16'h812e;
17'h3584:	data_out=16'h9b0;
17'h3585:	data_out=16'h5d1;
17'h3586:	data_out=16'h212;
17'h3587:	data_out=16'h43c;
17'h3588:	data_out=16'h8740;
17'h3589:	data_out=16'h8609;
17'h358a:	data_out=16'h89fe;
17'h358b:	data_out=16'h8a00;
17'h358c:	data_out=16'h9f6;
17'h358d:	data_out=16'h149;
17'h358e:	data_out=16'h59;
17'h358f:	data_out=16'h8040;
17'h3590:	data_out=16'h86eb;
17'h3591:	data_out=16'h53a;
17'h3592:	data_out=16'h8954;
17'h3593:	data_out=16'h31;
17'h3594:	data_out=16'h89fa;
17'h3595:	data_out=16'h81eb;
17'h3596:	data_out=16'h8190;
17'h3597:	data_out=16'h89f4;
17'h3598:	data_out=16'h23;
17'h3599:	data_out=16'h9fe;
17'h359a:	data_out=16'ha00;
17'h359b:	data_out=16'h88c5;
17'h359c:	data_out=16'h88b4;
17'h359d:	data_out=16'h89f1;
17'h359e:	data_out=16'h891f;
17'h359f:	data_out=16'h506;
17'h35a0:	data_out=16'h89fd;
17'h35a1:	data_out=16'h5f;
17'h35a2:	data_out=16'hf2;
17'h35a3:	data_out=16'h200;
17'h35a4:	data_out=16'h201;
17'h35a5:	data_out=16'h9ff;
17'h35a6:	data_out=16'h8852;
17'h35a7:	data_out=16'h89ff;
17'h35a8:	data_out=16'h61;
17'h35a9:	data_out=16'h8964;
17'h35aa:	data_out=16'h8632;
17'h35ab:	data_out=16'h8a00;
17'h35ac:	data_out=16'h81fb;
17'h35ad:	data_out=16'h8595;
17'h35ae:	data_out=16'h8441;
17'h35af:	data_out=16'h88de;
17'h35b0:	data_out=16'ha00;
17'h35b1:	data_out=16'h89ff;
17'h35b2:	data_out=16'ha00;
17'h35b3:	data_out=16'h89ff;
17'h35b4:	data_out=16'h8a00;
17'h35b5:	data_out=16'h9db;
17'h35b6:	data_out=16'h8861;
17'h35b7:	data_out=16'h8047;
17'h35b8:	data_out=16'h885d;
17'h35b9:	data_out=16'h89fe;
17'h35ba:	data_out=16'h883d;
17'h35bb:	data_out=16'h856e;
17'h35bc:	data_out=16'h8864;
17'h35bd:	data_out=16'h8887;
17'h35be:	data_out=16'h60;
17'h35bf:	data_out=16'h5cf;
17'h35c0:	data_out=16'ha00;
17'h35c1:	data_out=16'h80cc;
17'h35c2:	data_out=16'h9fa;
17'h35c3:	data_out=16'h38a;
17'h35c4:	data_out=16'h89e0;
17'h35c5:	data_out=16'h81f0;
17'h35c6:	data_out=16'h897c;
17'h35c7:	data_out=16'h8049;
17'h35c8:	data_out=16'h8408;
17'h35c9:	data_out=16'h9fe;
17'h35ca:	data_out=16'h9dd;
17'h35cb:	data_out=16'h993;
17'h35cc:	data_out=16'ha00;
17'h35cd:	data_out=16'h74;
17'h35ce:	data_out=16'h8642;
17'h35cf:	data_out=16'h922;
17'h35d0:	data_out=16'h9ea;
17'h35d1:	data_out=16'h19b;
17'h35d2:	data_out=16'h26c;
17'h35d3:	data_out=16'h89ef;
17'h35d4:	data_out=16'h89c7;
17'h35d5:	data_out=16'h8558;
17'h35d6:	data_out=16'h2e6;
17'h35d7:	data_out=16'h22c;
17'h35d8:	data_out=16'h82e6;
17'h35d9:	data_out=16'h9ff;
17'h35da:	data_out=16'h89f4;
17'h35db:	data_out=16'h89fc;
17'h35dc:	data_out=16'h89f1;
17'h35dd:	data_out=16'h220;
17'h35de:	data_out=16'h8796;
17'h35df:	data_out=16'h804e;
17'h35e0:	data_out=16'h89a4;
17'h35e1:	data_out=16'h892a;
17'h35e2:	data_out=16'h86c1;
17'h35e3:	data_out=16'h89ff;
17'h35e4:	data_out=16'h8a00;
17'h35e5:	data_out=16'h9f8;
17'h35e6:	data_out=16'h9e7;
17'h35e7:	data_out=16'h8a00;
17'h35e8:	data_out=16'h5f;
17'h35e9:	data_out=16'h8849;
17'h35ea:	data_out=16'h58;
17'h35eb:	data_out=16'ha00;
17'h35ec:	data_out=16'h8844;
17'h35ed:	data_out=16'h89ff;
17'h35ee:	data_out=16'h58;
17'h35ef:	data_out=16'ha00;
17'h35f0:	data_out=16'h59;
17'h35f1:	data_out=16'h81a0;
17'h35f2:	data_out=16'h2c2;
17'h35f3:	data_out=16'h500;
17'h35f4:	data_out=16'ha00;
17'h35f5:	data_out=16'h87bc;
17'h35f6:	data_out=16'h8a00;
17'h35f7:	data_out=16'h9fa;
17'h35f8:	data_out=16'h542;
17'h35f9:	data_out=16'h8437;
17'h35fa:	data_out=16'h89fb;
17'h35fb:	data_out=16'h61;
17'h35fc:	data_out=16'h7e;
17'h35fd:	data_out=16'h1a9;
17'h35fe:	data_out=16'h8966;
17'h35ff:	data_out=16'ha00;
17'h3600:	data_out=16'h89fc;
17'h3601:	data_out=16'h89fe;
17'h3602:	data_out=16'h8907;
17'h3603:	data_out=16'h833b;
17'h3604:	data_out=16'h9f9;
17'h3605:	data_out=16'h3c4;
17'h3606:	data_out=16'hde;
17'h3607:	data_out=16'h318;
17'h3608:	data_out=16'h89fe;
17'h3609:	data_out=16'h8211;
17'h360a:	data_out=16'h89ff;
17'h360b:	data_out=16'h8a00;
17'h360c:	data_out=16'h9fa;
17'h360d:	data_out=16'h84d7;
17'h360e:	data_out=16'h818c;
17'h360f:	data_out=16'h89c1;
17'h3610:	data_out=16'h8306;
17'h3611:	data_out=16'h4d8;
17'h3612:	data_out=16'h89ff;
17'h3613:	data_out=16'h844c;
17'h3614:	data_out=16'h8a00;
17'h3615:	data_out=16'h8320;
17'h3616:	data_out=16'h8589;
17'h3617:	data_out=16'h8a00;
17'h3618:	data_out=16'h8309;
17'h3619:	data_out=16'ha00;
17'h361a:	data_out=16'ha00;
17'h361b:	data_out=16'h8a00;
17'h361c:	data_out=16'h8a00;
17'h361d:	data_out=16'h89ff;
17'h361e:	data_out=16'h8a00;
17'h361f:	data_out=16'h817f;
17'h3620:	data_out=16'h89ff;
17'h3621:	data_out=16'h817c;
17'h3622:	data_out=16'h403;
17'h3623:	data_out=16'h804f;
17'h3624:	data_out=16'h804f;
17'h3625:	data_out=16'h93d;
17'h3626:	data_out=16'h89fe;
17'h3627:	data_out=16'h89ff;
17'h3628:	data_out=16'h816f;
17'h3629:	data_out=16'h89ff;
17'h362a:	data_out=16'h89ff;
17'h362b:	data_out=16'h8a00;
17'h362c:	data_out=16'h8462;
17'h362d:	data_out=16'h8405;
17'h362e:	data_out=16'h8a00;
17'h362f:	data_out=16'h8573;
17'h3630:	data_out=16'ha00;
17'h3631:	data_out=16'h89ff;
17'h3632:	data_out=16'ha00;
17'h3633:	data_out=16'h8a00;
17'h3634:	data_out=16'h86f1;
17'h3635:	data_out=16'h66c;
17'h3636:	data_out=16'h89fe;
17'h3637:	data_out=16'h891f;
17'h3638:	data_out=16'h88a7;
17'h3639:	data_out=16'h8a00;
17'h363a:	data_out=16'h84cc;
17'h363b:	data_out=16'h823b;
17'h363c:	data_out=16'h89fe;
17'h363d:	data_out=16'h8680;
17'h363e:	data_out=16'h816f;
17'h363f:	data_out=16'h3c2;
17'h3640:	data_out=16'ha00;
17'h3641:	data_out=16'h86d2;
17'h3642:	data_out=16'h9fc;
17'h3643:	data_out=16'h219;
17'h3644:	data_out=16'h86bc;
17'h3645:	data_out=16'h8339;
17'h3646:	data_out=16'h89fb;
17'h3647:	data_out=16'h818d;
17'h3648:	data_out=16'h8530;
17'h3649:	data_out=16'h95f;
17'h364a:	data_out=16'h778;
17'h364b:	data_out=16'h9f8;
17'h364c:	data_out=16'h979;
17'h364d:	data_out=16'h41b;
17'h364e:	data_out=16'h89fe;
17'h364f:	data_out=16'h6d4;
17'h3650:	data_out=16'h820;
17'h3651:	data_out=16'h86a1;
17'h3652:	data_out=16'h800a;
17'h3653:	data_out=16'h8a00;
17'h3654:	data_out=16'h8983;
17'h3655:	data_out=16'h8a00;
17'h3656:	data_out=16'h854f;
17'h3657:	data_out=16'h8459;
17'h3658:	data_out=16'h89fe;
17'h3659:	data_out=16'h7ce;
17'h365a:	data_out=16'h8a00;
17'h365b:	data_out=16'h89fe;
17'h365c:	data_out=16'h8696;
17'h365d:	data_out=16'h82ef;
17'h365e:	data_out=16'h846d;
17'h365f:	data_out=16'h8284;
17'h3660:	data_out=16'h8a00;
17'h3661:	data_out=16'h89da;
17'h3662:	data_out=16'h8a00;
17'h3663:	data_out=16'h8a00;
17'h3664:	data_out=16'h89b0;
17'h3665:	data_out=16'ha00;
17'h3666:	data_out=16'h9f8;
17'h3667:	data_out=16'h8a00;
17'h3668:	data_out=16'h8175;
17'h3669:	data_out=16'h89fe;
17'h366a:	data_out=16'h8197;
17'h366b:	data_out=16'h874;
17'h366c:	data_out=16'h89fb;
17'h366d:	data_out=16'h8a00;
17'h366e:	data_out=16'h8196;
17'h366f:	data_out=16'h80d;
17'h3670:	data_out=16'h8190;
17'h3671:	data_out=16'h8a00;
17'h3672:	data_out=16'h801d;
17'h3673:	data_out=16'h360;
17'h3674:	data_out=16'ha00;
17'h3675:	data_out=16'h89fe;
17'h3676:	data_out=16'h8a00;
17'h3677:	data_out=16'h6d0;
17'h3678:	data_out=16'h5e5;
17'h3679:	data_out=16'h89fb;
17'h367a:	data_out=16'h8a00;
17'h367b:	data_out=16'h816f;
17'h367c:	data_out=16'h8294;
17'h367d:	data_out=16'h8052;
17'h367e:	data_out=16'h857f;
17'h367f:	data_out=16'h84b;
17'h3680:	data_out=16'h80e8;
17'h3681:	data_out=16'h803a;
17'h3682:	data_out=16'h80f1;
17'h3683:	data_out=16'h80e8;
17'h3684:	data_out=16'h15f;
17'h3685:	data_out=16'h116;
17'h3686:	data_out=16'h80b7;
17'h3687:	data_out=16'h8192;
17'h3688:	data_out=16'h810d;
17'h3689:	data_out=16'h80ed;
17'h368a:	data_out=16'h8088;
17'h368b:	data_out=16'h8336;
17'h368c:	data_out=16'h190;
17'h368d:	data_out=16'h8096;
17'h368e:	data_out=16'h802f;
17'h368f:	data_out=16'h8122;
17'h3690:	data_out=16'h805b;
17'h3691:	data_out=16'h119;
17'h3692:	data_out=16'h83a8;
17'h3693:	data_out=16'h12;
17'h3694:	data_out=16'h81fd;
17'h3695:	data_out=16'h9a;
17'h3696:	data_out=16'h32;
17'h3697:	data_out=16'h827c;
17'h3698:	data_out=16'h8017;
17'h3699:	data_out=16'h2d9;
17'h369a:	data_out=16'h1f7;
17'h369b:	data_out=16'h8255;
17'h369c:	data_out=16'h36;
17'h369d:	data_out=16'h80bf;
17'h369e:	data_out=16'h8200;
17'h369f:	data_out=16'h3a;
17'h36a0:	data_out=16'h81;
17'h36a1:	data_out=16'h8036;
17'h36a2:	data_out=16'h80ce;
17'h36a3:	data_out=16'h80c4;
17'h36a4:	data_out=16'h80d7;
17'h36a5:	data_out=16'h803a;
17'h36a6:	data_out=16'h8385;
17'h36a7:	data_out=16'h80fd;
17'h36a8:	data_out=16'h8034;
17'h36a9:	data_out=16'h80f3;
17'h36aa:	data_out=16'h82f1;
17'h36ab:	data_out=16'h823b;
17'h36ac:	data_out=16'h8008;
17'h36ad:	data_out=16'h8149;
17'h36ae:	data_out=16'h8161;
17'h36af:	data_out=16'h80b0;
17'h36b0:	data_out=16'h1db;
17'h36b1:	data_out=16'h806a;
17'h36b2:	data_out=16'h1ec;
17'h36b3:	data_out=16'h819c;
17'h36b4:	data_out=16'h7b;
17'h36b5:	data_out=16'h25a;
17'h36b6:	data_out=16'h80a9;
17'h36b7:	data_out=16'h8102;
17'h36b8:	data_out=16'h261;
17'h36b9:	data_out=16'h819a;
17'h36ba:	data_out=16'h81aa;
17'h36bb:	data_out=16'h67;
17'h36bc:	data_out=16'h810e;
17'h36bd:	data_out=16'ha4;
17'h36be:	data_out=16'h8035;
17'h36bf:	data_out=16'h288;
17'h36c0:	data_out=16'h70;
17'h36c1:	data_out=16'h8030;
17'h36c2:	data_out=16'hd1;
17'h36c3:	data_out=16'h3d;
17'h36c4:	data_out=16'h1a8;
17'h36c5:	data_out=16'h1e;
17'h36c6:	data_out=16'h8282;
17'h36c7:	data_out=16'h81f3;
17'h36c8:	data_out=16'h81cc;
17'h36c9:	data_out=16'h801c;
17'h36ca:	data_out=16'h7f;
17'h36cb:	data_out=16'h3c;
17'h36cc:	data_out=16'h7;
17'h36cd:	data_out=16'h80b6;
17'h36ce:	data_out=16'h8060;
17'h36cf:	data_out=16'h8028;
17'h36d0:	data_out=16'h95;
17'h36d1:	data_out=16'hb6;
17'h36d2:	data_out=16'h80d6;
17'h36d3:	data_out=16'h81d3;
17'h36d4:	data_out=16'h39;
17'h36d5:	data_out=16'h8061;
17'h36d6:	data_out=16'h8143;
17'h36d7:	data_out=16'h811c;
17'h36d8:	data_out=16'h80b6;
17'h36d9:	data_out=16'h80c5;
17'h36da:	data_out=16'h82e7;
17'h36db:	data_out=16'h122;
17'h36dc:	data_out=16'h4a;
17'h36dd:	data_out=16'h8094;
17'h36de:	data_out=16'h8007;
17'h36df:	data_out=16'h8045;
17'h36e0:	data_out=16'h827c;
17'h36e1:	data_out=16'h1e8;
17'h36e2:	data_out=16'h8333;
17'h36e3:	data_out=16'h81a6;
17'h36e4:	data_out=16'h805f;
17'h36e5:	data_out=16'h1a0;
17'h36e6:	data_out=16'h1b8;
17'h36e7:	data_out=16'h82f1;
17'h36e8:	data_out=16'h8035;
17'h36e9:	data_out=16'h8111;
17'h36ea:	data_out=16'h803c;
17'h36eb:	data_out=16'h10e;
17'h36ec:	data_out=16'h81a5;
17'h36ed:	data_out=16'h81a0;
17'h36ee:	data_out=16'h8031;
17'h36ef:	data_out=16'h8078;
17'h36f0:	data_out=16'h8036;
17'h36f1:	data_out=16'h8118;
17'h36f2:	data_out=16'h4c;
17'h36f3:	data_out=16'h106;
17'h36f4:	data_out=16'h1db;
17'h36f5:	data_out=16'h808c;
17'h36f6:	data_out=16'h834d;
17'h36f7:	data_out=16'h1b1;
17'h36f8:	data_out=16'h80be;
17'h36f9:	data_out=16'h8153;
17'h36fa:	data_out=16'h81db;
17'h36fb:	data_out=16'h803b;
17'h36fc:	data_out=16'h8085;
17'h36fd:	data_out=16'h80e3;
17'h36fe:	data_out=16'h814f;
17'h36ff:	data_out=16'h18f;
17'h3700:	data_out=16'h822a;
17'h3701:	data_out=16'h8227;
17'h3702:	data_out=16'h81c3;
17'h3703:	data_out=16'h80c4;
17'h3704:	data_out=16'h17e;
17'h3705:	data_out=16'h11;
17'h3706:	data_out=16'hb;
17'h3707:	data_out=16'h10e;
17'h3708:	data_out=16'h8253;
17'h3709:	data_out=16'h8017;
17'h370a:	data_out=16'h81d8;
17'h370b:	data_out=16'h815e;
17'h370c:	data_out=16'h33b;
17'h370d:	data_out=16'h8051;
17'h370e:	data_out=16'h8055;
17'h370f:	data_out=16'h817d;
17'h3710:	data_out=16'h8044;
17'h3711:	data_out=16'h5f;
17'h3712:	data_out=16'h819b;
17'h3713:	data_out=16'h802a;
17'h3714:	data_out=16'h827c;
17'h3715:	data_out=16'h807d;
17'h3716:	data_out=16'h80d8;
17'h3717:	data_out=16'h8274;
17'h3718:	data_out=16'h8057;
17'h3719:	data_out=16'h270;
17'h371a:	data_out=16'h174;
17'h371b:	data_out=16'h81bb;
17'h371c:	data_out=16'h81df;
17'h371d:	data_out=16'h8258;
17'h371e:	data_out=16'h825b;
17'h371f:	data_out=16'h8077;
17'h3720:	data_out=16'h81a4;
17'h3721:	data_out=16'h8057;
17'h3722:	data_out=16'h1c;
17'h3723:	data_out=16'h807a;
17'h3724:	data_out=16'h807f;
17'h3725:	data_out=16'h17d;
17'h3726:	data_out=16'h829b;
17'h3727:	data_out=16'h8260;
17'h3728:	data_out=16'h8049;
17'h3729:	data_out=16'h810f;
17'h372a:	data_out=16'h8212;
17'h372b:	data_out=16'h8223;
17'h372c:	data_out=16'h809c;
17'h372d:	data_out=16'h8031;
17'h372e:	data_out=16'h81b5;
17'h372f:	data_out=16'h80fe;
17'h3730:	data_out=16'h12d;
17'h3731:	data_out=16'h81f2;
17'h3732:	data_out=16'h13d;
17'h3733:	data_out=16'h825d;
17'h3734:	data_out=16'h8111;
17'h3735:	data_out=16'h1b1;
17'h3736:	data_out=16'h81a0;
17'h3737:	data_out=16'h81c9;
17'h3738:	data_out=16'h818d;
17'h3739:	data_out=16'h8256;
17'h373a:	data_out=16'h8049;
17'h373b:	data_out=16'h8067;
17'h373c:	data_out=16'h8235;
17'h373d:	data_out=16'h81ae;
17'h373e:	data_out=16'h8049;
17'h373f:	data_out=16'h114;
17'h3740:	data_out=16'h156;
17'h3741:	data_out=16'h8149;
17'h3742:	data_out=16'h2df;
17'h3743:	data_out=16'h61;
17'h3744:	data_out=16'h8077;
17'h3745:	data_out=16'h80c1;
17'h3746:	data_out=16'h82a1;
17'h3747:	data_out=16'h8036;
17'h3748:	data_out=16'h80b2;
17'h3749:	data_out=16'h173;
17'h374a:	data_out=16'h1d4;
17'h374b:	data_out=16'h399;
17'h374c:	data_out=16'h246;
17'h374d:	data_out=16'h27;
17'h374e:	data_out=16'h80be;
17'h374f:	data_out=16'h215;
17'h3750:	data_out=16'hd4;
17'h3751:	data_out=16'h813e;
17'h3752:	data_out=16'h8060;
17'h3753:	data_out=16'h8249;
17'h3754:	data_out=16'h8162;
17'h3755:	data_out=16'h81cd;
17'h3756:	data_out=16'h819c;
17'h3757:	data_out=16'h811b;
17'h3758:	data_out=16'h8234;
17'h3759:	data_out=16'h4c;
17'h375a:	data_out=16'h826a;
17'h375b:	data_out=16'h8230;
17'h375c:	data_out=16'h80eb;
17'h375d:	data_out=16'h80de;
17'h375e:	data_out=16'h808c;
17'h375f:	data_out=16'h8065;
17'h3760:	data_out=16'h81b6;
17'h3761:	data_out=16'h80d6;
17'h3762:	data_out=16'h81ec;
17'h3763:	data_out=16'h823b;
17'h3764:	data_out=16'h8133;
17'h3765:	data_out=16'h291;
17'h3766:	data_out=16'h2a9;
17'h3767:	data_out=16'h81a7;
17'h3768:	data_out=16'h8050;
17'h3769:	data_out=16'h8212;
17'h376a:	data_out=16'h805b;
17'h376b:	data_out=16'hc3;
17'h376c:	data_out=16'h824c;
17'h376d:	data_out=16'h8267;
17'h376e:	data_out=16'h804e;
17'h376f:	data_out=16'h12;
17'h3770:	data_out=16'h805a;
17'h3771:	data_out=16'h81b3;
17'h3772:	data_out=16'h808f;
17'h3773:	data_out=16'h8032;
17'h3774:	data_out=16'h128;
17'h3775:	data_out=16'h8153;
17'h3776:	data_out=16'h824c;
17'h3777:	data_out=16'h1b3;
17'h3778:	data_out=16'h38;
17'h3779:	data_out=16'h81ff;
17'h377a:	data_out=16'h8266;
17'h377b:	data_out=16'h8050;
17'h377c:	data_out=16'h80b0;
17'h377d:	data_out=16'h800c;
17'h377e:	data_out=16'h80b9;
17'h377f:	data_out=16'h11c;
17'h3780:	data_out=16'h8004;
17'h3781:	data_out=16'h7;
17'h3782:	data_out=16'h8005;
17'h3783:	data_out=16'h4;
17'h3784:	data_out=16'h3;
17'h3785:	data_out=16'h8;
17'h3786:	data_out=16'h8005;
17'h3787:	data_out=16'h7;
17'h3788:	data_out=16'h8003;
17'h3789:	data_out=16'h8000;
17'h378a:	data_out=16'h2;
17'h378b:	data_out=16'h4;
17'h378c:	data_out=16'h2;
17'h378d:	data_out=16'h1;
17'h378e:	data_out=16'h5;
17'h378f:	data_out=16'h4;
17'h3790:	data_out=16'h8003;
17'h3791:	data_out=16'h2;
17'h3792:	data_out=16'h5;
17'h3793:	data_out=16'h8;
17'h3794:	data_out=16'h8;
17'h3795:	data_out=16'h8006;
17'h3796:	data_out=16'h4;
17'h3797:	data_out=16'h0;
17'h3798:	data_out=16'h8008;
17'h3799:	data_out=16'h8001;
17'h379a:	data_out=16'h1;
17'h379b:	data_out=16'h8;
17'h379c:	data_out=16'h8000;
17'h379d:	data_out=16'h8004;
17'h379e:	data_out=16'h3;
17'h379f:	data_out=16'h5;
17'h37a0:	data_out=16'h8007;
17'h37a1:	data_out=16'h8;
17'h37a2:	data_out=16'h0;
17'h37a3:	data_out=16'h5;
17'h37a4:	data_out=16'h6;
17'h37a5:	data_out=16'h5;
17'h37a6:	data_out=16'h3;
17'h37a7:	data_out=16'h8006;
17'h37a8:	data_out=16'h8005;
17'h37a9:	data_out=16'h8004;
17'h37aa:	data_out=16'h7;
17'h37ab:	data_out=16'h6;
17'h37ac:	data_out=16'h6;
17'h37ad:	data_out=16'h3;
17'h37ae:	data_out=16'h1;
17'h37af:	data_out=16'h8006;
17'h37b0:	data_out=16'h8004;
17'h37b1:	data_out=16'h8003;
17'h37b2:	data_out=16'h8008;
17'h37b3:	data_out=16'h8005;
17'h37b4:	data_out=16'h8000;
17'h37b5:	data_out=16'h5;
17'h37b6:	data_out=16'h4;
17'h37b7:	data_out=16'h1;
17'h37b8:	data_out=16'h8005;
17'h37b9:	data_out=16'h8004;
17'h37ba:	data_out=16'h8000;
17'h37bb:	data_out=16'h4;
17'h37bc:	data_out=16'h2;
17'h37bd:	data_out=16'h8006;
17'h37be:	data_out=16'h0;
17'h37bf:	data_out=16'h4;
17'h37c0:	data_out=16'h8008;
17'h37c1:	data_out=16'h8009;
17'h37c2:	data_out=16'h0;
17'h37c3:	data_out=16'h8;
17'h37c4:	data_out=16'h5;
17'h37c5:	data_out=16'h8006;
17'h37c6:	data_out=16'h8007;
17'h37c7:	data_out=16'h8009;
17'h37c8:	data_out=16'h8001;
17'h37c9:	data_out=16'h9;
17'h37ca:	data_out=16'h6;
17'h37cb:	data_out=16'h8005;
17'h37cc:	data_out=16'h3;
17'h37cd:	data_out=16'h8002;
17'h37ce:	data_out=16'h8002;
17'h37cf:	data_out=16'h8;
17'h37d0:	data_out=16'h4;
17'h37d1:	data_out=16'h0;
17'h37d2:	data_out=16'h8007;
17'h37d3:	data_out=16'h8005;
17'h37d4:	data_out=16'h8004;
17'h37d5:	data_out=16'h6;
17'h37d6:	data_out=16'h5;
17'h37d7:	data_out=16'h0;
17'h37d8:	data_out=16'h8006;
17'h37d9:	data_out=16'h8005;
17'h37da:	data_out=16'h8005;
17'h37db:	data_out=16'h4;
17'h37dc:	data_out=16'h8002;
17'h37dd:	data_out=16'h4;
17'h37de:	data_out=16'h8001;
17'h37df:	data_out=16'h8000;
17'h37e0:	data_out=16'h4;
17'h37e1:	data_out=16'h9;
17'h37e2:	data_out=16'h8002;
17'h37e3:	data_out=16'h8000;
17'h37e4:	data_out=16'h8006;
17'h37e5:	data_out=16'h8000;
17'h37e6:	data_out=16'h8000;
17'h37e7:	data_out=16'h2;
17'h37e8:	data_out=16'h8000;
17'h37e9:	data_out=16'h8003;
17'h37ea:	data_out=16'h6;
17'h37eb:	data_out=16'h8007;
17'h37ec:	data_out=16'h4;
17'h37ed:	data_out=16'h8005;
17'h37ee:	data_out=16'h8008;
17'h37ef:	data_out=16'h8001;
17'h37f0:	data_out=16'h5;
17'h37f1:	data_out=16'h8006;
17'h37f2:	data_out=16'h3;
17'h37f3:	data_out=16'h8008;
17'h37f4:	data_out=16'h8009;
17'h37f5:	data_out=16'h8002;
17'h37f6:	data_out=16'h1;
17'h37f7:	data_out=16'h8006;
17'h37f8:	data_out=16'h3;
17'h37f9:	data_out=16'h5;
17'h37fa:	data_out=16'h7;
17'h37fb:	data_out=16'h8009;
17'h37fc:	data_out=16'h8001;
17'h37fd:	data_out=16'h8002;
17'h37fe:	data_out=16'h0;
17'h37ff:	data_out=16'h8006;
17'h3800:	data_out=16'h8002;
17'h3801:	data_out=16'h7;
17'h3802:	data_out=16'h3;
17'h3803:	data_out=16'h0;
17'h3804:	data_out=16'h8002;
17'h3805:	data_out=16'h8006;
17'h3806:	data_out=16'h8007;
17'h3807:	data_out=16'h7;
17'h3808:	data_out=16'h8000;
17'h3809:	data_out=16'h8;
17'h380a:	data_out=16'h8009;
17'h380b:	data_out=16'h8005;
17'h380c:	data_out=16'h8005;
17'h380d:	data_out=16'h8008;
17'h380e:	data_out=16'h3;
17'h380f:	data_out=16'h8;
17'h3810:	data_out=16'h8005;
17'h3811:	data_out=16'h8003;
17'h3812:	data_out=16'h9;
17'h3813:	data_out=16'h8005;
17'h3814:	data_out=16'h5;
17'h3815:	data_out=16'h1;
17'h3816:	data_out=16'h8002;
17'h3817:	data_out=16'h8002;
17'h3818:	data_out=16'h8004;
17'h3819:	data_out=16'h8003;
17'h381a:	data_out=16'h8001;
17'h381b:	data_out=16'h5;
17'h381c:	data_out=16'h4;
17'h381d:	data_out=16'h8;
17'h381e:	data_out=16'h8;
17'h381f:	data_out=16'h8008;
17'h3820:	data_out=16'h6;
17'h3821:	data_out=16'h2;
17'h3822:	data_out=16'h2;
17'h3823:	data_out=16'h8005;
17'h3824:	data_out=16'h5;
17'h3825:	data_out=16'h4;
17'h3826:	data_out=16'h8007;
17'h3827:	data_out=16'h8004;
17'h3828:	data_out=16'h3;
17'h3829:	data_out=16'h8006;
17'h382a:	data_out=16'h8000;
17'h382b:	data_out=16'h7;
17'h382c:	data_out=16'h8005;
17'h382d:	data_out=16'h8006;
17'h382e:	data_out=16'h6;
17'h382f:	data_out=16'h8001;
17'h3830:	data_out=16'h8000;
17'h3831:	data_out=16'h6;
17'h3832:	data_out=16'h3;
17'h3833:	data_out=16'h8005;
17'h3834:	data_out=16'h8003;
17'h3835:	data_out=16'h8007;
17'h3836:	data_out=16'h3;
17'h3837:	data_out=16'h2;
17'h3838:	data_out=16'h8001;
17'h3839:	data_out=16'h8007;
17'h383a:	data_out=16'h8002;
17'h383b:	data_out=16'h8007;
17'h383c:	data_out=16'h8009;
17'h383d:	data_out=16'h8004;
17'h383e:	data_out=16'h8005;
17'h383f:	data_out=16'h7;
17'h3840:	data_out=16'h8;
17'h3841:	data_out=16'h6;
17'h3842:	data_out=16'h8007;
17'h3843:	data_out=16'h3;
17'h3844:	data_out=16'h0;
17'h3845:	data_out=16'h8004;
17'h3846:	data_out=16'h8;
17'h3847:	data_out=16'h8006;
17'h3848:	data_out=16'h8001;
17'h3849:	data_out=16'h8002;
17'h384a:	data_out=16'h8009;
17'h384b:	data_out=16'h3;
17'h384c:	data_out=16'h1;
17'h384d:	data_out=16'h6;
17'h384e:	data_out=16'h8008;
17'h384f:	data_out=16'h8008;
17'h3850:	data_out=16'h3;
17'h3851:	data_out=16'h5;
17'h3852:	data_out=16'h8003;
17'h3853:	data_out=16'h9;
17'h3854:	data_out=16'h7;
17'h3855:	data_out=16'h9;
17'h3856:	data_out=16'h2;
17'h3857:	data_out=16'h8004;
17'h3858:	data_out=16'h8008;
17'h3859:	data_out=16'h8009;
17'h385a:	data_out=16'h8001;
17'h385b:	data_out=16'h8007;
17'h385c:	data_out=16'h8003;
17'h385d:	data_out=16'h3;
17'h385e:	data_out=16'h9;
17'h385f:	data_out=16'h8005;
17'h3860:	data_out=16'h8001;
17'h3861:	data_out=16'h8007;
17'h3862:	data_out=16'h7;
17'h3863:	data_out=16'h9;
17'h3864:	data_out=16'h8002;
17'h3865:	data_out=16'h6;
17'h3866:	data_out=16'h8007;
17'h3867:	data_out=16'h6;
17'h3868:	data_out=16'h8004;
17'h3869:	data_out=16'h8006;
17'h386a:	data_out=16'h8001;
17'h386b:	data_out=16'h6;
17'h386c:	data_out=16'h8009;
17'h386d:	data_out=16'h1;
17'h386e:	data_out=16'h7;
17'h386f:	data_out=16'h3;
17'h3870:	data_out=16'h8003;
17'h3871:	data_out=16'h8005;
17'h3872:	data_out=16'h3;
17'h3873:	data_out=16'h8006;
17'h3874:	data_out=16'h8006;
17'h3875:	data_out=16'h8004;
17'h3876:	data_out=16'h0;
17'h3877:	data_out=16'h8004;
17'h3878:	data_out=16'h8003;
17'h3879:	data_out=16'h8;
17'h387a:	data_out=16'h8003;
17'h387b:	data_out=16'h2;
17'h387c:	data_out=16'h2;
17'h387d:	data_out=16'h8003;
17'h387e:	data_out=16'h6;
17'h387f:	data_out=16'h8008;
17'h3880:	data_out=16'h8003;
17'h3881:	data_out=16'h9;
17'h3882:	data_out=16'h4;
17'h3883:	data_out=16'hf;
17'h3884:	data_out=16'h5;
17'h3885:	data_out=16'h8001;
17'h3886:	data_out=16'h9;
17'h3887:	data_out=16'h10;
17'h3888:	data_out=16'h5;
17'h3889:	data_out=16'h8005;
17'h388a:	data_out=16'h9;
17'h388b:	data_out=16'h9;
17'h388c:	data_out=16'hc;
17'h388d:	data_out=16'ha;
17'h388e:	data_out=16'h8005;
17'h388f:	data_out=16'h13;
17'h3890:	data_out=16'hc;
17'h3891:	data_out=16'h8;
17'h3892:	data_out=16'h8;
17'h3893:	data_out=16'h15;
17'h3894:	data_out=16'h4;
17'h3895:	data_out=16'h5;
17'h3896:	data_out=16'h1;
17'h3897:	data_out=16'hd;
17'h3898:	data_out=16'h8;
17'h3899:	data_out=16'h3;
17'h389a:	data_out=16'hd;
17'h389b:	data_out=16'h5;
17'h389c:	data_out=16'hc;
17'h389d:	data_out=16'hc;
17'h389e:	data_out=16'h6;
17'h389f:	data_out=16'h5;
17'h38a0:	data_out=16'h1;
17'h38a1:	data_out=16'h8001;
17'h38a2:	data_out=16'h8000;
17'h38a3:	data_out=16'h8004;
17'h38a4:	data_out=16'h2;
17'h38a5:	data_out=16'he;
17'h38a6:	data_out=16'h8000;
17'h38a7:	data_out=16'hb;
17'h38a8:	data_out=16'hc;
17'h38a9:	data_out=16'h10;
17'h38aa:	data_out=16'h9;
17'h38ab:	data_out=16'h6;
17'h38ac:	data_out=16'h2;
17'h38ad:	data_out=16'h4;
17'h38ae:	data_out=16'h13;
17'h38af:	data_out=16'h8001;
17'h38b0:	data_out=16'h12;
17'h38b1:	data_out=16'h9;
17'h38b2:	data_out=16'h2;
17'h38b3:	data_out=16'h13;
17'h38b4:	data_out=16'h5;
17'h38b5:	data_out=16'h5;
17'h38b6:	data_out=16'h5;
17'h38b7:	data_out=16'h8;
17'h38b8:	data_out=16'h9;
17'h38b9:	data_out=16'h3;
17'h38ba:	data_out=16'h4;
17'h38bb:	data_out=16'ha;
17'h38bc:	data_out=16'h8;
17'h38bd:	data_out=16'h2;
17'h38be:	data_out=16'h8001;
17'h38bf:	data_out=16'h9;
17'h38c0:	data_out=16'h8002;
17'h38c1:	data_out=16'hb;
17'h38c2:	data_out=16'h12;
17'h38c3:	data_out=16'h5;
17'h38c4:	data_out=16'h4;
17'h38c5:	data_out=16'h8;
17'h38c6:	data_out=16'h4;
17'h38c7:	data_out=16'h5;
17'h38c8:	data_out=16'hf;
17'h38c9:	data_out=16'h6;
17'h38ca:	data_out=16'h3;
17'h38cb:	data_out=16'h16;
17'h38cc:	data_out=16'hf;
17'h38cd:	data_out=16'h6;
17'h38ce:	data_out=16'h2;
17'h38cf:	data_out=16'hd;
17'h38d0:	data_out=16'h7;
17'h38d1:	data_out=16'h1;
17'h38d2:	data_out=16'h4;
17'h38d3:	data_out=16'h8001;
17'h38d4:	data_out=16'h4;
17'h38d5:	data_out=16'h15;
17'h38d6:	data_out=16'h6;
17'h38d7:	data_out=16'h6;
17'h38d8:	data_out=16'h8;
17'h38d9:	data_out=16'h9;
17'h38da:	data_out=16'h9;
17'h38db:	data_out=16'h8001;
17'h38dc:	data_out=16'h5;
17'h38dd:	data_out=16'hb;
17'h38de:	data_out=16'h12;
17'h38df:	data_out=16'h5;
17'h38e0:	data_out=16'h4;
17'h38e1:	data_out=16'hb;
17'h38e2:	data_out=16'h13;
17'h38e3:	data_out=16'ha;
17'h38e4:	data_out=16'h6;
17'h38e5:	data_out=16'h2;
17'h38e6:	data_out=16'h9;
17'h38e7:	data_out=16'h6;
17'h38e8:	data_out=16'h7;
17'h38e9:	data_out=16'h12;
17'h38ea:	data_out=16'h8003;
17'h38eb:	data_out=16'h1;
17'h38ec:	data_out=16'h8;
17'h38ed:	data_out=16'h4;
17'h38ee:	data_out=16'h8005;
17'h38ef:	data_out=16'h8000;
17'h38f0:	data_out=16'h8001;
17'h38f1:	data_out=16'h12;
17'h38f2:	data_out=16'h1;
17'h38f3:	data_out=16'h9;
17'h38f4:	data_out=16'hc;
17'h38f5:	data_out=16'ha;
17'h38f6:	data_out=16'h8003;
17'h38f7:	data_out=16'hf;
17'h38f8:	data_out=16'h8003;
17'h38f9:	data_out=16'h12;
17'h38fa:	data_out=16'h7;
17'h38fb:	data_out=16'h4;
17'h38fc:	data_out=16'h8002;
17'h38fd:	data_out=16'h8002;
17'h38fe:	data_out=16'he;
17'h38ff:	data_out=16'h1;
17'h3900:	data_out=16'h802f;
17'h3901:	data_out=16'h38;
17'h3902:	data_out=16'h7;
17'h3903:	data_out=16'hd;
17'h3904:	data_out=16'h8033;
17'h3905:	data_out=16'ha;
17'h3906:	data_out=16'h5;
17'h3907:	data_out=16'h8009;
17'h3908:	data_out=16'h800c;
17'h3909:	data_out=16'h805e;
17'h390a:	data_out=16'h1;
17'h390b:	data_out=16'h6e;
17'h390c:	data_out=16'h8053;
17'h390d:	data_out=16'h28;
17'h390e:	data_out=16'hd;
17'h390f:	data_out=16'h48;
17'h3910:	data_out=16'h803b;
17'h3911:	data_out=16'h8029;
17'h3912:	data_out=16'h3d;
17'h3913:	data_out=16'h2d;
17'h3914:	data_out=16'h9e;
17'h3915:	data_out=16'h24;
17'h3916:	data_out=16'h29;
17'h3917:	data_out=16'hb1;
17'h3918:	data_out=16'h8028;
17'h3919:	data_out=16'h805b;
17'h391a:	data_out=16'h802f;
17'h391b:	data_out=16'h5e;
17'h391c:	data_out=16'h31;
17'h391d:	data_out=16'h13;
17'h391e:	data_out=16'h53;
17'h391f:	data_out=16'h28;
17'h3920:	data_out=16'h1f;
17'h3921:	data_out=16'h1;
17'h3922:	data_out=16'h8018;
17'h3923:	data_out=16'h8034;
17'h3924:	data_out=16'h802a;
17'h3925:	data_out=16'h802d;
17'h3926:	data_out=16'h801f;
17'h3927:	data_out=16'h1b;
17'h3928:	data_out=16'hd;
17'h3929:	data_out=16'h2f;
17'h392a:	data_out=16'h8007;
17'h392b:	data_out=16'h802d;
17'h392c:	data_out=16'h2f;
17'h392d:	data_out=16'h8022;
17'h392e:	data_out=16'h1c;
17'h392f:	data_out=16'h30;
17'h3930:	data_out=16'h1d;
17'h3931:	data_out=16'h0;
17'h3932:	data_out=16'h29;
17'h3933:	data_out=16'h8d;
17'h3934:	data_out=16'h800a;
17'h3935:	data_out=16'h8021;
17'h3936:	data_out=16'h28;
17'h3937:	data_out=16'h19;
17'h3938:	data_out=16'h8018;
17'h3939:	data_out=16'h60;
17'h393a:	data_out=16'h803a;
17'h393b:	data_out=16'h801f;
17'h393c:	data_out=16'h2c;
17'h393d:	data_out=16'h8025;
17'h393e:	data_out=16'h2;
17'h393f:	data_out=16'h8000;
17'h3940:	data_out=16'h802d;
17'h3941:	data_out=16'h29;
17'h3942:	data_out=16'h8044;
17'h3943:	data_out=16'h8004;
17'h3944:	data_out=16'h8001;
17'h3945:	data_out=16'h8006;
17'h3946:	data_out=16'h3a;
17'h3947:	data_out=16'h802d;
17'h3948:	data_out=16'h8004;
17'h3949:	data_out=16'h8041;
17'h394a:	data_out=16'h8012;
17'h394b:	data_out=16'h803f;
17'h394c:	data_out=16'h8043;
17'h394d:	data_out=16'h8008;
17'h394e:	data_out=16'h5;
17'h394f:	data_out=16'h8045;
17'h3950:	data_out=16'h802c;
17'h3951:	data_out=16'h53;
17'h3952:	data_out=16'h801a;
17'h3953:	data_out=16'h4d;
17'h3954:	data_out=16'h49;
17'h3955:	data_out=16'h32;
17'h3956:	data_out=16'h43;
17'h3957:	data_out=16'h801a;
17'h3958:	data_out=16'hb;
17'h3959:	data_out=16'h802e;
17'h395a:	data_out=16'h35;
17'h395b:	data_out=16'h6b;
17'h395c:	data_out=16'h17;
17'h395d:	data_out=16'h0;
17'h395e:	data_out=16'h32;
17'h395f:	data_out=16'h8018;
17'h3960:	data_out=16'h800d;
17'h3961:	data_out=16'h3d;
17'h3962:	data_out=16'h59;
17'h3963:	data_out=16'h91;
17'h3964:	data_out=16'h801b;
17'h3965:	data_out=16'h8030;
17'h3966:	data_out=16'h8051;
17'h3967:	data_out=16'h800d;
17'h3968:	data_out=16'h7;
17'h3969:	data_out=16'h10;
17'h396a:	data_out=16'h2;
17'h396b:	data_out=16'h801a;
17'h396c:	data_out=16'h6;
17'h396d:	data_out=16'h88;
17'h396e:	data_out=16'h4;
17'h396f:	data_out=16'h15;
17'h3970:	data_out=16'h8001;
17'h3971:	data_out=16'h9;
17'h3972:	data_out=16'h800a;
17'h3973:	data_out=16'h14;
17'h3974:	data_out=16'h1d;
17'h3975:	data_out=16'h28;
17'h3976:	data_out=16'h8010;
17'h3977:	data_out=16'h8046;
17'h3978:	data_out=16'h7;
17'h3979:	data_out=16'h19;
17'h397a:	data_out=16'ha4;
17'h397b:	data_out=16'h4;
17'h397c:	data_out=16'h11;
17'h397d:	data_out=16'h42;
17'h397e:	data_out=16'h803b;
17'h397f:	data_out=16'h8024;
17'h3980:	data_out=16'h807a;
17'h3981:	data_out=16'h68;
17'h3982:	data_out=16'ha2;
17'h3983:	data_out=16'h2e;
17'h3984:	data_out=16'h7f;
17'h3985:	data_out=16'hf2;
17'h3986:	data_out=16'h801e;
17'h3987:	data_out=16'h8051;
17'h3988:	data_out=16'h26;
17'h3989:	data_out=16'h80e1;
17'h398a:	data_out=16'h2d;
17'h398b:	data_out=16'hda;
17'h398c:	data_out=16'he3;
17'h398d:	data_out=16'h29;
17'h398e:	data_out=16'h8012;
17'h398f:	data_out=16'h2b;
17'h3990:	data_out=16'h80af;
17'h3991:	data_out=16'h82;
17'h3992:	data_out=16'h25;
17'h3993:	data_out=16'h16;
17'h3994:	data_out=16'hf8;
17'h3995:	data_out=16'h8040;
17'h3996:	data_out=16'h8027;
17'h3997:	data_out=16'h136;
17'h3998:	data_out=16'h8066;
17'h3999:	data_out=16'h1a;
17'h399a:	data_out=16'h83;
17'h399b:	data_out=16'h124;
17'h399c:	data_out=16'h139;
17'h399d:	data_out=16'hc5;
17'h399e:	data_out=16'hcc;
17'h399f:	data_out=16'h5a;
17'h39a0:	data_out=16'hf2;
17'h39a1:	data_out=16'h800f;
17'h39a2:	data_out=16'h8023;
17'h39a3:	data_out=16'h8145;
17'h39a4:	data_out=16'h8149;
17'h39a5:	data_out=16'h802d;
17'h39a6:	data_out=16'h8093;
17'h39a7:	data_out=16'h106;
17'h39a8:	data_out=16'h8008;
17'h39a9:	data_out=16'he;
17'h39aa:	data_out=16'h8046;
17'h39ab:	data_out=16'h67;
17'h39ac:	data_out=16'hc;
17'h39ad:	data_out=16'h8024;
17'h39ae:	data_out=16'hf;
17'h39af:	data_out=16'h96;
17'h39b0:	data_out=16'hc5;
17'h39b1:	data_out=16'h78;
17'h39b2:	data_out=16'hc3;
17'h39b3:	data_out=16'he4;
17'h39b4:	data_out=16'h801b;
17'h39b5:	data_out=16'hd0;
17'h39b6:	data_out=16'h32;
17'h39b7:	data_out=16'hab;
17'h39b8:	data_out=16'h36;
17'h39b9:	data_out=16'h7f;
17'h39ba:	data_out=16'h80d4;
17'h39bb:	data_out=16'h5d;
17'h39bc:	data_out=16'h10e;
17'h39bd:	data_out=16'h8036;
17'h39be:	data_out=16'h8008;
17'h39bf:	data_out=16'hc3;
17'h39c0:	data_out=16'h8021;
17'h39c1:	data_out=16'h111;
17'h39c2:	data_out=16'h8077;
17'h39c3:	data_out=16'h71;
17'h39c4:	data_out=16'h78;
17'h39c5:	data_out=16'h807b;
17'h39c6:	data_out=16'h117;
17'h39c7:	data_out=16'h809f;
17'h39c8:	data_out=16'h19;
17'h39c9:	data_out=16'h803f;
17'h39ca:	data_out=16'h2a;
17'h39cb:	data_out=16'h31;
17'h39cc:	data_out=16'h8064;
17'h39cd:	data_out=16'h800d;
17'h39ce:	data_out=16'h43;
17'h39cf:	data_out=16'h807d;
17'h39d0:	data_out=16'h12;
17'h39d1:	data_out=16'h5f;
17'h39d2:	data_out=16'h8155;
17'h39d3:	data_out=16'h20d;
17'h39d4:	data_out=16'h7b;
17'h39d5:	data_out=16'hdb;
17'h39d6:	data_out=16'h6;
17'h39d7:	data_out=16'h8065;
17'h39d8:	data_out=16'hce;
17'h39d9:	data_out=16'h8044;
17'h39da:	data_out=16'h178;
17'h39db:	data_out=16'hc6;
17'h39dc:	data_out=16'hf1;
17'h39dd:	data_out=16'h1a;
17'h39de:	data_out=16'haa;
17'h39df:	data_out=16'h801e;
17'h39e0:	data_out=16'h809b;
17'h39e1:	data_out=16'ha3;
17'h39e2:	data_out=16'hfe;
17'h39e3:	data_out=16'hf3;
17'h39e4:	data_out=16'h8019;
17'h39e5:	data_out=16'h20;
17'h39e6:	data_out=16'h33;
17'h39e7:	data_out=16'h29;
17'h39e8:	data_out=16'h800c;
17'h39e9:	data_out=16'h29;
17'h39ea:	data_out=16'h8009;
17'h39eb:	data_out=16'haa;
17'h39ec:	data_out=16'h8037;
17'h39ed:	data_out=16'hf6;
17'h39ee:	data_out=16'h8010;
17'h39ef:	data_out=16'h90;
17'h39f0:	data_out=16'h800d;
17'h39f1:	data_out=16'h8043;
17'h39f2:	data_out=16'h26;
17'h39f3:	data_out=16'h6c;
17'h39f4:	data_out=16'hc9;
17'h39f5:	data_out=16'h18a;
17'h39f6:	data_out=16'h8025;
17'h39f7:	data_out=16'h8028;
17'h39f8:	data_out=16'h59;
17'h39f9:	data_out=16'h8011;
17'h39fa:	data_out=16'hfb;
17'h39fb:	data_out=16'h8002;
17'h39fc:	data_out=16'h8027;
17'h39fd:	data_out=16'h31;
17'h39fe:	data_out=16'h807f;
17'h39ff:	data_out=16'h8050;
17'h3a00:	data_out=16'h86b3;
17'h3a01:	data_out=16'h85ae;
17'h3a02:	data_out=16'h82df;
17'h3a03:	data_out=16'h819f;
17'h3a04:	data_out=16'h2e;
17'h3a05:	data_out=16'h1a2;
17'h3a06:	data_out=16'h17e;
17'h3a07:	data_out=16'hac;
17'h3a08:	data_out=16'h8511;
17'h3a09:	data_out=16'h80f4;
17'h3a0a:	data_out=16'h8654;
17'h3a0b:	data_out=16'h294;
17'h3a0c:	data_out=16'h131;
17'h3a0d:	data_out=16'h30;
17'h3a0e:	data_out=16'h80b6;
17'h3a0f:	data_out=16'h8281;
17'h3a10:	data_out=16'h82e3;
17'h3a11:	data_out=16'h818c;
17'h3a12:	data_out=16'h5;
17'h3a13:	data_out=16'h805c;
17'h3a14:	data_out=16'h8136;
17'h3a15:	data_out=16'h828f;
17'h3a16:	data_out=16'h82ee;
17'h3a17:	data_out=16'h801e;
17'h3a18:	data_out=16'h8103;
17'h3a19:	data_out=16'h11c;
17'h3a1a:	data_out=16'h174;
17'h3a1b:	data_out=16'he8;
17'h3a1c:	data_out=16'h8217;
17'h3a1d:	data_out=16'h84f2;
17'h3a1e:	data_out=16'h80d1;
17'h3a1f:	data_out=16'h12b;
17'h3a20:	data_out=16'h81cd;
17'h3a21:	data_out=16'h80a4;
17'h3a22:	data_out=16'h90;
17'h3a23:	data_out=16'h83bb;
17'h3a24:	data_out=16'h83bb;
17'h3a25:	data_out=16'h36;
17'h3a26:	data_out=16'h83a7;
17'h3a27:	data_out=16'h83de;
17'h3a28:	data_out=16'h8085;
17'h3a29:	data_out=16'h82f5;
17'h3a2a:	data_out=16'h82b1;
17'h3a2b:	data_out=16'hc3;
17'h3a2c:	data_out=16'h8241;
17'h3a2d:	data_out=16'h84b0;
17'h3a2e:	data_out=16'h80d2;
17'h3a2f:	data_out=16'h8186;
17'h3a30:	data_out=16'h282;
17'h3a31:	data_out=16'h80e0;
17'h3a32:	data_out=16'h253;
17'h3a33:	data_out=16'h812c;
17'h3a34:	data_out=16'h839b;
17'h3a35:	data_out=16'h807b;
17'h3a36:	data_out=16'h851b;
17'h3a37:	data_out=16'h829b;
17'h3a38:	data_out=16'h838b;
17'h3a39:	data_out=16'h816f;
17'h3a3a:	data_out=16'h82e1;
17'h3a3b:	data_out=16'h8113;
17'h3a3c:	data_out=16'h840f;
17'h3a3d:	data_out=16'h8418;
17'h3a3e:	data_out=16'h8086;
17'h3a3f:	data_out=16'h122;
17'h3a40:	data_out=16'h104;
17'h3a41:	data_out=16'h80be;
17'h3a42:	data_out=16'h80d2;
17'h3a43:	data_out=16'h222;
17'h3a44:	data_out=16'h8272;
17'h3a45:	data_out=16'h8297;
17'h3a46:	data_out=16'h8173;
17'h3a47:	data_out=16'h8134;
17'h3a48:	data_out=16'h23c;
17'h3a49:	data_out=16'h12;
17'h3a4a:	data_out=16'h20e;
17'h3a4b:	data_out=16'hfb;
17'h3a4c:	data_out=16'hdf;
17'h3a4d:	data_out=16'h52;
17'h3a4e:	data_out=16'h8236;
17'h3a4f:	data_out=16'h73;
17'h3a50:	data_out=16'hb6;
17'h3a51:	data_out=16'h81c5;
17'h3a52:	data_out=16'h845e;
17'h3a53:	data_out=16'hf1;
17'h3a54:	data_out=16'h83ce;
17'h3a55:	data_out=16'h82dc;
17'h3a56:	data_out=16'h83a9;
17'h3a57:	data_out=16'h83d4;
17'h3a58:	data_out=16'h83f6;
17'h3a59:	data_out=16'h822c;
17'h3a5a:	data_out=16'h260;
17'h3a5b:	data_out=16'h83c1;
17'h3a5c:	data_out=16'h8161;
17'h3a5d:	data_out=16'h829b;
17'h3a5e:	data_out=16'h80cb;
17'h3a5f:	data_out=16'h815e;
17'h3a60:	data_out=16'h852a;
17'h3a61:	data_out=16'h82c5;
17'h3a62:	data_out=16'h145;
17'h3a63:	data_out=16'h8117;
17'h3a64:	data_out=16'h8274;
17'h3a65:	data_out=16'hef;
17'h3a66:	data_out=16'h12b;
17'h3a67:	data_out=16'h68;
17'h3a68:	data_out=16'h809f;
17'h3a69:	data_out=16'h85c4;
17'h3a6a:	data_out=16'h80d1;
17'h3a6b:	data_out=16'h9c;
17'h3a6c:	data_out=16'h88b0;
17'h3a6d:	data_out=16'h80f3;
17'h3a6e:	data_out=16'h80d3;
17'h3a6f:	data_out=16'h263;
17'h3a70:	data_out=16'h80ca;
17'h3a71:	data_out=16'h8008;
17'h3a72:	data_out=16'h8197;
17'h3a73:	data_out=16'h815f;
17'h3a74:	data_out=16'h291;
17'h3a75:	data_out=16'h804c;
17'h3a76:	data_out=16'h8006;
17'h3a77:	data_out=16'h8153;
17'h3a78:	data_out=16'h25d;
17'h3a79:	data_out=16'h81cc;
17'h3a7a:	data_out=16'h8114;
17'h3a7b:	data_out=16'h807a;
17'h3a7c:	data_out=16'h80d0;
17'h3a7d:	data_out=16'h2ce;
17'h3a7e:	data_out=16'h80e3;
17'h3a7f:	data_out=16'h80a5;
17'h3a80:	data_out=16'h8a00;
17'h3a81:	data_out=16'h8a00;
17'h3a82:	data_out=16'h89ff;
17'h3a83:	data_out=16'h81bf;
17'h3a84:	data_out=16'h77d;
17'h3a85:	data_out=16'h9ff;
17'h3a86:	data_out=16'h9b5;
17'h3a87:	data_out=16'h83d1;
17'h3a88:	data_out=16'h89fe;
17'h3a89:	data_out=16'h89fc;
17'h3a8a:	data_out=16'h8a00;
17'h3a8b:	data_out=16'h77f;
17'h3a8c:	data_out=16'h582;
17'h3a8d:	data_out=16'h337;
17'h3a8e:	data_out=16'h835e;
17'h3a8f:	data_out=16'h8a00;
17'h3a90:	data_out=16'h89ff;
17'h3a91:	data_out=16'h1b6;
17'h3a92:	data_out=16'h88f4;
17'h3a93:	data_out=16'h93;
17'h3a94:	data_out=16'h8025;
17'h3a95:	data_out=16'h8688;
17'h3a96:	data_out=16'h88e9;
17'h3a97:	data_out=16'h24b;
17'h3a98:	data_out=16'h86a4;
17'h3a99:	data_out=16'ha00;
17'h3a9a:	data_out=16'ha00;
17'h3a9b:	data_out=16'h9a3;
17'h3a9c:	data_out=16'h6d;
17'h3a9d:	data_out=16'h8a00;
17'h3a9e:	data_out=16'h8477;
17'h3a9f:	data_out=16'h80e7;
17'h3aa0:	data_out=16'h21d;
17'h3aa1:	data_out=16'h830a;
17'h3aa2:	data_out=16'h862a;
17'h3aa3:	data_out=16'h8a00;
17'h3aa4:	data_out=16'h8a00;
17'h3aa5:	data_out=16'h868c;
17'h3aa6:	data_out=16'h8a00;
17'h3aa7:	data_out=16'h860a;
17'h3aa8:	data_out=16'h8292;
17'h3aa9:	data_out=16'h8783;
17'h3aaa:	data_out=16'h8a00;
17'h3aab:	data_out=16'h9fe;
17'h3aac:	data_out=16'h8788;
17'h3aad:	data_out=16'h8a00;
17'h3aae:	data_out=16'h89f9;
17'h3aaf:	data_out=16'h43;
17'h3ab0:	data_out=16'h979;
17'h3ab1:	data_out=16'h1e8;
17'h3ab2:	data_out=16'h91c;
17'h3ab3:	data_out=16'h822d;
17'h3ab4:	data_out=16'h897a;
17'h3ab5:	data_out=16'h636;
17'h3ab6:	data_out=16'h8a00;
17'h3ab7:	data_out=16'h89fe;
17'h3ab8:	data_out=16'h8078;
17'h3ab9:	data_out=16'h829e;
17'h3aba:	data_out=16'h8a00;
17'h3abb:	data_out=16'h8390;
17'h3abc:	data_out=16'h89ff;
17'h3abd:	data_out=16'h8a00;
17'h3abe:	data_out=16'h8290;
17'h3abf:	data_out=16'h9ff;
17'h3ac0:	data_out=16'h820b;
17'h3ac1:	data_out=16'h854e;
17'h3ac2:	data_out=16'h89fe;
17'h3ac3:	data_out=16'ha00;
17'h3ac4:	data_out=16'h8399;
17'h3ac5:	data_out=16'h86bc;
17'h3ac6:	data_out=16'h883b;
17'h3ac7:	data_out=16'h8a00;
17'h3ac8:	data_out=16'h8053;
17'h3ac9:	data_out=16'h8610;
17'h3aca:	data_out=16'h149;
17'h3acb:	data_out=16'h8376;
17'h3acc:	data_out=16'h8907;
17'h3acd:	data_out=16'h85b8;
17'h3ace:	data_out=16'h893b;
17'h3acf:	data_out=16'h89ff;
17'h3ad0:	data_out=16'h8249;
17'h3ad1:	data_out=16'h81df;
17'h3ad2:	data_out=16'h89ff;
17'h3ad3:	data_out=16'ha00;
17'h3ad4:	data_out=16'h88a9;
17'h3ad5:	data_out=16'h88a3;
17'h3ad6:	data_out=16'h8a00;
17'h3ad7:	data_out=16'h8a00;
17'h3ad8:	data_out=16'h89f3;
17'h3ad9:	data_out=16'h89e2;
17'h3ada:	data_out=16'h9ff;
17'h3adb:	data_out=16'h82f1;
17'h3adc:	data_out=16'h853;
17'h3add:	data_out=16'h8a00;
17'h3ade:	data_out=16'h800b;
17'h3adf:	data_out=16'h859f;
17'h3ae0:	data_out=16'h8a00;
17'h3ae1:	data_out=16'h8264;
17'h3ae2:	data_out=16'h99c;
17'h3ae3:	data_out=16'h8103;
17'h3ae4:	data_out=16'h846f;
17'h3ae5:	data_out=16'h55c;
17'h3ae6:	data_out=16'ha00;
17'h3ae7:	data_out=16'h877b;
17'h3ae8:	data_out=16'h82cd;
17'h3ae9:	data_out=16'h8a00;
17'h3aea:	data_out=16'h83ae;
17'h3aeb:	data_out=16'h86a;
17'h3aec:	data_out=16'h8a00;
17'h3aed:	data_out=16'h8183;
17'h3aee:	data_out=16'h83ac;
17'h3aef:	data_out=16'ha00;
17'h3af0:	data_out=16'h837d;
17'h3af1:	data_out=16'h89fe;
17'h3af2:	data_out=16'h822c;
17'h3af3:	data_out=16'h29b;
17'h3af4:	data_out=16'h9ac;
17'h3af5:	data_out=16'ha00;
17'h3af6:	data_out=16'h41f;
17'h3af7:	data_out=16'h890c;
17'h3af8:	data_out=16'ha00;
17'h3af9:	data_out=16'h8a00;
17'h3afa:	data_out=16'h802b;
17'h3afb:	data_out=16'h8290;
17'h3afc:	data_out=16'h8414;
17'h3afd:	data_out=16'ha00;
17'h3afe:	data_out=16'h8a00;
17'h3aff:	data_out=16'h8729;
17'h3b00:	data_out=16'h8a00;
17'h3b01:	data_out=16'h8a00;
17'h3b02:	data_out=16'h89ff;
17'h3b03:	data_out=16'h4b;
17'h3b04:	data_out=16'h9ff;
17'h3b05:	data_out=16'ha00;
17'h3b06:	data_out=16'ha00;
17'h3b07:	data_out=16'h57b;
17'h3b08:	data_out=16'h89fe;
17'h3b09:	data_out=16'h8035;
17'h3b0a:	data_out=16'h8a00;
17'h3b0b:	data_out=16'h8e5;
17'h3b0c:	data_out=16'ha00;
17'h3b0d:	data_out=16'h84cf;
17'h3b0e:	data_out=16'h8257;
17'h3b0f:	data_out=16'h89fe;
17'h3b10:	data_out=16'h8280;
17'h3b11:	data_out=16'h79b;
17'h3b12:	data_out=16'h82c2;
17'h3b13:	data_out=16'h810a;
17'h3b14:	data_out=16'h8055;
17'h3b15:	data_out=16'h8354;
17'h3b16:	data_out=16'h884b;
17'h3b17:	data_out=16'h8126;
17'h3b18:	data_out=16'h8608;
17'h3b19:	data_out=16'ha00;
17'h3b1a:	data_out=16'ha00;
17'h3b1b:	data_out=16'h899;
17'h3b1c:	data_out=16'h355;
17'h3b1d:	data_out=16'h853b;
17'h3b1e:	data_out=16'h8404;
17'h3b1f:	data_out=16'h6bc;
17'h3b20:	data_out=16'h9c6;
17'h3b21:	data_out=16'h81b4;
17'h3b22:	data_out=16'h824;
17'h3b23:	data_out=16'h8a00;
17'h3b24:	data_out=16'h8a00;
17'h3b25:	data_out=16'h219;
17'h3b26:	data_out=16'h8a00;
17'h3b27:	data_out=16'h63;
17'h3b28:	data_out=16'h807d;
17'h3b29:	data_out=16'h86b0;
17'h3b2a:	data_out=16'h89ff;
17'h3b2b:	data_out=16'ha00;
17'h3b2c:	data_out=16'h863d;
17'h3b2d:	data_out=16'h8a00;
17'h3b2e:	data_out=16'h890f;
17'h3b2f:	data_out=16'h869;
17'h3b30:	data_out=16'ha00;
17'h3b31:	data_out=16'h318;
17'h3b32:	data_out=16'ha00;
17'h3b33:	data_out=16'h800a;
17'h3b34:	data_out=16'h8507;
17'h3b35:	data_out=16'h873;
17'h3b36:	data_out=16'h89ff;
17'h3b37:	data_out=16'h89fd;
17'h3b38:	data_out=16'h9ff;
17'h3b39:	data_out=16'h806d;
17'h3b3a:	data_out=16'h82a4;
17'h3b3b:	data_out=16'hd0;
17'h3b3c:	data_out=16'h89fd;
17'h3b3d:	data_out=16'h466;
17'h3b3e:	data_out=16'h8062;
17'h3b3f:	data_out=16'ha00;
17'h3b40:	data_out=16'ha00;
17'h3b41:	data_out=16'h89ff;
17'h3b42:	data_out=16'h89fe;
17'h3b43:	data_out=16'ha00;
17'h3b44:	data_out=16'hb2;
17'h3b45:	data_out=16'h82f3;
17'h3b46:	data_out=16'h88f9;
17'h3b47:	data_out=16'h831a;
17'h3b48:	data_out=16'h703;
17'h3b49:	data_out=16'h370;
17'h3b4a:	data_out=16'h841;
17'h3b4b:	data_out=16'h89fb;
17'h3b4c:	data_out=16'h8833;
17'h3b4d:	data_out=16'h92e;
17'h3b4e:	data_out=16'h8859;
17'h3b4f:	data_out=16'h858a;
17'h3b50:	data_out=16'h9ff;
17'h3b51:	data_out=16'h8661;
17'h3b52:	data_out=16'h89f2;
17'h3b53:	data_out=16'ha00;
17'h3b54:	data_out=16'h271;
17'h3b55:	data_out=16'h89dc;
17'h3b56:	data_out=16'h89d1;
17'h3b57:	data_out=16'h874e;
17'h3b58:	data_out=16'h89fd;
17'h3b59:	data_out=16'h30a;
17'h3b5a:	data_out=16'h438;
17'h3b5b:	data_out=16'h806a;
17'h3b5c:	data_out=16'h9ba;
17'h3b5d:	data_out=16'h8a00;
17'h3b5e:	data_out=16'h7ff;
17'h3b5f:	data_out=16'h83c8;
17'h3b60:	data_out=16'h8a00;
17'h3b61:	data_out=16'h82;
17'h3b62:	data_out=16'h23d;
17'h3b63:	data_out=16'hb5;
17'h3b64:	data_out=16'h140;
17'h3b65:	data_out=16'ha00;
17'h3b66:	data_out=16'ha00;
17'h3b67:	data_out=16'h1cc;
17'h3b68:	data_out=16'h8134;
17'h3b69:	data_out=16'h8a00;
17'h3b6a:	data_out=16'h831e;
17'h3b6b:	data_out=16'h9f9;
17'h3b6c:	data_out=16'h8a00;
17'h3b6d:	data_out=16'h78;
17'h3b6e:	data_out=16'h831d;
17'h3b6f:	data_out=16'ha00;
17'h3b70:	data_out=16'h827d;
17'h3b71:	data_out=16'h89fd;
17'h3b72:	data_out=16'h207;
17'h3b73:	data_out=16'h6fe;
17'h3b74:	data_out=16'ha00;
17'h3b75:	data_out=16'h495;
17'h3b76:	data_out=16'ha00;
17'h3b77:	data_out=16'h3c6;
17'h3b78:	data_out=16'ha00;
17'h3b79:	data_out=16'h8a00;
17'h3b7a:	data_out=16'h63;
17'h3b7b:	data_out=16'h8049;
17'h3b7c:	data_out=16'h8347;
17'h3b7d:	data_out=16'ha00;
17'h3b7e:	data_out=16'ha4;
17'h3b7f:	data_out=16'h46f;
17'h3b80:	data_out=16'h8a00;
17'h3b81:	data_out=16'h8a00;
17'h3b82:	data_out=16'h8a00;
17'h3b83:	data_out=16'h89fe;
17'h3b84:	data_out=16'h9fa;
17'h3b85:	data_out=16'h9ca;
17'h3b86:	data_out=16'h89e;
17'h3b87:	data_out=16'ha00;
17'h3b88:	data_out=16'h8a00;
17'h3b89:	data_out=16'h1a3;
17'h3b8a:	data_out=16'h88ae;
17'h3b8b:	data_out=16'h643;
17'h3b8c:	data_out=16'ha00;
17'h3b8d:	data_out=16'h89ff;
17'h3b8e:	data_out=16'h197;
17'h3b8f:	data_out=16'h89fd;
17'h3b90:	data_out=16'h8378;
17'h3b91:	data_out=16'h6aa;
17'h3b92:	data_out=16'h88aa;
17'h3b93:	data_out=16'h89fc;
17'h3b94:	data_out=16'h8761;
17'h3b95:	data_out=16'h86f9;
17'h3b96:	data_out=16'h8a00;
17'h3b97:	data_out=16'h89f0;
17'h3b98:	data_out=16'h8a00;
17'h3b99:	data_out=16'ha00;
17'h3b9a:	data_out=16'ha00;
17'h3b9b:	data_out=16'h26b;
17'h3b9c:	data_out=16'ha8;
17'h3b9d:	data_out=16'h83b1;
17'h3b9e:	data_out=16'h89ff;
17'h3b9f:	data_out=16'h701;
17'h3ba0:	data_out=16'h908;
17'h3ba1:	data_out=16'h1eb;
17'h3ba2:	data_out=16'h9f3;
17'h3ba3:	data_out=16'h89e5;
17'h3ba4:	data_out=16'h89df;
17'h3ba5:	data_out=16'h1d5;
17'h3ba6:	data_out=16'h8a00;
17'h3ba7:	data_out=16'h54;
17'h3ba8:	data_out=16'h24b;
17'h3ba9:	data_out=16'h875a;
17'h3baa:	data_out=16'h8a00;
17'h3bab:	data_out=16'ha00;
17'h3bac:	data_out=16'h8a00;
17'h3bad:	data_out=16'h8754;
17'h3bae:	data_out=16'h8841;
17'h3baf:	data_out=16'h7fa;
17'h3bb0:	data_out=16'ha00;
17'h3bb1:	data_out=16'h659;
17'h3bb2:	data_out=16'ha00;
17'h3bb3:	data_out=16'h8606;
17'h3bb4:	data_out=16'h41;
17'h3bb5:	data_out=16'h67e;
17'h3bb6:	data_out=16'h8a00;
17'h3bb7:	data_out=16'h89ff;
17'h3bb8:	data_out=16'h9ff;
17'h3bb9:	data_out=16'h86b2;
17'h3bba:	data_out=16'h81a3;
17'h3bbb:	data_out=16'h4f7;
17'h3bbc:	data_out=16'h89fa;
17'h3bbd:	data_out=16'h313;
17'h3bbe:	data_out=16'h24c;
17'h3bbf:	data_out=16'h9c7;
17'h3bc0:	data_out=16'h9ff;
17'h3bc1:	data_out=16'h8a00;
17'h3bc2:	data_out=16'h89f9;
17'h3bc3:	data_out=16'h9e3;
17'h3bc4:	data_out=16'h82ec;
17'h3bc5:	data_out=16'h86c3;
17'h3bc6:	data_out=16'h87e5;
17'h3bc7:	data_out=16'h84f3;
17'h3bc8:	data_out=16'h9f6;
17'h3bc9:	data_out=16'h4bc;
17'h3bca:	data_out=16'ha00;
17'h3bcb:	data_out=16'h89fa;
17'h3bcc:	data_out=16'h8a00;
17'h3bcd:	data_out=16'h9f5;
17'h3bce:	data_out=16'h868c;
17'h3bcf:	data_out=16'h8995;
17'h3bd0:	data_out=16'h9f3;
17'h3bd1:	data_out=16'h89ff;
17'h3bd2:	data_out=16'h884d;
17'h3bd3:	data_out=16'ha00;
17'h3bd4:	data_out=16'h1c9;
17'h3bd5:	data_out=16'h89fa;
17'h3bd6:	data_out=16'h8a00;
17'h3bd7:	data_out=16'h8a00;
17'h3bd8:	data_out=16'h89fe;
17'h3bd9:	data_out=16'h4b6;
17'h3bda:	data_out=16'h8343;
17'h3bdb:	data_out=16'h41a;
17'h3bdc:	data_out=16'h7c3;
17'h3bdd:	data_out=16'h8a00;
17'h3bde:	data_out=16'h7b0;
17'h3bdf:	data_out=16'h8600;
17'h3be0:	data_out=16'h8a00;
17'h3be1:	data_out=16'h8185;
17'h3be2:	data_out=16'h89c5;
17'h3be3:	data_out=16'h84f2;
17'h3be4:	data_out=16'h446;
17'h3be5:	data_out=16'ha00;
17'h3be6:	data_out=16'ha00;
17'h3be7:	data_out=16'h59c;
17'h3be8:	data_out=16'h21a;
17'h3be9:	data_out=16'h8a00;
17'h3bea:	data_out=16'h157;
17'h3beb:	data_out=16'h99e;
17'h3bec:	data_out=16'h8a00;
17'h3bed:	data_out=16'h852d;
17'h3bee:	data_out=16'h157;
17'h3bef:	data_out=16'ha00;
17'h3bf0:	data_out=16'h17e;
17'h3bf1:	data_out=16'h89fc;
17'h3bf2:	data_out=16'h179;
17'h3bf3:	data_out=16'h570;
17'h3bf4:	data_out=16'ha00;
17'h3bf5:	data_out=16'h118;
17'h3bf6:	data_out=16'ha00;
17'h3bf7:	data_out=16'h3ab;
17'h3bf8:	data_out=16'ha00;
17'h3bf9:	data_out=16'h8971;
17'h3bfa:	data_out=16'h8614;
17'h3bfb:	data_out=16'h24a;
17'h3bfc:	data_out=16'h8544;
17'h3bfd:	data_out=16'ha00;
17'h3bfe:	data_out=16'h81c0;
17'h3bff:	data_out=16'h5ce;
17'h3c00:	data_out=16'h8a00;
17'h3c01:	data_out=16'h8a00;
17'h3c02:	data_out=16'h8a00;
17'h3c03:	data_out=16'h89fc;
17'h3c04:	data_out=16'ha00;
17'h3c05:	data_out=16'h9f3;
17'h3c06:	data_out=16'h244;
17'h3c07:	data_out=16'ha00;
17'h3c08:	data_out=16'h8a00;
17'h3c09:	data_out=16'h86b2;
17'h3c0a:	data_out=16'ha2;
17'h3c0b:	data_out=16'h87ab;
17'h3c0c:	data_out=16'ha00;
17'h3c0d:	data_out=16'h89fe;
17'h3c0e:	data_out=16'h8033;
17'h3c0f:	data_out=16'h89ff;
17'h3c10:	data_out=16'h8553;
17'h3c11:	data_out=16'h573;
17'h3c12:	data_out=16'h8a00;
17'h3c13:	data_out=16'h89f8;
17'h3c14:	data_out=16'h89f3;
17'h3c15:	data_out=16'h89ff;
17'h3c16:	data_out=16'h89f9;
17'h3c17:	data_out=16'h89ea;
17'h3c18:	data_out=16'h8a00;
17'h3c19:	data_out=16'ha00;
17'h3c1a:	data_out=16'ha00;
17'h3c1b:	data_out=16'h8414;
17'h3c1c:	data_out=16'h285;
17'h3c1d:	data_out=16'h8879;
17'h3c1e:	data_out=16'h89fa;
17'h3c1f:	data_out=16'h8360;
17'h3c20:	data_out=16'h82a;
17'h3c21:	data_out=16'h38;
17'h3c22:	data_out=16'h998;
17'h3c23:	data_out=16'h89f8;
17'h3c24:	data_out=16'h89f8;
17'h3c25:	data_out=16'h8927;
17'h3c26:	data_out=16'h8a00;
17'h3c27:	data_out=16'h87fd;
17'h3c28:	data_out=16'hd7;
17'h3c29:	data_out=16'h880c;
17'h3c2a:	data_out=16'h8a00;
17'h3c2b:	data_out=16'ha00;
17'h3c2c:	data_out=16'h89f9;
17'h3c2d:	data_out=16'h8653;
17'h3c2e:	data_out=16'h88ed;
17'h3c2f:	data_out=16'h5d6;
17'h3c30:	data_out=16'h9ff;
17'h3c31:	data_out=16'h826;
17'h3c32:	data_out=16'ha00;
17'h3c33:	data_out=16'h89ef;
17'h3c34:	data_out=16'h46e;
17'h3c35:	data_out=16'h425;
17'h3c36:	data_out=16'h8a00;
17'h3c37:	data_out=16'h89ff;
17'h3c38:	data_out=16'h9ff;
17'h3c39:	data_out=16'h89f2;
17'h3c3a:	data_out=16'h884c;
17'h3c3b:	data_out=16'h9fd;
17'h3c3c:	data_out=16'h89f1;
17'h3c3d:	data_out=16'h8960;
17'h3c3e:	data_out=16'hd9;
17'h3c3f:	data_out=16'h9f2;
17'h3c40:	data_out=16'ha00;
17'h3c41:	data_out=16'h8a00;
17'h3c42:	data_out=16'h89e7;
17'h3c43:	data_out=16'h8ef;
17'h3c44:	data_out=16'h86cf;
17'h3c45:	data_out=16'h89ff;
17'h3c46:	data_out=16'h876a;
17'h3c47:	data_out=16'h89fe;
17'h3c48:	data_out=16'h1de;
17'h3c49:	data_out=16'h8828;
17'h3c4a:	data_out=16'ha00;
17'h3c4b:	data_out=16'h89fc;
17'h3c4c:	data_out=16'h8a00;
17'h3c4d:	data_out=16'h9f4;
17'h3c4e:	data_out=16'h83d5;
17'h3c4f:	data_out=16'h8a00;
17'h3c50:	data_out=16'h9eb;
17'h3c51:	data_out=16'h89ff;
17'h3c52:	data_out=16'h88d9;
17'h3c53:	data_out=16'ha00;
17'h3c54:	data_out=16'h8572;
17'h3c55:	data_out=16'h89fc;
17'h3c56:	data_out=16'h8a00;
17'h3c57:	data_out=16'h89fb;
17'h3c58:	data_out=16'h89ff;
17'h3c59:	data_out=16'h251;
17'h3c5a:	data_out=16'h856d;
17'h3c5b:	data_out=16'h9af;
17'h3c5c:	data_out=16'h9d2;
17'h3c5d:	data_out=16'h89fc;
17'h3c5e:	data_out=16'h5bf;
17'h3c5f:	data_out=16'h89fe;
17'h3c60:	data_out=16'h8a00;
17'h3c61:	data_out=16'h366;
17'h3c62:	data_out=16'h89f9;
17'h3c63:	data_out=16'h8946;
17'h3c64:	data_out=16'h8332;
17'h3c65:	data_out=16'h9fe;
17'h3c66:	data_out=16'ha00;
17'h3c67:	data_out=16'h38c;
17'h3c68:	data_out=16'h7c;
17'h3c69:	data_out=16'h8a00;
17'h3c6a:	data_out=16'h806c;
17'h3c6b:	data_out=16'h990;
17'h3c6c:	data_out=16'h89fe;
17'h3c6d:	data_out=16'h8976;
17'h3c6e:	data_out=16'h806c;
17'h3c6f:	data_out=16'ha00;
17'h3c70:	data_out=16'h8050;
17'h3c71:	data_out=16'h89fd;
17'h3c72:	data_out=16'h86f;
17'h3c73:	data_out=16'h9fb;
17'h3c74:	data_out=16'h9fe;
17'h3c75:	data_out=16'h134;
17'h3c76:	data_out=16'ha00;
17'h3c77:	data_out=16'h89fd;
17'h3c78:	data_out=16'ha00;
17'h3c79:	data_out=16'h8828;
17'h3c7a:	data_out=16'h89f1;
17'h3c7b:	data_out=16'hd5;
17'h3c7c:	data_out=16'h89ff;
17'h3c7d:	data_out=16'ha00;
17'h3c7e:	data_out=16'h8a00;
17'h3c7f:	data_out=16'h8435;
17'h3c80:	data_out=16'h89eb;
17'h3c81:	data_out=16'h6b6;
17'h3c82:	data_out=16'h8a00;
17'h3c83:	data_out=16'h89fe;
17'h3c84:	data_out=16'ha00;
17'h3c85:	data_out=16'h9ff;
17'h3c86:	data_out=16'h89fd;
17'h3c87:	data_out=16'h741;
17'h3c88:	data_out=16'h89f7;
17'h3c89:	data_out=16'h89ff;
17'h3c8a:	data_out=16'ha00;
17'h3c8b:	data_out=16'h8926;
17'h3c8c:	data_out=16'h83e;
17'h3c8d:	data_out=16'h8a00;
17'h3c8e:	data_out=16'h831a;
17'h3c8f:	data_out=16'h8a00;
17'h3c90:	data_out=16'h806b;
17'h3c91:	data_out=16'h7a6;
17'h3c92:	data_out=16'h8a00;
17'h3c93:	data_out=16'h89fb;
17'h3c94:	data_out=16'h89f1;
17'h3c95:	data_out=16'h88d1;
17'h3c96:	data_out=16'h89f6;
17'h3c97:	data_out=16'h89f1;
17'h3c98:	data_out=16'h89fe;
17'h3c99:	data_out=16'ha00;
17'h3c9a:	data_out=16'ha00;
17'h3c9b:	data_out=16'h89fb;
17'h3c9c:	data_out=16'h680;
17'h3c9d:	data_out=16'h790;
17'h3c9e:	data_out=16'h89f9;
17'h3c9f:	data_out=16'h84a0;
17'h3ca0:	data_out=16'h99c;
17'h3ca1:	data_out=16'h82c2;
17'h3ca2:	data_out=16'h29b;
17'h3ca3:	data_out=16'h87df;
17'h3ca4:	data_out=16'h87dc;
17'h3ca5:	data_out=16'h89e9;
17'h3ca6:	data_out=16'h8a00;
17'h3ca7:	data_out=16'h958;
17'h3ca8:	data_out=16'h8228;
17'h3ca9:	data_out=16'h876c;
17'h3caa:	data_out=16'h8a00;
17'h3cab:	data_out=16'ha00;
17'h3cac:	data_out=16'h89ef;
17'h3cad:	data_out=16'h8922;
17'h3cae:	data_out=16'h89d2;
17'h3caf:	data_out=16'h99d;
17'h3cb0:	data_out=16'ha00;
17'h3cb1:	data_out=16'h9f5;
17'h3cb2:	data_out=16'ha00;
17'h3cb3:	data_out=16'h8968;
17'h3cb4:	data_out=16'h9fe;
17'h3cb5:	data_out=16'h888;
17'h3cb6:	data_out=16'h89f8;
17'h3cb7:	data_out=16'h89fe;
17'h3cb8:	data_out=16'ha00;
17'h3cb9:	data_out=16'h89ec;
17'h3cba:	data_out=16'h87bb;
17'h3cbb:	data_out=16'ha00;
17'h3cbc:	data_out=16'h89f9;
17'h3cbd:	data_out=16'h89d;
17'h3cbe:	data_out=16'h8228;
17'h3cbf:	data_out=16'h9ff;
17'h3cc0:	data_out=16'ha00;
17'h3cc1:	data_out=16'h8a00;
17'h3cc2:	data_out=16'h89f2;
17'h3cc3:	data_out=16'h675;
17'h3cc4:	data_out=16'h835;
17'h3cc5:	data_out=16'h89a6;
17'h3cc6:	data_out=16'h8a00;
17'h3cc7:	data_out=16'h89fd;
17'h3cc8:	data_out=16'h887b;
17'h3cc9:	data_out=16'h871b;
17'h3cca:	data_out=16'h442;
17'h3ccb:	data_out=16'h8a00;
17'h3ccc:	data_out=16'h8a00;
17'h3ccd:	data_out=16'h997;
17'h3cce:	data_out=16'h817e;
17'h3ccf:	data_out=16'h8a00;
17'h3cd0:	data_out=16'h9f6;
17'h3cd1:	data_out=16'h8a00;
17'h3cd2:	data_out=16'h83cd;
17'h3cd3:	data_out=16'ha00;
17'h3cd4:	data_out=16'h991;
17'h3cd5:	data_out=16'h89fd;
17'h3cd6:	data_out=16'h8a00;
17'h3cd7:	data_out=16'h8980;
17'h3cd8:	data_out=16'h89fc;
17'h3cd9:	data_out=16'h9f6;
17'h3cda:	data_out=16'h89f4;
17'h3cdb:	data_out=16'ha00;
17'h3cdc:	data_out=16'h9d1;
17'h3cdd:	data_out=16'h88f2;
17'h3cde:	data_out=16'h756;
17'h3cdf:	data_out=16'h89b5;
17'h3ce0:	data_out=16'h89ff;
17'h3ce1:	data_out=16'ha00;
17'h3ce2:	data_out=16'h89f8;
17'h3ce3:	data_out=16'h886c;
17'h3ce4:	data_out=16'h31;
17'h3ce5:	data_out=16'ha00;
17'h3ce6:	data_out=16'ha00;
17'h3ce7:	data_out=16'h958;
17'h3ce8:	data_out=16'h8285;
17'h3ce9:	data_out=16'h8a00;
17'h3cea:	data_out=16'h8349;
17'h3ceb:	data_out=16'h9db;
17'h3cec:	data_out=16'h89e8;
17'h3ced:	data_out=16'h8892;
17'h3cee:	data_out=16'h8349;
17'h3cef:	data_out=16'ha00;
17'h3cf0:	data_out=16'h8332;
17'h3cf1:	data_out=16'h89fe;
17'h3cf2:	data_out=16'h8f9;
17'h3cf3:	data_out=16'h9fd;
17'h3cf4:	data_out=16'h9fd;
17'h3cf5:	data_out=16'h804f;
17'h3cf6:	data_out=16'ha00;
17'h3cf7:	data_out=16'h8a00;
17'h3cf8:	data_out=16'ha00;
17'h3cf9:	data_out=16'h86e8;
17'h3cfa:	data_out=16'h89ee;
17'h3cfb:	data_out=16'h822c;
17'h3cfc:	data_out=16'h89fc;
17'h3cfd:	data_out=16'ha00;
17'h3cfe:	data_out=16'h8a00;
17'h3cff:	data_out=16'h8003;
17'h3d00:	data_out=16'h89f5;
17'h3d01:	data_out=16'h9ef;
17'h3d02:	data_out=16'h89f6;
17'h3d03:	data_out=16'h8a00;
17'h3d04:	data_out=16'ha00;
17'h3d05:	data_out=16'ha00;
17'h3d06:	data_out=16'h89fa;
17'h3d07:	data_out=16'h54b;
17'h3d08:	data_out=16'h89e1;
17'h3d09:	data_out=16'h8a00;
17'h3d0a:	data_out=16'ha00;
17'h3d0b:	data_out=16'h89f4;
17'h3d0c:	data_out=16'h9fe;
17'h3d0d:	data_out=16'h8a00;
17'h3d0e:	data_out=16'h828c;
17'h3d0f:	data_out=16'h8a00;
17'h3d10:	data_out=16'h873e;
17'h3d11:	data_out=16'h598;
17'h3d12:	data_out=16'h8a00;
17'h3d13:	data_out=16'h8a00;
17'h3d14:	data_out=16'h89ec;
17'h3d15:	data_out=16'h85f1;
17'h3d16:	data_out=16'h89e1;
17'h3d17:	data_out=16'h89e8;
17'h3d18:	data_out=16'h89ff;
17'h3d19:	data_out=16'ha00;
17'h3d1a:	data_out=16'ha00;
17'h3d1b:	data_out=16'h89e6;
17'h3d1c:	data_out=16'h6f2;
17'h3d1d:	data_out=16'h5ca;
17'h3d1e:	data_out=16'h89fa;
17'h3d1f:	data_out=16'h87d6;
17'h3d20:	data_out=16'h9c2;
17'h3d21:	data_out=16'h8223;
17'h3d22:	data_out=16'h89fe;
17'h3d23:	data_out=16'h8714;
17'h3d24:	data_out=16'h8710;
17'h3d25:	data_out=16'h89fb;
17'h3d26:	data_out=16'h89ff;
17'h3d27:	data_out=16'h73c;
17'h3d28:	data_out=16'h8156;
17'h3d29:	data_out=16'h887e;
17'h3d2a:	data_out=16'h89ff;
17'h3d2b:	data_out=16'ha00;
17'h3d2c:	data_out=16'h89e0;
17'h3d2d:	data_out=16'h89ff;
17'h3d2e:	data_out=16'h89d9;
17'h3d2f:	data_out=16'h8015;
17'h3d30:	data_out=16'ha00;
17'h3d31:	data_out=16'h9ef;
17'h3d32:	data_out=16'ha00;
17'h3d33:	data_out=16'h89f0;
17'h3d34:	data_out=16'h9f5;
17'h3d35:	data_out=16'h88b;
17'h3d36:	data_out=16'h89dc;
17'h3d37:	data_out=16'h89e4;
17'h3d38:	data_out=16'h9e5;
17'h3d39:	data_out=16'h89f7;
17'h3d3a:	data_out=16'h89ff;
17'h3d3b:	data_out=16'ha00;
17'h3d3c:	data_out=16'h8970;
17'h3d3d:	data_out=16'h152;
17'h3d3e:	data_out=16'h8155;
17'h3d3f:	data_out=16'ha00;
17'h3d40:	data_out=16'ha00;
17'h3d41:	data_out=16'h89f1;
17'h3d42:	data_out=16'h89ff;
17'h3d43:	data_out=16'h50a;
17'h3d44:	data_out=16'h7d2;
17'h3d45:	data_out=16'h8754;
17'h3d46:	data_out=16'h89fe;
17'h3d47:	data_out=16'h8a00;
17'h3d48:	data_out=16'h8a00;
17'h3d49:	data_out=16'h89f7;
17'h3d4a:	data_out=16'h4b5;
17'h3d4b:	data_out=16'h8a00;
17'h3d4c:	data_out=16'h8a00;
17'h3d4d:	data_out=16'h89ea;
17'h3d4e:	data_out=16'hd3;
17'h3d4f:	data_out=16'h8a00;
17'h3d50:	data_out=16'h9d5;
17'h3d51:	data_out=16'h8a00;
17'h3d52:	data_out=16'h82e2;
17'h3d53:	data_out=16'ha00;
17'h3d54:	data_out=16'h9c5;
17'h3d55:	data_out=16'h89f7;
17'h3d56:	data_out=16'h89f2;
17'h3d57:	data_out=16'h89fa;
17'h3d58:	data_out=16'h89ef;
17'h3d59:	data_out=16'h9f1;
17'h3d5a:	data_out=16'h89e6;
17'h3d5b:	data_out=16'ha00;
17'h3d5c:	data_out=16'h9e7;
17'h3d5d:	data_out=16'h88b8;
17'h3d5e:	data_out=16'h8299;
17'h3d5f:	data_out=16'h89ff;
17'h3d60:	data_out=16'h89ff;
17'h3d61:	data_out=16'ha00;
17'h3d62:	data_out=16'h89ef;
17'h3d63:	data_out=16'h89e4;
17'h3d64:	data_out=16'h89fd;
17'h3d65:	data_out=16'ha00;
17'h3d66:	data_out=16'ha00;
17'h3d67:	data_out=16'h65f;
17'h3d68:	data_out=16'h81df;
17'h3d69:	data_out=16'h8a00;
17'h3d6a:	data_out=16'h82be;
17'h3d6b:	data_out=16'h9e5;
17'h3d6c:	data_out=16'h89eb;
17'h3d6d:	data_out=16'h89e9;
17'h3d6e:	data_out=16'h82be;
17'h3d6f:	data_out=16'ha00;
17'h3d70:	data_out=16'h82a8;
17'h3d71:	data_out=16'h89f9;
17'h3d72:	data_out=16'h9aa;
17'h3d73:	data_out=16'ha00;
17'h3d74:	data_out=16'ha00;
17'h3d75:	data_out=16'h3df;
17'h3d76:	data_out=16'ha00;
17'h3d77:	data_out=16'h89ff;
17'h3d78:	data_out=16'ha00;
17'h3d79:	data_out=16'h873c;
17'h3d7a:	data_out=16'h89e4;
17'h3d7b:	data_out=16'h8158;
17'h3d7c:	data_out=16'h89fd;
17'h3d7d:	data_out=16'ha00;
17'h3d7e:	data_out=16'h8a00;
17'h3d7f:	data_out=16'h2b4;
17'h3d80:	data_out=16'h89fc;
17'h3d81:	data_out=16'h9f3;
17'h3d82:	data_out=16'h89b1;
17'h3d83:	data_out=16'h8a00;
17'h3d84:	data_out=16'ha00;
17'h3d85:	data_out=16'ha00;
17'h3d86:	data_out=16'h89fe;
17'h3d87:	data_out=16'h184;
17'h3d88:	data_out=16'h899b;
17'h3d89:	data_out=16'h89ff;
17'h3d8a:	data_out=16'ha00;
17'h3d8b:	data_out=16'h89d9;
17'h3d8c:	data_out=16'h48a;
17'h3d8d:	data_out=16'h8a00;
17'h3d8e:	data_out=16'h8249;
17'h3d8f:	data_out=16'h89f1;
17'h3d90:	data_out=16'h8642;
17'h3d91:	data_out=16'h8a6;
17'h3d92:	data_out=16'h8a00;
17'h3d93:	data_out=16'h8a00;
17'h3d94:	data_out=16'h89ed;
17'h3d95:	data_out=16'h848a;
17'h3d96:	data_out=16'h89ff;
17'h3d97:	data_out=16'h89ed;
17'h3d98:	data_out=16'h89fb;
17'h3d99:	data_out=16'ha00;
17'h3d9a:	data_out=16'ha00;
17'h3d9b:	data_out=16'h89d1;
17'h3d9c:	data_out=16'h6a5;
17'h3d9d:	data_out=16'h9f3;
17'h3d9e:	data_out=16'h89fd;
17'h3d9f:	data_out=16'h87b5;
17'h3da0:	data_out=16'h9e4;
17'h3da1:	data_out=16'h8205;
17'h3da2:	data_out=16'h89ee;
17'h3da3:	data_out=16'h8748;
17'h3da4:	data_out=16'h874a;
17'h3da5:	data_out=16'h89f3;
17'h3da6:	data_out=16'h89ff;
17'h3da7:	data_out=16'h9e5;
17'h3da8:	data_out=16'h810c;
17'h3da9:	data_out=16'h88b0;
17'h3daa:	data_out=16'h89da;
17'h3dab:	data_out=16'ha00;
17'h3dac:	data_out=16'h89ff;
17'h3dad:	data_out=16'h89f9;
17'h3dae:	data_out=16'h8992;
17'h3daf:	data_out=16'h9ed;
17'h3db0:	data_out=16'ha00;
17'h3db1:	data_out=16'h9dc;
17'h3db2:	data_out=16'ha00;
17'h3db3:	data_out=16'h89f6;
17'h3db4:	data_out=16'h9f0;
17'h3db5:	data_out=16'h9de;
17'h3db6:	data_out=16'h8981;
17'h3db7:	data_out=16'h8985;
17'h3db8:	data_out=16'h9a5;
17'h3db9:	data_out=16'h89fa;
17'h3dba:	data_out=16'h89f8;
17'h3dbb:	data_out=16'ha00;
17'h3dbc:	data_out=16'h8725;
17'h3dbd:	data_out=16'h963;
17'h3dbe:	data_out=16'h8108;
17'h3dbf:	data_out=16'ha00;
17'h3dc0:	data_out=16'ha00;
17'h3dc1:	data_out=16'h89dd;
17'h3dc2:	data_out=16'h89f2;
17'h3dc3:	data_out=16'h8108;
17'h3dc4:	data_out=16'h916;
17'h3dc5:	data_out=16'h8651;
17'h3dc6:	data_out=16'h8497;
17'h3dc7:	data_out=16'h89ff;
17'h3dc8:	data_out=16'h8a00;
17'h3dc9:	data_out=16'h89ef;
17'h3dca:	data_out=16'h839;
17'h3dcb:	data_out=16'h8a00;
17'h3dcc:	data_out=16'h89fc;
17'h3dcd:	data_out=16'h89c7;
17'h3dce:	data_out=16'h38b;
17'h3dcf:	data_out=16'h89f4;
17'h3dd0:	data_out=16'h1e5;
17'h3dd1:	data_out=16'h8a00;
17'h3dd2:	data_out=16'h8394;
17'h3dd3:	data_out=16'ha00;
17'h3dd4:	data_out=16'h9f0;
17'h3dd5:	data_out=16'h8a00;
17'h3dd6:	data_out=16'h89bd;
17'h3dd7:	data_out=16'h892b;
17'h3dd8:	data_out=16'h89ec;
17'h3dd9:	data_out=16'h9ef;
17'h3dda:	data_out=16'h89e9;
17'h3ddb:	data_out=16'ha00;
17'h3ddc:	data_out=16'h9d1;
17'h3ddd:	data_out=16'h8598;
17'h3dde:	data_out=16'h9c4;
17'h3ddf:	data_out=16'h89f8;
17'h3de0:	data_out=16'h89d5;
17'h3de1:	data_out=16'ha00;
17'h3de2:	data_out=16'h89dc;
17'h3de3:	data_out=16'h89cf;
17'h3de4:	data_out=16'h9c8;
17'h3de5:	data_out=16'ha00;
17'h3de6:	data_out=16'ha00;
17'h3de7:	data_out=16'h9fa;
17'h3de8:	data_out=16'h81c2;
17'h3de9:	data_out=16'h89f4;
17'h3dea:	data_out=16'h826a;
17'h3deb:	data_out=16'h9e1;
17'h3dec:	data_out=16'h89b7;
17'h3ded:	data_out=16'h89de;
17'h3dee:	data_out=16'h826b;
17'h3def:	data_out=16'ha00;
17'h3df0:	data_out=16'h8262;
17'h3df1:	data_out=16'h89ee;
17'h3df2:	data_out=16'h9d1;
17'h3df3:	data_out=16'ha00;
17'h3df4:	data_out=16'ha00;
17'h3df5:	data_out=16'h33e;
17'h3df6:	data_out=16'ha00;
17'h3df7:	data_out=16'h89ff;
17'h3df8:	data_out=16'ha00;
17'h3df9:	data_out=16'h87ba;
17'h3dfa:	data_out=16'h89d6;
17'h3dfb:	data_out=16'h810a;
17'h3dfc:	data_out=16'h89f9;
17'h3dfd:	data_out=16'h751;
17'h3dfe:	data_out=16'h8a00;
17'h3dff:	data_out=16'h82f2;
17'h3e00:	data_out=16'h89fd;
17'h3e01:	data_out=16'h9f5;
17'h3e02:	data_out=16'h89df;
17'h3e03:	data_out=16'h8a00;
17'h3e04:	data_out=16'ha00;
17'h3e05:	data_out=16'ha00;
17'h3e06:	data_out=16'h89f1;
17'h3e07:	data_out=16'h86d9;
17'h3e08:	data_out=16'h89dc;
17'h3e09:	data_out=16'h89fc;
17'h3e0a:	data_out=16'ha00;
17'h3e0b:	data_out=16'h89f0;
17'h3e0c:	data_out=16'h8996;
17'h3e0d:	data_out=16'h8a00;
17'h3e0e:	data_out=16'h839d;
17'h3e0f:	data_out=16'h89ee;
17'h3e10:	data_out=16'h890c;
17'h3e11:	data_out=16'h74d;
17'h3e12:	data_out=16'h8a00;
17'h3e13:	data_out=16'h89ff;
17'h3e14:	data_out=16'h89fb;
17'h3e15:	data_out=16'h859f;
17'h3e16:	data_out=16'h89ff;
17'h3e17:	data_out=16'h89fd;
17'h3e18:	data_out=16'h8a00;
17'h3e19:	data_out=16'ha00;
17'h3e1a:	data_out=16'ha00;
17'h3e1b:	data_out=16'h89e3;
17'h3e1c:	data_out=16'h4a8;
17'h3e1d:	data_out=16'h9ea;
17'h3e1e:	data_out=16'h89fc;
17'h3e1f:	data_out=16'h85d4;
17'h3e20:	data_out=16'h9ad;
17'h3e21:	data_out=16'h8341;
17'h3e22:	data_out=16'h89d4;
17'h3e23:	data_out=16'h8993;
17'h3e24:	data_out=16'h8993;
17'h3e25:	data_out=16'h89d5;
17'h3e26:	data_out=16'h89de;
17'h3e27:	data_out=16'h95f;
17'h3e28:	data_out=16'h81ff;
17'h3e29:	data_out=16'h8563;
17'h3e2a:	data_out=16'h89ec;
17'h3e2b:	data_out=16'ha00;
17'h3e2c:	data_out=16'h89ff;
17'h3e2d:	data_out=16'h89fc;
17'h3e2e:	data_out=16'h89b9;
17'h3e2f:	data_out=16'h9cd;
17'h3e30:	data_out=16'ha00;
17'h3e31:	data_out=16'h9cd;
17'h3e32:	data_out=16'ha00;
17'h3e33:	data_out=16'h89fa;
17'h3e34:	data_out=16'h9ef;
17'h3e35:	data_out=16'h88c;
17'h3e36:	data_out=16'h89e0;
17'h3e37:	data_out=16'h89d7;
17'h3e38:	data_out=16'h970;
17'h3e39:	data_out=16'h89fc;
17'h3e3a:	data_out=16'h89fd;
17'h3e3b:	data_out=16'ha00;
17'h3e3c:	data_out=16'h84d5;
17'h3e3d:	data_out=16'h8fc;
17'h3e3e:	data_out=16'h81f8;
17'h3e3f:	data_out=16'ha00;
17'h3e40:	data_out=16'ha00;
17'h3e41:	data_out=16'h89de;
17'h3e42:	data_out=16'h89e7;
17'h3e43:	data_out=16'ha00;
17'h3e44:	data_out=16'h8bd;
17'h3e45:	data_out=16'h8724;
17'h3e46:	data_out=16'h8919;
17'h3e47:	data_out=16'h89ff;
17'h3e48:	data_out=16'h89ff;
17'h3e49:	data_out=16'h89d6;
17'h3e4a:	data_out=16'h24a;
17'h3e4b:	data_out=16'h8a00;
17'h3e4c:	data_out=16'h89e2;
17'h3e4d:	data_out=16'h88b3;
17'h3e4e:	data_out=16'haf;
17'h3e4f:	data_out=16'h89e9;
17'h3e50:	data_out=16'h21c;
17'h3e51:	data_out=16'h8a00;
17'h3e52:	data_out=16'h868a;
17'h3e53:	data_out=16'h9e9;
17'h3e54:	data_out=16'h9cf;
17'h3e55:	data_out=16'h89fb;
17'h3e56:	data_out=16'h89ca;
17'h3e57:	data_out=16'h89f2;
17'h3e58:	data_out=16'h89f2;
17'h3e59:	data_out=16'h9f5;
17'h3e5a:	data_out=16'h89f3;
17'h3e5b:	data_out=16'ha00;
17'h3e5c:	data_out=16'h9c2;
17'h3e5d:	data_out=16'h879a;
17'h3e5e:	data_out=16'h9c5;
17'h3e5f:	data_out=16'h89fe;
17'h3e60:	data_out=16'h89cd;
17'h3e61:	data_out=16'ha00;
17'h3e62:	data_out=16'h89ef;
17'h3e63:	data_out=16'h89df;
17'h3e64:	data_out=16'h99c;
17'h3e65:	data_out=16'ha00;
17'h3e66:	data_out=16'ha00;
17'h3e67:	data_out=16'h9f2;
17'h3e68:	data_out=16'h82df;
17'h3e69:	data_out=16'h8a00;
17'h3e6a:	data_out=16'h83d7;
17'h3e6b:	data_out=16'h9bf;
17'h3e6c:	data_out=16'h89fc;
17'h3e6d:	data_out=16'h89ed;
17'h3e6e:	data_out=16'h83d6;
17'h3e6f:	data_out=16'ha00;
17'h3e70:	data_out=16'h83be;
17'h3e71:	data_out=16'h89f1;
17'h3e72:	data_out=16'h9d8;
17'h3e73:	data_out=16'ha00;
17'h3e74:	data_out=16'ha00;
17'h3e75:	data_out=16'h752;
17'h3e76:	data_out=16'ha00;
17'h3e77:	data_out=16'h89fb;
17'h3e78:	data_out=16'ha00;
17'h3e79:	data_out=16'h89d5;
17'h3e7a:	data_out=16'h89e5;
17'h3e7b:	data_out=16'h81f8;
17'h3e7c:	data_out=16'h89fd;
17'h3e7d:	data_out=16'h9d8;
17'h3e7e:	data_out=16'h8a00;
17'h3e7f:	data_out=16'h82ac;
17'h3e80:	data_out=16'h89fd;
17'h3e81:	data_out=16'h9fa;
17'h3e82:	data_out=16'h89c8;
17'h3e83:	data_out=16'h89fc;
17'h3e84:	data_out=16'ha00;
17'h3e85:	data_out=16'ha00;
17'h3e86:	data_out=16'h89ee;
17'h3e87:	data_out=16'h88da;
17'h3e88:	data_out=16'h89cd;
17'h3e89:	data_out=16'h89fb;
17'h3e8a:	data_out=16'ha00;
17'h3e8b:	data_out=16'h81f6;
17'h3e8c:	data_out=16'h89c7;
17'h3e8d:	data_out=16'h8a00;
17'h3e8e:	data_out=16'h89e3;
17'h3e8f:	data_out=16'h89df;
17'h3e90:	data_out=16'h89e3;
17'h3e91:	data_out=16'h744;
17'h3e92:	data_out=16'h8a00;
17'h3e93:	data_out=16'h89f9;
17'h3e94:	data_out=16'h89de;
17'h3e95:	data_out=16'h89de;
17'h3e96:	data_out=16'h89fd;
17'h3e97:	data_out=16'h89b9;
17'h3e98:	data_out=16'h8a00;
17'h3e99:	data_out=16'ha00;
17'h3e9a:	data_out=16'ha00;
17'h3e9b:	data_out=16'h89de;
17'h3e9c:	data_out=16'h64;
17'h3e9d:	data_out=16'h9ef;
17'h3e9e:	data_out=16'h89f6;
17'h3e9f:	data_out=16'h812f;
17'h3ea0:	data_out=16'h9d4;
17'h3ea1:	data_out=16'h89d1;
17'h3ea2:	data_out=16'h89e1;
17'h3ea3:	data_out=16'h899d;
17'h3ea4:	data_out=16'h899e;
17'h3ea5:	data_out=16'h89e1;
17'h3ea6:	data_out=16'h89e2;
17'h3ea7:	data_out=16'h9af;
17'h3ea8:	data_out=16'h8993;
17'h3ea9:	data_out=16'h8863;
17'h3eaa:	data_out=16'h89df;
17'h3eab:	data_out=16'ha00;
17'h3eac:	data_out=16'h89fd;
17'h3ead:	data_out=16'h89fb;
17'h3eae:	data_out=16'h89a9;
17'h3eaf:	data_out=16'h9d2;
17'h3eb0:	data_out=16'ha00;
17'h3eb1:	data_out=16'h9ea;
17'h3eb2:	data_out=16'ha00;
17'h3eb3:	data_out=16'h89f5;
17'h3eb4:	data_out=16'h9f3;
17'h3eb5:	data_out=16'h983;
17'h3eb6:	data_out=16'h89cf;
17'h3eb7:	data_out=16'h89b6;
17'h3eb8:	data_out=16'h837;
17'h3eb9:	data_out=16'h89f7;
17'h3eba:	data_out=16'h89fa;
17'h3ebb:	data_out=16'ha00;
17'h3ebc:	data_out=16'h8649;
17'h3ebd:	data_out=16'h7ee;
17'h3ebe:	data_out=16'h8991;
17'h3ebf:	data_out=16'ha00;
17'h3ec0:	data_out=16'ha00;
17'h3ec1:	data_out=16'h89cb;
17'h3ec2:	data_out=16'h8a00;
17'h3ec3:	data_out=16'ha00;
17'h3ec4:	data_out=16'h9ec;
17'h3ec5:	data_out=16'h89f3;
17'h3ec6:	data_out=16'h89d7;
17'h3ec7:	data_out=16'h89fe;
17'h3ec8:	data_out=16'h89fb;
17'h3ec9:	data_out=16'h89e3;
17'h3eca:	data_out=16'h28f;
17'h3ecb:	data_out=16'h8a00;
17'h3ecc:	data_out=16'h89f6;
17'h3ecd:	data_out=16'h89cc;
17'h3ece:	data_out=16'h8363;
17'h3ecf:	data_out=16'h8a00;
17'h3ed0:	data_out=16'h2b4;
17'h3ed1:	data_out=16'h8a00;
17'h3ed2:	data_out=16'h8993;
17'h3ed3:	data_out=16'h9ff;
17'h3ed4:	data_out=16'h9df;
17'h3ed5:	data_out=16'h89e1;
17'h3ed6:	data_out=16'h89c3;
17'h3ed7:	data_out=16'h89d8;
17'h3ed8:	data_out=16'h89f3;
17'h3ed9:	data_out=16'h9f5;
17'h3eda:	data_out=16'h89e3;
17'h3edb:	data_out=16'ha00;
17'h3edc:	data_out=16'h9e0;
17'h3edd:	data_out=16'h89c5;
17'h3ede:	data_out=16'h983;
17'h3edf:	data_out=16'h89fd;
17'h3ee0:	data_out=16'h89ca;
17'h3ee1:	data_out=16'ha00;
17'h3ee2:	data_out=16'h89b1;
17'h3ee3:	data_out=16'h89ca;
17'h3ee4:	data_out=16'h9d2;
17'h3ee5:	data_out=16'ha00;
17'h3ee6:	data_out=16'ha00;
17'h3ee7:	data_out=16'h9fb;
17'h3ee8:	data_out=16'h89b8;
17'h3ee9:	data_out=16'h8a00;
17'h3eea:	data_out=16'h89e4;
17'h3eeb:	data_out=16'h9cf;
17'h3eec:	data_out=16'h89fd;
17'h3eed:	data_out=16'h89da;
17'h3eee:	data_out=16'h89e4;
17'h3eef:	data_out=16'ha00;
17'h3ef0:	data_out=16'h89e3;
17'h3ef1:	data_out=16'h89df;
17'h3ef2:	data_out=16'h9db;
17'h3ef3:	data_out=16'ha00;
17'h3ef4:	data_out=16'h9ff;
17'h3ef5:	data_out=16'h839;
17'h3ef6:	data_out=16'ha00;
17'h3ef7:	data_out=16'h89fb;
17'h3ef8:	data_out=16'ha00;
17'h3ef9:	data_out=16'h89df;
17'h3efa:	data_out=16'h89c7;
17'h3efb:	data_out=16'h8991;
17'h3efc:	data_out=16'h89fd;
17'h3efd:	data_out=16'ha00;
17'h3efe:	data_out=16'h8a00;
17'h3eff:	data_out=16'h8527;
17'h3f00:	data_out=16'h89fb;
17'h3f01:	data_out=16'h9ee;
17'h3f02:	data_out=16'h89ab;
17'h3f03:	data_out=16'h89fc;
17'h3f04:	data_out=16'ha00;
17'h3f05:	data_out=16'ha00;
17'h3f06:	data_out=16'h89ed;
17'h3f07:	data_out=16'h89df;
17'h3f08:	data_out=16'h89ba;
17'h3f09:	data_out=16'h89ff;
17'h3f0a:	data_out=16'ha00;
17'h3f0b:	data_out=16'h89fc;
17'h3f0c:	data_out=16'h89f6;
17'h3f0d:	data_out=16'h8a00;
17'h3f0e:	data_out=16'h89c9;
17'h3f0f:	data_out=16'h89e9;
17'h3f10:	data_out=16'h89f0;
17'h3f11:	data_out=16'h615;
17'h3f12:	data_out=16'h8a00;
17'h3f13:	data_out=16'h89be;
17'h3f14:	data_out=16'h89f3;
17'h3f15:	data_out=16'h88f4;
17'h3f16:	data_out=16'h89b9;
17'h3f17:	data_out=16'h89cc;
17'h3f18:	data_out=16'h8a00;
17'h3f19:	data_out=16'ha00;
17'h3f1a:	data_out=16'ha00;
17'h3f1b:	data_out=16'h89bb;
17'h3f1c:	data_out=16'h84bd;
17'h3f1d:	data_out=16'h9cb;
17'h3f1e:	data_out=16'h89f7;
17'h3f1f:	data_out=16'h8395;
17'h3f20:	data_out=16'h9e0;
17'h3f21:	data_out=16'h89bd;
17'h3f22:	data_out=16'h89f4;
17'h3f23:	data_out=16'h88b1;
17'h3f24:	data_out=16'h88c0;
17'h3f25:	data_out=16'h89e7;
17'h3f26:	data_out=16'h8a00;
17'h3f27:	data_out=16'h9d3;
17'h3f28:	data_out=16'h8981;
17'h3f29:	data_out=16'h89d8;
17'h3f2a:	data_out=16'h89d5;
17'h3f2b:	data_out=16'h9f5;
17'h3f2c:	data_out=16'h89be;
17'h3f2d:	data_out=16'h8a00;
17'h3f2e:	data_out=16'h89c7;
17'h3f2f:	data_out=16'h88e5;
17'h3f30:	data_out=16'ha00;
17'h3f31:	data_out=16'h9e8;
17'h3f32:	data_out=16'ha00;
17'h3f33:	data_out=16'h89f5;
17'h3f34:	data_out=16'h9d2;
17'h3f35:	data_out=16'h9da;
17'h3f36:	data_out=16'h89b8;
17'h3f37:	data_out=16'h899b;
17'h3f38:	data_out=16'h8013;
17'h3f39:	data_out=16'h89f9;
17'h3f3a:	data_out=16'h89fd;
17'h3f3b:	data_out=16'ha00;
17'h3f3c:	data_out=16'h8795;
17'h3f3d:	data_out=16'h87a6;
17'h3f3e:	data_out=16'h8980;
17'h3f3f:	data_out=16'ha00;
17'h3f40:	data_out=16'ha00;
17'h3f41:	data_out=16'h89aa;
17'h3f42:	data_out=16'h8a00;
17'h3f43:	data_out=16'ha00;
17'h3f44:	data_out=16'h9fc;
17'h3f45:	data_out=16'h88f6;
17'h3f46:	data_out=16'h89da;
17'h3f47:	data_out=16'h8a00;
17'h3f48:	data_out=16'h89fc;
17'h3f49:	data_out=16'h89e6;
17'h3f4a:	data_out=16'h118;
17'h3f4b:	data_out=16'h8a00;
17'h3f4c:	data_out=16'h89f4;
17'h3f4d:	data_out=16'h89e2;
17'h3f4e:	data_out=16'h89bf;
17'h3f4f:	data_out=16'h8a00;
17'h3f50:	data_out=16'h1d2;
17'h3f51:	data_out=16'h8a00;
17'h3f52:	data_out=16'h89ac;
17'h3f53:	data_out=16'h4f5;
17'h3f54:	data_out=16'h87c1;
17'h3f55:	data_out=16'h89e4;
17'h3f56:	data_out=16'h8989;
17'h3f57:	data_out=16'h89b4;
17'h3f58:	data_out=16'h89cd;
17'h3f59:	data_out=16'ha00;
17'h3f5a:	data_out=16'h89de;
17'h3f5b:	data_out=16'ha00;
17'h3f5c:	data_out=16'h9fa;
17'h3f5d:	data_out=16'h899b;
17'h3f5e:	data_out=16'h88af;
17'h3f5f:	data_out=16'h89fc;
17'h3f60:	data_out=16'h8a00;
17'h3f61:	data_out=16'ha00;
17'h3f62:	data_out=16'h89d5;
17'h3f63:	data_out=16'h89ec;
17'h3f64:	data_out=16'h99e;
17'h3f65:	data_out=16'ha00;
17'h3f66:	data_out=16'ha00;
17'h3f67:	data_out=16'h9f0;
17'h3f68:	data_out=16'h89a7;
17'h3f69:	data_out=16'h8a00;
17'h3f6a:	data_out=16'h89c9;
17'h3f6b:	data_out=16'h9fe;
17'h3f6c:	data_out=16'h89c2;
17'h3f6d:	data_out=16'h89f3;
17'h3f6e:	data_out=16'h89c9;
17'h3f6f:	data_out=16'ha00;
17'h3f70:	data_out=16'h89c8;
17'h3f71:	data_out=16'h89e0;
17'h3f72:	data_out=16'h9f9;
17'h3f73:	data_out=16'ha00;
17'h3f74:	data_out=16'ha00;
17'h3f75:	data_out=16'h9ff;
17'h3f76:	data_out=16'h9fb;
17'h3f77:	data_out=16'h8a00;
17'h3f78:	data_out=16'ha00;
17'h3f79:	data_out=16'h89f0;
17'h3f7a:	data_out=16'h89ef;
17'h3f7b:	data_out=16'h897f;
17'h3f7c:	data_out=16'h89ff;
17'h3f7d:	data_out=16'ha00;
17'h3f7e:	data_out=16'h8a00;
17'h3f7f:	data_out=16'h8242;
17'h3f80:	data_out=16'h89fd;
17'h3f81:	data_out=16'h9f2;
17'h3f82:	data_out=16'h899b;
17'h3f83:	data_out=16'h8a00;
17'h3f84:	data_out=16'ha00;
17'h3f85:	data_out=16'ha00;
17'h3f86:	data_out=16'h899b;
17'h3f87:	data_out=16'h89df;
17'h3f88:	data_out=16'h89bb;
17'h3f89:	data_out=16'h8a00;
17'h3f8a:	data_out=16'ha00;
17'h3f8b:	data_out=16'h8a00;
17'h3f8c:	data_out=16'h89ec;
17'h3f8d:	data_out=16'h8a00;
17'h3f8e:	data_out=16'h897b;
17'h3f8f:	data_out=16'h89d2;
17'h3f90:	data_out=16'h89fc;
17'h3f91:	data_out=16'h46b;
17'h3f92:	data_out=16'h8a00;
17'h3f93:	data_out=16'h86cb;
17'h3f94:	data_out=16'h89e8;
17'h3f95:	data_out=16'h8917;
17'h3f96:	data_out=16'h8981;
17'h3f97:	data_out=16'h89cf;
17'h3f98:	data_out=16'h8a00;
17'h3f99:	data_out=16'ha00;
17'h3f9a:	data_out=16'ha00;
17'h3f9b:	data_out=16'h89a8;
17'h3f9c:	data_out=16'h89d5;
17'h3f9d:	data_out=16'h9c0;
17'h3f9e:	data_out=16'h89e7;
17'h3f9f:	data_out=16'h8684;
17'h3fa0:	data_out=16'h83df;
17'h3fa1:	data_out=16'h896f;
17'h3fa2:	data_out=16'h89fe;
17'h3fa3:	data_out=16'h9fa;
17'h3fa4:	data_out=16'h9fa;
17'h3fa5:	data_out=16'h89ef;
17'h3fa6:	data_out=16'h8a00;
17'h3fa7:	data_out=16'h631;
17'h3fa8:	data_out=16'h8924;
17'h3fa9:	data_out=16'h89e5;
17'h3faa:	data_out=16'h89a5;
17'h3fab:	data_out=16'h9d5;
17'h3fac:	data_out=16'h899c;
17'h3fad:	data_out=16'h8a00;
17'h3fae:	data_out=16'h89c8;
17'h3faf:	data_out=16'h8990;
17'h3fb0:	data_out=16'ha00;
17'h3fb1:	data_out=16'ha00;
17'h3fb2:	data_out=16'ha00;
17'h3fb3:	data_out=16'h89fb;
17'h3fb4:	data_out=16'h9d1;
17'h3fb5:	data_out=16'h8ac;
17'h3fb6:	data_out=16'h89a4;
17'h3fb7:	data_out=16'h898c;
17'h3fb8:	data_out=16'h89fd;
17'h3fb9:	data_out=16'h89ff;
17'h3fba:	data_out=16'h8a00;
17'h3fbb:	data_out=16'ha00;
17'h3fbc:	data_out=16'h83e8;
17'h3fbd:	data_out=16'h89cb;
17'h3fbe:	data_out=16'h8921;
17'h3fbf:	data_out=16'ha00;
17'h3fc0:	data_out=16'ha00;
17'h3fc1:	data_out=16'h899c;
17'h3fc2:	data_out=16'h8a00;
17'h3fc3:	data_out=16'ha00;
17'h3fc4:	data_out=16'ha00;
17'h3fc5:	data_out=16'h8912;
17'h3fc6:	data_out=16'h89dd;
17'h3fc7:	data_out=16'h8a00;
17'h3fc8:	data_out=16'h89fe;
17'h3fc9:	data_out=16'h89f7;
17'h3fca:	data_out=16'h472;
17'h3fcb:	data_out=16'h8a00;
17'h3fcc:	data_out=16'h89f8;
17'h3fcd:	data_out=16'h89f4;
17'h3fce:	data_out=16'h89e5;
17'h3fcf:	data_out=16'h8a00;
17'h3fd0:	data_out=16'h81e0;
17'h3fd1:	data_out=16'h89e2;
17'h3fd2:	data_out=16'h77c;
17'h3fd3:	data_out=16'h121;
17'h3fd4:	data_out=16'h89a4;
17'h3fd5:	data_out=16'h89be;
17'h3fd6:	data_out=16'h897d;
17'h3fd7:	data_out=16'h89d1;
17'h3fd8:	data_out=16'h89a8;
17'h3fd9:	data_out=16'ha00;
17'h3fda:	data_out=16'h89c9;
17'h3fdb:	data_out=16'ha00;
17'h3fdc:	data_out=16'h9fb;
17'h3fdd:	data_out=16'h89ab;
17'h3fde:	data_out=16'h88ec;
17'h3fdf:	data_out=16'h89ff;
17'h3fe0:	data_out=16'h8a00;
17'h3fe1:	data_out=16'ha00;
17'h3fe2:	data_out=16'h89b1;
17'h3fe3:	data_out=16'h89f1;
17'h3fe4:	data_out=16'h89b7;
17'h3fe5:	data_out=16'ha00;
17'h3fe6:	data_out=16'ha00;
17'h3fe7:	data_out=16'h5;
17'h3fe8:	data_out=16'h8956;
17'h3fe9:	data_out=16'h8a00;
17'h3fea:	data_out=16'h8983;
17'h3feb:	data_out=16'ha00;
17'h3fec:	data_out=16'h89f5;
17'h3fed:	data_out=16'h89f7;
17'h3fee:	data_out=16'h8983;
17'h3fef:	data_out=16'ha00;
17'h3ff0:	data_out=16'h897d;
17'h3ff1:	data_out=16'h89c5;
17'h3ff2:	data_out=16'ha00;
17'h3ff3:	data_out=16'ha00;
17'h3ff4:	data_out=16'ha00;
17'h3ff5:	data_out=16'ha00;
17'h3ff6:	data_out=16'h9cc;
17'h3ff7:	data_out=16'h8a00;
17'h3ff8:	data_out=16'ha00;
17'h3ff9:	data_out=16'h8a00;
17'h3ffa:	data_out=16'h89da;
17'h3ffb:	data_out=16'h8920;
17'h3ffc:	data_out=16'h8a00;
17'h3ffd:	data_out=16'h780;
17'h3ffe:	data_out=16'h8a00;
17'h3fff:	data_out=16'h8390;
17'h4000:	data_out=16'h8a00;
17'h4001:	data_out=16'h9fc;
17'h4002:	data_out=16'h899b;
17'h4003:	data_out=16'h8a00;
17'h4004:	data_out=16'ha00;
17'h4005:	data_out=16'ha00;
17'h4006:	data_out=16'h850;
17'h4007:	data_out=16'h8534;
17'h4008:	data_out=16'h89d5;
17'h4009:	data_out=16'h89fd;
17'h400a:	data_out=16'ha00;
17'h400b:	data_out=16'h8a00;
17'h400c:	data_out=16'h89f1;
17'h400d:	data_out=16'h8a00;
17'h400e:	data_out=16'h1be;
17'h400f:	data_out=16'h89de;
17'h4010:	data_out=16'h89fa;
17'h4011:	data_out=16'h5f4;
17'h4012:	data_out=16'h8a00;
17'h4013:	data_out=16'h839c;
17'h4014:	data_out=16'h8a00;
17'h4015:	data_out=16'h89eb;
17'h4016:	data_out=16'h89e1;
17'h4017:	data_out=16'h89ec;
17'h4018:	data_out=16'h8a00;
17'h4019:	data_out=16'ha00;
17'h401a:	data_out=16'ha00;
17'h401b:	data_out=16'h89d6;
17'h401c:	data_out=16'h89f6;
17'h401d:	data_out=16'h8cc;
17'h401e:	data_out=16'h8a00;
17'h401f:	data_out=16'h8948;
17'h4020:	data_out=16'h8904;
17'h4021:	data_out=16'h25a;
17'h4022:	data_out=16'h89fb;
17'h4023:	data_out=16'ha00;
17'h4024:	data_out=16'ha00;
17'h4025:	data_out=16'h8909;
17'h4026:	data_out=16'h8a00;
17'h4027:	data_out=16'h59a;
17'h4028:	data_out=16'h42b;
17'h4029:	data_out=16'h89e6;
17'h402a:	data_out=16'h89ba;
17'h402b:	data_out=16'h7ce;
17'h402c:	data_out=16'h89f0;
17'h402d:	data_out=16'h8a00;
17'h402e:	data_out=16'h89d0;
17'h402f:	data_out=16'h89cc;
17'h4030:	data_out=16'ha00;
17'h4031:	data_out=16'ha00;
17'h4032:	data_out=16'ha00;
17'h4033:	data_out=16'h8a00;
17'h4034:	data_out=16'h874;
17'h4035:	data_out=16'h837;
17'h4036:	data_out=16'h89bd;
17'h4037:	data_out=16'h898f;
17'h4038:	data_out=16'h89fb;
17'h4039:	data_out=16'h8a00;
17'h403a:	data_out=16'h89fd;
17'h403b:	data_out=16'ha00;
17'h403c:	data_out=16'h427;
17'h403d:	data_out=16'h89f1;
17'h403e:	data_out=16'h43d;
17'h403f:	data_out=16'ha00;
17'h4040:	data_out=16'ha00;
17'h4041:	data_out=16'h89ba;
17'h4042:	data_out=16'h8a00;
17'h4043:	data_out=16'ha00;
17'h4044:	data_out=16'ha00;
17'h4045:	data_out=16'h89eb;
17'h4046:	data_out=16'h89e1;
17'h4047:	data_out=16'h8a00;
17'h4048:	data_out=16'h85de;
17'h4049:	data_out=16'h89e9;
17'h404a:	data_out=16'ha00;
17'h404b:	data_out=16'h8a00;
17'h404c:	data_out=16'h89dc;
17'h404d:	data_out=16'h88fc;
17'h404e:	data_out=16'h89fb;
17'h404f:	data_out=16'h89fe;
17'h4050:	data_out=16'h857e;
17'h4051:	data_out=16'h8a00;
17'h4052:	data_out=16'h9d4;
17'h4053:	data_out=16'h751;
17'h4054:	data_out=16'h89c8;
17'h4055:	data_out=16'h89e0;
17'h4056:	data_out=16'h8980;
17'h4057:	data_out=16'h89bd;
17'h4058:	data_out=16'h89c4;
17'h4059:	data_out=16'ha00;
17'h405a:	data_out=16'h89d9;
17'h405b:	data_out=16'ha00;
17'h405c:	data_out=16'h9f8;
17'h405d:	data_out=16'h89b3;
17'h405e:	data_out=16'h8812;
17'h405f:	data_out=16'h8a00;
17'h4060:	data_out=16'h8a00;
17'h4061:	data_out=16'ha00;
17'h4062:	data_out=16'h89eb;
17'h4063:	data_out=16'h8a00;
17'h4064:	data_out=16'h89ff;
17'h4065:	data_out=16'ha00;
17'h4066:	data_out=16'ha00;
17'h4067:	data_out=16'h9c8;
17'h4068:	data_out=16'h2d8;
17'h4069:	data_out=16'h8a00;
17'h406a:	data_out=16'h13d;
17'h406b:	data_out=16'ha00;
17'h406c:	data_out=16'h89ff;
17'h406d:	data_out=16'h8a00;
17'h406e:	data_out=16'h144;
17'h406f:	data_out=16'ha00;
17'h4070:	data_out=16'h199;
17'h4071:	data_out=16'h89cd;
17'h4072:	data_out=16'ha00;
17'h4073:	data_out=16'ha00;
17'h4074:	data_out=16'ha00;
17'h4075:	data_out=16'ha00;
17'h4076:	data_out=16'h898;
17'h4077:	data_out=16'h8a00;
17'h4078:	data_out=16'ha00;
17'h4079:	data_out=16'h8a00;
17'h407a:	data_out=16'h89fb;
17'h407b:	data_out=16'h446;
17'h407c:	data_out=16'h89ff;
17'h407d:	data_out=16'h99d;
17'h407e:	data_out=16'h8a00;
17'h407f:	data_out=16'h822f;
17'h4080:	data_out=16'h8a00;
17'h4081:	data_out=16'h9ff;
17'h4082:	data_out=16'h89a6;
17'h4083:	data_out=16'h8a00;
17'h4084:	data_out=16'ha00;
17'h4085:	data_out=16'ha00;
17'h4086:	data_out=16'h7c9;
17'h4087:	data_out=16'h936;
17'h4088:	data_out=16'h89ea;
17'h4089:	data_out=16'h89fc;
17'h408a:	data_out=16'ha00;
17'h408b:	data_out=16'h8a00;
17'h408c:	data_out=16'h30e;
17'h408d:	data_out=16'h8a00;
17'h408e:	data_out=16'h9d4;
17'h408f:	data_out=16'h89e6;
17'h4090:	data_out=16'h89fc;
17'h4091:	data_out=16'h9f5;
17'h4092:	data_out=16'h8a00;
17'h4093:	data_out=16'h863b;
17'h4094:	data_out=16'h89ff;
17'h4095:	data_out=16'h89f3;
17'h4096:	data_out=16'h89fe;
17'h4097:	data_out=16'h89ff;
17'h4098:	data_out=16'h8a00;
17'h4099:	data_out=16'ha00;
17'h409a:	data_out=16'ha00;
17'h409b:	data_out=16'h89ff;
17'h409c:	data_out=16'h8a00;
17'h409d:	data_out=16'h86c;
17'h409e:	data_out=16'h89ff;
17'h409f:	data_out=16'h89fc;
17'h40a0:	data_out=16'h89e0;
17'h40a1:	data_out=16'h9ff;
17'h40a2:	data_out=16'h81d;
17'h40a3:	data_out=16'ha00;
17'h40a4:	data_out=16'ha00;
17'h40a5:	data_out=16'h408;
17'h40a6:	data_out=16'h89f0;
17'h40a7:	data_out=16'h875;
17'h40a8:	data_out=16'h9ff;
17'h40a9:	data_out=16'h89f2;
17'h40aa:	data_out=16'h89cb;
17'h40ab:	data_out=16'h625;
17'h40ac:	data_out=16'h89fe;
17'h40ad:	data_out=16'h89ff;
17'h40ae:	data_out=16'h89f3;
17'h40af:	data_out=16'h89fd;
17'h40b0:	data_out=16'ha00;
17'h40b1:	data_out=16'ha00;
17'h40b2:	data_out=16'ha00;
17'h40b3:	data_out=16'h8a00;
17'h40b4:	data_out=16'h8952;
17'h40b5:	data_out=16'h9ec;
17'h40b6:	data_out=16'h89d5;
17'h40b7:	data_out=16'h87b0;
17'h40b8:	data_out=16'h890e;
17'h40b9:	data_out=16'h8a00;
17'h40ba:	data_out=16'h89fa;
17'h40bb:	data_out=16'ha00;
17'h40bc:	data_out=16'hd3;
17'h40bd:	data_out=16'h89f4;
17'h40be:	data_out=16'h9ff;
17'h40bf:	data_out=16'ha00;
17'h40c0:	data_out=16'ha00;
17'h40c1:	data_out=16'h89eb;
17'h40c2:	data_out=16'h8a00;
17'h40c3:	data_out=16'h9f6;
17'h40c4:	data_out=16'ha00;
17'h40c5:	data_out=16'h89f5;
17'h40c6:	data_out=16'h89b5;
17'h40c7:	data_out=16'h8a00;
17'h40c8:	data_out=16'h35d;
17'h40c9:	data_out=16'h562;
17'h40ca:	data_out=16'ha00;
17'h40cb:	data_out=16'h8a00;
17'h40cc:	data_out=16'h9d7;
17'h40cd:	data_out=16'h95d;
17'h40ce:	data_out=16'h8a00;
17'h40cf:	data_out=16'h8090;
17'h40d0:	data_out=16'h89fc;
17'h40d1:	data_out=16'h8a00;
17'h40d2:	data_out=16'h9ef;
17'h40d3:	data_out=16'h83a;
17'h40d4:	data_out=16'h89f0;
17'h40d5:	data_out=16'h89ff;
17'h40d6:	data_out=16'h86ef;
17'h40d7:	data_out=16'h89ac;
17'h40d8:	data_out=16'h89f3;
17'h40d9:	data_out=16'ha00;
17'h40da:	data_out=16'h8a00;
17'h40db:	data_out=16'ha00;
17'h40dc:	data_out=16'h86b7;
17'h40dd:	data_out=16'h880a;
17'h40de:	data_out=16'h8908;
17'h40df:	data_out=16'h89ff;
17'h40e0:	data_out=16'h89fd;
17'h40e1:	data_out=16'ha00;
17'h40e2:	data_out=16'h89fe;
17'h40e3:	data_out=16'h89ff;
17'h40e4:	data_out=16'h89fe;
17'h40e5:	data_out=16'ha00;
17'h40e6:	data_out=16'ha00;
17'h40e7:	data_out=16'h9af;
17'h40e8:	data_out=16'h9ff;
17'h40e9:	data_out=16'h8a00;
17'h40ea:	data_out=16'h968;
17'h40eb:	data_out=16'h9d7;
17'h40ec:	data_out=16'h89ff;
17'h40ed:	data_out=16'h89ff;
17'h40ee:	data_out=16'h96f;
17'h40ef:	data_out=16'ha00;
17'h40f0:	data_out=16'h9ba;
17'h40f1:	data_out=16'h89de;
17'h40f2:	data_out=16'h9f7;
17'h40f3:	data_out=16'ha00;
17'h40f4:	data_out=16'ha00;
17'h40f5:	data_out=16'ha00;
17'h40f6:	data_out=16'h853;
17'h40f7:	data_out=16'h89fd;
17'h40f8:	data_out=16'ha00;
17'h40f9:	data_out=16'h8a00;
17'h40fa:	data_out=16'h89ff;
17'h40fb:	data_out=16'h9ff;
17'h40fc:	data_out=16'h8a00;
17'h40fd:	data_out=16'h3e8;
17'h40fe:	data_out=16'h8a00;
17'h40ff:	data_out=16'h6bd;
17'h4100:	data_out=16'h89fa;
17'h4101:	data_out=16'h5ca;
17'h4102:	data_out=16'h8761;
17'h4103:	data_out=16'h8a00;
17'h4104:	data_out=16'h9fe;
17'h4105:	data_out=16'ha00;
17'h4106:	data_out=16'h7ea;
17'h4107:	data_out=16'h9e2;
17'h4108:	data_out=16'h89bf;
17'h4109:	data_out=16'h89fe;
17'h410a:	data_out=16'ha00;
17'h410b:	data_out=16'h89ff;
17'h410c:	data_out=16'h748;
17'h410d:	data_out=16'h8a00;
17'h410e:	data_out=16'h9ff;
17'h410f:	data_out=16'h89c7;
17'h4110:	data_out=16'h89fd;
17'h4111:	data_out=16'ha00;
17'h4112:	data_out=16'h8a00;
17'h4113:	data_out=16'h89d3;
17'h4114:	data_out=16'h89fe;
17'h4115:	data_out=16'h89e1;
17'h4116:	data_out=16'h89f5;
17'h4117:	data_out=16'h89fe;
17'h4118:	data_out=16'h8a00;
17'h4119:	data_out=16'ha00;
17'h411a:	data_out=16'ha00;
17'h411b:	data_out=16'h89e8;
17'h411c:	data_out=16'h86f2;
17'h411d:	data_out=16'h69b;
17'h411e:	data_out=16'h89fe;
17'h411f:	data_out=16'h89fc;
17'h4120:	data_out=16'h8994;
17'h4121:	data_out=16'h9ff;
17'h4122:	data_out=16'h45b;
17'h4123:	data_out=16'ha00;
17'h4124:	data_out=16'ha00;
17'h4125:	data_out=16'h3a8;
17'h4126:	data_out=16'h89e4;
17'h4127:	data_out=16'h5d5;
17'h4128:	data_out=16'ha00;
17'h4129:	data_out=16'h89e8;
17'h412a:	data_out=16'h89b1;
17'h412b:	data_out=16'h89e9;
17'h412c:	data_out=16'h89fe;
17'h412d:	data_out=16'h89ff;
17'h412e:	data_out=16'h89e3;
17'h412f:	data_out=16'h8831;
17'h4130:	data_out=16'ha00;
17'h4131:	data_out=16'ha00;
17'h4132:	data_out=16'ha00;
17'h4133:	data_out=16'h89ff;
17'h4134:	data_out=16'h89be;
17'h4135:	data_out=16'h9e2;
17'h4136:	data_out=16'h89bc;
17'h4137:	data_out=16'h8534;
17'h4138:	data_out=16'h80e2;
17'h4139:	data_out=16'h89ff;
17'h413a:	data_out=16'h89fd;
17'h413b:	data_out=16'ha00;
17'h413c:	data_out=16'h80fb;
17'h413d:	data_out=16'h89df;
17'h413e:	data_out=16'ha00;
17'h413f:	data_out=16'ha00;
17'h4140:	data_out=16'ha00;
17'h4141:	data_out=16'h89f3;
17'h4142:	data_out=16'h8a00;
17'h4143:	data_out=16'h9f8;
17'h4144:	data_out=16'ha00;
17'h4145:	data_out=16'h89e3;
17'h4146:	data_out=16'h89c0;
17'h4147:	data_out=16'h8a00;
17'h4148:	data_out=16'h450;
17'h4149:	data_out=16'h39b;
17'h414a:	data_out=16'h9fb;
17'h414b:	data_out=16'h8a00;
17'h414c:	data_out=16'h9eb;
17'h414d:	data_out=16'h940;
17'h414e:	data_out=16'h89fe;
17'h414f:	data_out=16'h812b;
17'h4150:	data_out=16'h84a2;
17'h4151:	data_out=16'h89ff;
17'h4152:	data_out=16'ha00;
17'h4153:	data_out=16'h7da;
17'h4154:	data_out=16'h89bb;
17'h4155:	data_out=16'h89f5;
17'h4156:	data_out=16'h860f;
17'h4157:	data_out=16'h89aa;
17'h4158:	data_out=16'h89ea;
17'h4159:	data_out=16'ha00;
17'h415a:	data_out=16'h89ff;
17'h415b:	data_out=16'h9f5;
17'h415c:	data_out=16'h87c1;
17'h415d:	data_out=16'h8701;
17'h415e:	data_out=16'h8671;
17'h415f:	data_out=16'h89ff;
17'h4160:	data_out=16'h89ec;
17'h4161:	data_out=16'ha00;
17'h4162:	data_out=16'h89fe;
17'h4163:	data_out=16'h89fe;
17'h4164:	data_out=16'h89fc;
17'h4165:	data_out=16'ha00;
17'h4166:	data_out=16'ha00;
17'h4167:	data_out=16'h89cb;
17'h4168:	data_out=16'ha00;
17'h4169:	data_out=16'h8a00;
17'h416a:	data_out=16'h9ff;
17'h416b:	data_out=16'h9f0;
17'h416c:	data_out=16'h89fa;
17'h416d:	data_out=16'h89fe;
17'h416e:	data_out=16'h9ff;
17'h416f:	data_out=16'ha00;
17'h4170:	data_out=16'h9ff;
17'h4171:	data_out=16'h89c8;
17'h4172:	data_out=16'h9fe;
17'h4173:	data_out=16'ha00;
17'h4174:	data_out=16'ha00;
17'h4175:	data_out=16'ha00;
17'h4176:	data_out=16'h89ec;
17'h4177:	data_out=16'h894b;
17'h4178:	data_out=16'ha00;
17'h4179:	data_out=16'h8a00;
17'h417a:	data_out=16'h89fe;
17'h417b:	data_out=16'ha00;
17'h417c:	data_out=16'h89f4;
17'h417d:	data_out=16'h4e1;
17'h417e:	data_out=16'h8a00;
17'h417f:	data_out=16'h9df;
17'h4180:	data_out=16'h89fd;
17'h4181:	data_out=16'h83bf;
17'h4182:	data_out=16'h8981;
17'h4183:	data_out=16'h89fe;
17'h4184:	data_out=16'h98b;
17'h4185:	data_out=16'ha00;
17'h4186:	data_out=16'h852;
17'h4187:	data_out=16'h9f5;
17'h4188:	data_out=16'h89d8;
17'h4189:	data_out=16'h89ed;
17'h418a:	data_out=16'ha00;
17'h418b:	data_out=16'h8a00;
17'h418c:	data_out=16'h8aa;
17'h418d:	data_out=16'h89df;
17'h418e:	data_out=16'h30c;
17'h418f:	data_out=16'h89ad;
17'h4190:	data_out=16'h8a00;
17'h4191:	data_out=16'h9ee;
17'h4192:	data_out=16'h8a00;
17'h4193:	data_out=16'h89d3;
17'h4194:	data_out=16'h89fe;
17'h4195:	data_out=16'h89ad;
17'h4196:	data_out=16'h36d;
17'h4197:	data_out=16'h89f7;
17'h4198:	data_out=16'h89e8;
17'h4199:	data_out=16'h9fe;
17'h419a:	data_out=16'ha00;
17'h419b:	data_out=16'h89f3;
17'h419c:	data_out=16'h8556;
17'h419d:	data_out=16'h847c;
17'h419e:	data_out=16'h89fd;
17'h419f:	data_out=16'h89d5;
17'h41a0:	data_out=16'h89bb;
17'h41a1:	data_out=16'h333;
17'h41a2:	data_out=16'h86d2;
17'h41a3:	data_out=16'ha00;
17'h41a4:	data_out=16'ha00;
17'h41a5:	data_out=16'h824e;
17'h41a6:	data_out=16'h89dc;
17'h41a7:	data_out=16'h89f3;
17'h41a8:	data_out=16'h3a3;
17'h41a9:	data_out=16'h89f1;
17'h41aa:	data_out=16'h89b2;
17'h41ab:	data_out=16'h89f8;
17'h41ac:	data_out=16'h4ba;
17'h41ad:	data_out=16'h89ff;
17'h41ae:	data_out=16'h89e8;
17'h41af:	data_out=16'h89e1;
17'h41b0:	data_out=16'ha00;
17'h41b1:	data_out=16'ha00;
17'h41b2:	data_out=16'ha00;
17'h41b3:	data_out=16'h89ff;
17'h41b4:	data_out=16'h89df;
17'h41b5:	data_out=16'h88c7;
17'h41b6:	data_out=16'h89ce;
17'h41b7:	data_out=16'h8987;
17'h41b8:	data_out=16'h8711;
17'h41b9:	data_out=16'h8a00;
17'h41ba:	data_out=16'h89fe;
17'h41bb:	data_out=16'ha00;
17'h41bc:	data_out=16'h89cc;
17'h41bd:	data_out=16'h89c4;
17'h41be:	data_out=16'h3ac;
17'h41bf:	data_out=16'ha00;
17'h41c0:	data_out=16'ha00;
17'h41c1:	data_out=16'h8a00;
17'h41c2:	data_out=16'h89f6;
17'h41c3:	data_out=16'h9fe;
17'h41c4:	data_out=16'ha00;
17'h41c5:	data_out=16'h89ad;
17'h41c6:	data_out=16'h8a00;
17'h41c7:	data_out=16'h8a00;
17'h41c8:	data_out=16'h8654;
17'h41c9:	data_out=16'h8176;
17'h41ca:	data_out=16'h9ee;
17'h41cb:	data_out=16'h8a00;
17'h41cc:	data_out=16'h9fc;
17'h41cd:	data_out=16'h84a3;
17'h41ce:	data_out=16'h8a00;
17'h41cf:	data_out=16'h80a1;
17'h41d0:	data_out=16'h1ee;
17'h41d1:	data_out=16'h89b9;
17'h41d2:	data_out=16'ha00;
17'h41d3:	data_out=16'h89da;
17'h41d4:	data_out=16'h89e9;
17'h41d5:	data_out=16'h89c8;
17'h41d6:	data_out=16'h8881;
17'h41d7:	data_out=16'h8999;
17'h41d8:	data_out=16'h89dd;
17'h41d9:	data_out=16'ha00;
17'h41da:	data_out=16'h8a00;
17'h41db:	data_out=16'h727;
17'h41dc:	data_out=16'h89bd;
17'h41dd:	data_out=16'h8956;
17'h41de:	data_out=16'h89bc;
17'h41df:	data_out=16'h89ff;
17'h41e0:	data_out=16'h89d7;
17'h41e1:	data_out=16'ha00;
17'h41e2:	data_out=16'h89fe;
17'h41e3:	data_out=16'h89ff;
17'h41e4:	data_out=16'h8a00;
17'h41e5:	data_out=16'ha00;
17'h41e6:	data_out=16'ha00;
17'h41e7:	data_out=16'h89f3;
17'h41e8:	data_out=16'h32f;
17'h41e9:	data_out=16'h8a00;
17'h41ea:	data_out=16'h2dd;
17'h41eb:	data_out=16'h9fd;
17'h41ec:	data_out=16'h89f6;
17'h41ed:	data_out=16'h89ff;
17'h41ee:	data_out=16'h2e2;
17'h41ef:	data_out=16'ha00;
17'h41f0:	data_out=16'h305;
17'h41f1:	data_out=16'h8990;
17'h41f2:	data_out=16'ha00;
17'h41f3:	data_out=16'ha00;
17'h41f4:	data_out=16'ha00;
17'h41f5:	data_out=16'ha00;
17'h41f6:	data_out=16'h89ff;
17'h41f7:	data_out=16'h89ea;
17'h41f8:	data_out=16'ha00;
17'h41f9:	data_out=16'h8a00;
17'h41fa:	data_out=16'h89ff;
17'h41fb:	data_out=16'h3b3;
17'h41fc:	data_out=16'h89e1;
17'h41fd:	data_out=16'h651;
17'h41fe:	data_out=16'h8a00;
17'h41ff:	data_out=16'h9e5;
17'h4200:	data_out=16'h89fc;
17'h4201:	data_out=16'h89fa;
17'h4202:	data_out=16'h89da;
17'h4203:	data_out=16'h89ff;
17'h4204:	data_out=16'h567;
17'h4205:	data_out=16'ha00;
17'h4206:	data_out=16'h86c;
17'h4207:	data_out=16'h9f8;
17'h4208:	data_out=16'h8a00;
17'h4209:	data_out=16'h89fc;
17'h420a:	data_out=16'h9f0;
17'h420b:	data_out=16'h8a00;
17'h420c:	data_out=16'h589;
17'h420d:	data_out=16'h891d;
17'h420e:	data_out=16'h812f;
17'h420f:	data_out=16'h89f6;
17'h4210:	data_out=16'h8a00;
17'h4211:	data_out=16'h3c8;
17'h4212:	data_out=16'h8a00;
17'h4213:	data_out=16'h87fb;
17'h4214:	data_out=16'h8a00;
17'h4215:	data_out=16'h82ab;
17'h4216:	data_out=16'h79e;
17'h4217:	data_out=16'h89ff;
17'h4218:	data_out=16'h89d9;
17'h4219:	data_out=16'h9a4;
17'h421a:	data_out=16'h9f5;
17'h421b:	data_out=16'h8a00;
17'h421c:	data_out=16'h8a00;
17'h421d:	data_out=16'h89ff;
17'h421e:	data_out=16'h89ff;
17'h421f:	data_out=16'h89f7;
17'h4220:	data_out=16'h89f8;
17'h4221:	data_out=16'h8130;
17'h4222:	data_out=16'h8a00;
17'h4223:	data_out=16'ha00;
17'h4224:	data_out=16'ha00;
17'h4225:	data_out=16'h8480;
17'h4226:	data_out=16'h8a00;
17'h4227:	data_out=16'h89fc;
17'h4228:	data_out=16'h818c;
17'h4229:	data_out=16'h8a00;
17'h422a:	data_out=16'h89ff;
17'h422b:	data_out=16'h89fc;
17'h422c:	data_out=16'h822;
17'h422d:	data_out=16'h8a00;
17'h422e:	data_out=16'h8a00;
17'h422f:	data_out=16'h89ff;
17'h4230:	data_out=16'h9ff;
17'h4231:	data_out=16'ha00;
17'h4232:	data_out=16'h9f8;
17'h4233:	data_out=16'h8a00;
17'h4234:	data_out=16'h89f1;
17'h4235:	data_out=16'h89fb;
17'h4236:	data_out=16'h8a00;
17'h4237:	data_out=16'h89e8;
17'h4238:	data_out=16'h8a00;
17'h4239:	data_out=16'h8a00;
17'h423a:	data_out=16'h89f2;
17'h423b:	data_out=16'h8fa;
17'h423c:	data_out=16'h89ff;
17'h423d:	data_out=16'h89d3;
17'h423e:	data_out=16'h818f;
17'h423f:	data_out=16'h9ff;
17'h4240:	data_out=16'h9fd;
17'h4241:	data_out=16'h8a00;
17'h4242:	data_out=16'h8a00;
17'h4243:	data_out=16'h9fe;
17'h4244:	data_out=16'h87cf;
17'h4245:	data_out=16'h8284;
17'h4246:	data_out=16'h8a00;
17'h4247:	data_out=16'h8a00;
17'h4248:	data_out=16'h8a00;
17'h4249:	data_out=16'h82c5;
17'h424a:	data_out=16'hab;
17'h424b:	data_out=16'h8a00;
17'h424c:	data_out=16'h9fa;
17'h424d:	data_out=16'h8816;
17'h424e:	data_out=16'h8a00;
17'h424f:	data_out=16'h6a8;
17'h4250:	data_out=16'h38d;
17'h4251:	data_out=16'h8918;
17'h4252:	data_out=16'h9f4;
17'h4253:	data_out=16'h8a00;
17'h4254:	data_out=16'h89fd;
17'h4255:	data_out=16'h89e2;
17'h4256:	data_out=16'h89ea;
17'h4257:	data_out=16'h89a3;
17'h4258:	data_out=16'h89fa;
17'h4259:	data_out=16'h9ef;
17'h425a:	data_out=16'h8a00;
17'h425b:	data_out=16'h89fa;
17'h425c:	data_out=16'h89f4;
17'h425d:	data_out=16'h89a6;
17'h425e:	data_out=16'h89e5;
17'h425f:	data_out=16'h8a00;
17'h4260:	data_out=16'h89fc;
17'h4261:	data_out=16'h9fa;
17'h4262:	data_out=16'h8a00;
17'h4263:	data_out=16'h8a00;
17'h4264:	data_out=16'h8a00;
17'h4265:	data_out=16'ha00;
17'h4266:	data_out=16'h9f6;
17'h4267:	data_out=16'h89fe;
17'h4268:	data_out=16'h8159;
17'h4269:	data_out=16'h8a00;
17'h426a:	data_out=16'h8132;
17'h426b:	data_out=16'h9f2;
17'h426c:	data_out=16'h89d5;
17'h426d:	data_out=16'h8a00;
17'h426e:	data_out=16'h8130;
17'h426f:	data_out=16'ha00;
17'h4270:	data_out=16'h812b;
17'h4271:	data_out=16'h89cb;
17'h4272:	data_out=16'h9f1;
17'h4273:	data_out=16'h9fc;
17'h4274:	data_out=16'ha00;
17'h4275:	data_out=16'ha00;
17'h4276:	data_out=16'h8a00;
17'h4277:	data_out=16'h8a00;
17'h4278:	data_out=16'h9f2;
17'h4279:	data_out=16'h8a00;
17'h427a:	data_out=16'h8a00;
17'h427b:	data_out=16'h818e;
17'h427c:	data_out=16'h89d5;
17'h427d:	data_out=16'h654;
17'h427e:	data_out=16'h8a00;
17'h427f:	data_out=16'h9f0;
17'h4280:	data_out=16'h2ef;
17'h4281:	data_out=16'h89e5;
17'h4282:	data_out=16'h884b;
17'h4283:	data_out=16'h89fe;
17'h4284:	data_out=16'h9c5;
17'h4285:	data_out=16'h9f5;
17'h4286:	data_out=16'h8968;
17'h4287:	data_out=16'h9ff;
17'h4288:	data_out=16'h89fe;
17'h4289:	data_out=16'h89ff;
17'h428a:	data_out=16'h9f9;
17'h428b:	data_out=16'h8a00;
17'h428c:	data_out=16'h94d;
17'h428d:	data_out=16'h9c1;
17'h428e:	data_out=16'h6a3;
17'h428f:	data_out=16'h895c;
17'h4290:	data_out=16'h89fe;
17'h4291:	data_out=16'h8141;
17'h4292:	data_out=16'h89f1;
17'h4293:	data_out=16'h8455;
17'h4294:	data_out=16'h8a00;
17'h4295:	data_out=16'h9f6;
17'h4296:	data_out=16'h9ed;
17'h4297:	data_out=16'h89ff;
17'h4298:	data_out=16'h9fa;
17'h4299:	data_out=16'h9e6;
17'h429a:	data_out=16'h9ee;
17'h429b:	data_out=16'h8a00;
17'h429c:	data_out=16'h89ff;
17'h429d:	data_out=16'h8a00;
17'h429e:	data_out=16'h89fd;
17'h429f:	data_out=16'h87f4;
17'h42a0:	data_out=16'h89da;
17'h42a1:	data_out=16'h641;
17'h42a2:	data_out=16'h89ff;
17'h42a3:	data_out=16'ha00;
17'h42a4:	data_out=16'ha00;
17'h42a5:	data_out=16'h85ac;
17'h42a6:	data_out=16'h89ff;
17'h42a7:	data_out=16'h89fe;
17'h42a8:	data_out=16'h522;
17'h42a9:	data_out=16'h89f7;
17'h42aa:	data_out=16'h89f1;
17'h42ab:	data_out=16'h8a00;
17'h42ac:	data_out=16'h9eb;
17'h42ad:	data_out=16'h8a00;
17'h42ae:	data_out=16'h8a00;
17'h42af:	data_out=16'h89fe;
17'h42b0:	data_out=16'ha00;
17'h42b1:	data_out=16'h8347;
17'h42b2:	data_out=16'h9f1;
17'h42b3:	data_out=16'h8a00;
17'h42b4:	data_out=16'h89f3;
17'h42b5:	data_out=16'h89fc;
17'h42b6:	data_out=16'h89fd;
17'h42b7:	data_out=16'h899e;
17'h42b8:	data_out=16'h89ff;
17'h42b9:	data_out=16'h8a00;
17'h42ba:	data_out=16'h89fe;
17'h42bb:	data_out=16'h88b;
17'h42bc:	data_out=16'h89ff;
17'h42bd:	data_out=16'h8544;
17'h42be:	data_out=16'h519;
17'h42bf:	data_out=16'h9f5;
17'h42c0:	data_out=16'h9ec;
17'h42c1:	data_out=16'h89ff;
17'h42c2:	data_out=16'h8a00;
17'h42c3:	data_out=16'h9f7;
17'h42c4:	data_out=16'h833f;
17'h42c5:	data_out=16'h9f6;
17'h42c6:	data_out=16'h8a00;
17'h42c7:	data_out=16'h8a00;
17'h42c8:	data_out=16'h8a00;
17'h42c9:	data_out=16'h8379;
17'h42ca:	data_out=16'h778;
17'h42cb:	data_out=16'h8a00;
17'h42cc:	data_out=16'h9f3;
17'h42cd:	data_out=16'h89fe;
17'h42ce:	data_out=16'h8a00;
17'h42cf:	data_out=16'h997;
17'h42d0:	data_out=16'h6ba;
17'h42d1:	data_out=16'h5d6;
17'h42d2:	data_out=16'h9fe;
17'h42d3:	data_out=16'h8a00;
17'h42d4:	data_out=16'h89fc;
17'h42d5:	data_out=16'h89fa;
17'h42d6:	data_out=16'h7d3;
17'h42d7:	data_out=16'h858a;
17'h42d8:	data_out=16'h8035;
17'h42d9:	data_out=16'h9ec;
17'h42da:	data_out=16'h8a00;
17'h42db:	data_out=16'h812d;
17'h42dc:	data_out=16'h8a00;
17'h42dd:	data_out=16'h142;
17'h42de:	data_out=16'h89de;
17'h42df:	data_out=16'h824d;
17'h42e0:	data_out=16'h89ff;
17'h42e1:	data_out=16'h9fb;
17'h42e2:	data_out=16'h8a00;
17'h42e3:	data_out=16'h8a00;
17'h42e4:	data_out=16'h8a00;
17'h42e5:	data_out=16'ha00;
17'h42e6:	data_out=16'h9e7;
17'h42e7:	data_out=16'h89fe;
17'h42e8:	data_out=16'h5d5;
17'h42e9:	data_out=16'h8a00;
17'h42ea:	data_out=16'h6e8;
17'h42eb:	data_out=16'h9e7;
17'h42ec:	data_out=16'h9f1;
17'h42ed:	data_out=16'h8a00;
17'h42ee:	data_out=16'h6e9;
17'h42ef:	data_out=16'h9ee;
17'h42f0:	data_out=16'h6c6;
17'h42f1:	data_out=16'h2ab;
17'h42f2:	data_out=16'h9eb;
17'h42f3:	data_out=16'h9f0;
17'h42f4:	data_out=16'ha00;
17'h42f5:	data_out=16'h791;
17'h42f6:	data_out=16'h8a00;
17'h42f7:	data_out=16'h89fe;
17'h42f8:	data_out=16'h9e5;
17'h42f9:	data_out=16'h895a;
17'h42fa:	data_out=16'h8a00;
17'h42fb:	data_out=16'h518;
17'h42fc:	data_out=16'h9fc;
17'h42fd:	data_out=16'h848f;
17'h42fe:	data_out=16'h8a00;
17'h42ff:	data_out=16'h9f1;
17'h4300:	data_out=16'h1bf;
17'h4301:	data_out=16'h89ff;
17'h4302:	data_out=16'h8321;
17'h4303:	data_out=16'h89ff;
17'h4304:	data_out=16'h9d0;
17'h4305:	data_out=16'h413;
17'h4306:	data_out=16'h850c;
17'h4307:	data_out=16'ha00;
17'h4308:	data_out=16'h83c6;
17'h4309:	data_out=16'h899a;
17'h430a:	data_out=16'h82cb;
17'h430b:	data_out=16'h8a00;
17'h430c:	data_out=16'h9f2;
17'h430d:	data_out=16'h9f1;
17'h430e:	data_out=16'h7b6;
17'h430f:	data_out=16'h6ee;
17'h4310:	data_out=16'h89ff;
17'h4311:	data_out=16'h8a00;
17'h4312:	data_out=16'h8973;
17'h4313:	data_out=16'h878c;
17'h4314:	data_out=16'h8a00;
17'h4315:	data_out=16'h9f6;
17'h4316:	data_out=16'h9e8;
17'h4317:	data_out=16'h8a00;
17'h4318:	data_out=16'h9fb;
17'h4319:	data_out=16'h9e7;
17'h431a:	data_out=16'h9e4;
17'h431b:	data_out=16'h8a00;
17'h431c:	data_out=16'h89ff;
17'h431d:	data_out=16'h8a00;
17'h431e:	data_out=16'h89fe;
17'h431f:	data_out=16'h817c;
17'h4320:	data_out=16'h89ff;
17'h4321:	data_out=16'h75e;
17'h4322:	data_out=16'h89ff;
17'h4323:	data_out=16'ha00;
17'h4324:	data_out=16'ha00;
17'h4325:	data_out=16'h38d;
17'h4326:	data_out=16'h8253;
17'h4327:	data_out=16'h8a00;
17'h4328:	data_out=16'h65f;
17'h4329:	data_out=16'h89f4;
17'h432a:	data_out=16'h8447;
17'h432b:	data_out=16'h8a00;
17'h432c:	data_out=16'h9e8;
17'h432d:	data_out=16'h89ff;
17'h432e:	data_out=16'h89ff;
17'h432f:	data_out=16'h89ff;
17'h4330:	data_out=16'ha00;
17'h4331:	data_out=16'h89d6;
17'h4332:	data_out=16'h9e8;
17'h4333:	data_out=16'h8a00;
17'h4334:	data_out=16'h89f7;
17'h4335:	data_out=16'h877f;
17'h4336:	data_out=16'h89c7;
17'h4337:	data_out=16'h890b;
17'h4338:	data_out=16'h8a00;
17'h4339:	data_out=16'h8a00;
17'h433a:	data_out=16'h88ef;
17'h433b:	data_out=16'h5de;
17'h433c:	data_out=16'h8a00;
17'h433d:	data_out=16'h8981;
17'h433e:	data_out=16'h657;
17'h433f:	data_out=16'h44c;
17'h4340:	data_out=16'h9e5;
17'h4341:	data_out=16'h89f9;
17'h4342:	data_out=16'h53d;
17'h4343:	data_out=16'h611;
17'h4344:	data_out=16'h89d1;
17'h4345:	data_out=16'h9f5;
17'h4346:	data_out=16'h8a00;
17'h4347:	data_out=16'h95;
17'h4348:	data_out=16'h89ff;
17'h4349:	data_out=16'h440;
17'h434a:	data_out=16'h84c;
17'h434b:	data_out=16'h8166;
17'h434c:	data_out=16'h9fb;
17'h434d:	data_out=16'h89ff;
17'h434e:	data_out=16'h8a00;
17'h434f:	data_out=16'h9f8;
17'h4350:	data_out=16'h558;
17'h4351:	data_out=16'h9ed;
17'h4352:	data_out=16'ha00;
17'h4353:	data_out=16'h8a00;
17'h4354:	data_out=16'h8a00;
17'h4355:	data_out=16'h898a;
17'h4356:	data_out=16'h722;
17'h4357:	data_out=16'h8491;
17'h4358:	data_out=16'h482;
17'h4359:	data_out=16'h9e5;
17'h435a:	data_out=16'h8a00;
17'h435b:	data_out=16'h89ff;
17'h435c:	data_out=16'h8a00;
17'h435d:	data_out=16'h251;
17'h435e:	data_out=16'h89fe;
17'h435f:	data_out=16'h65b;
17'h4360:	data_out=16'h89ec;
17'h4361:	data_out=16'h87f1;
17'h4362:	data_out=16'h8a00;
17'h4363:	data_out=16'h8a00;
17'h4364:	data_out=16'h8a00;
17'h4365:	data_out=16'h9fa;
17'h4366:	data_out=16'h96a;
17'h4367:	data_out=16'h8a00;
17'h4368:	data_out=16'h702;
17'h4369:	data_out=16'h85e1;
17'h436a:	data_out=16'h7f1;
17'h436b:	data_out=16'h884;
17'h436c:	data_out=16'h9ed;
17'h436d:	data_out=16'h8a00;
17'h436e:	data_out=16'h7f2;
17'h436f:	data_out=16'h948;
17'h4370:	data_out=16'h7d4;
17'h4371:	data_out=16'h9e0;
17'h4372:	data_out=16'h89bc;
17'h4373:	data_out=16'h891e;
17'h4374:	data_out=16'ha00;
17'h4375:	data_out=16'h89c1;
17'h4376:	data_out=16'h8a00;
17'h4377:	data_out=16'h75b;
17'h4378:	data_out=16'h276;
17'h4379:	data_out=16'h48e;
17'h437a:	data_out=16'h8a00;
17'h437b:	data_out=16'h656;
17'h437c:	data_out=16'h9fc;
17'h437d:	data_out=16'h85ab;
17'h437e:	data_out=16'h8a00;
17'h437f:	data_out=16'h9e7;
17'h4380:	data_out=16'h8150;
17'h4381:	data_out=16'h8a00;
17'h4382:	data_out=16'h9f8;
17'h4383:	data_out=16'h89af;
17'h4384:	data_out=16'h80d;
17'h4385:	data_out=16'h84b8;
17'h4386:	data_out=16'h3cd;
17'h4387:	data_out=16'ha00;
17'h4388:	data_out=16'h940;
17'h4389:	data_out=16'h9f0;
17'h438a:	data_out=16'h89fb;
17'h438b:	data_out=16'h8a00;
17'h438c:	data_out=16'ha00;
17'h438d:	data_out=16'ha00;
17'h438e:	data_out=16'h686;
17'h438f:	data_out=16'h9f7;
17'h4390:	data_out=16'h224;
17'h4391:	data_out=16'h8815;
17'h4392:	data_out=16'h87c6;
17'h4393:	data_out=16'h814d;
17'h4394:	data_out=16'h8a00;
17'h4395:	data_out=16'ha00;
17'h4396:	data_out=16'h9ff;
17'h4397:	data_out=16'h8a00;
17'h4398:	data_out=16'ha00;
17'h4399:	data_out=16'h72f;
17'h439a:	data_out=16'h903;
17'h439b:	data_out=16'h8a00;
17'h439c:	data_out=16'h8a00;
17'h439d:	data_out=16'h8a00;
17'h439e:	data_out=16'h89dd;
17'h439f:	data_out=16'h690;
17'h43a0:	data_out=16'h8a00;
17'h43a1:	data_out=16'h64a;
17'h43a2:	data_out=16'h85eb;
17'h43a3:	data_out=16'ha00;
17'h43a4:	data_out=16'ha00;
17'h43a5:	data_out=16'ha00;
17'h43a6:	data_out=16'h769;
17'h43a7:	data_out=16'h8a00;
17'h43a8:	data_out=16'h592;
17'h43a9:	data_out=16'h8a00;
17'h43aa:	data_out=16'h9f6;
17'h43ab:	data_out=16'h8a00;
17'h43ac:	data_out=16'h9fe;
17'h43ad:	data_out=16'h8a00;
17'h43ae:	data_out=16'h516;
17'h43af:	data_out=16'h8a00;
17'h43b0:	data_out=16'h4e4;
17'h43b1:	data_out=16'h89f7;
17'h43b2:	data_out=16'h38c;
17'h43b3:	data_out=16'h8a00;
17'h43b4:	data_out=16'h89fb;
17'h43b5:	data_out=16'h2b2;
17'h43b6:	data_out=16'h8dc;
17'h43b7:	data_out=16'h847;
17'h43b8:	data_out=16'h8a00;
17'h43b9:	data_out=16'h8a00;
17'h43ba:	data_out=16'ha00;
17'h43bb:	data_out=16'h4d9;
17'h43bc:	data_out=16'h8a00;
17'h43bd:	data_out=16'h82f7;
17'h43be:	data_out=16'h58b;
17'h43bf:	data_out=16'h848f;
17'h43c0:	data_out=16'h9e1;
17'h43c1:	data_out=16'h82c8;
17'h43c2:	data_out=16'ha00;
17'h43c3:	data_out=16'h42;
17'h43c4:	data_out=16'h8933;
17'h43c5:	data_out=16'ha00;
17'h43c6:	data_out=16'h8a00;
17'h43c7:	data_out=16'ha00;
17'h43c8:	data_out=16'h88d2;
17'h43c9:	data_out=16'h9ff;
17'h43ca:	data_out=16'h84a;
17'h43cb:	data_out=16'h9ef;
17'h43cc:	data_out=16'ha00;
17'h43cd:	data_out=16'h8781;
17'h43ce:	data_out=16'h8c0;
17'h43cf:	data_out=16'ha00;
17'h43d0:	data_out=16'h811;
17'h43d1:	data_out=16'h9f7;
17'h43d2:	data_out=16'ha00;
17'h43d3:	data_out=16'h8a00;
17'h43d4:	data_out=16'h8a00;
17'h43d5:	data_out=16'h7d1;
17'h43d6:	data_out=16'h9ff;
17'h43d7:	data_out=16'h9f8;
17'h43d8:	data_out=16'h99a;
17'h43d9:	data_out=16'h9ed;
17'h43da:	data_out=16'h8a00;
17'h43db:	data_out=16'h8a00;
17'h43dc:	data_out=16'h8a00;
17'h43dd:	data_out=16'h9ef;
17'h43de:	data_out=16'h8a00;
17'h43df:	data_out=16'h9ec;
17'h43e0:	data_out=16'h258;
17'h43e1:	data_out=16'h8a00;
17'h43e2:	data_out=16'h8a00;
17'h43e3:	data_out=16'h8a00;
17'h43e4:	data_out=16'h8a00;
17'h43e5:	data_out=16'ha00;
17'h43e6:	data_out=16'h705;
17'h43e7:	data_out=16'h8a00;
17'h43e8:	data_out=16'h60b;
17'h43e9:	data_out=16'h9fe;
17'h43ea:	data_out=16'h6b1;
17'h43eb:	data_out=16'h893;
17'h43ec:	data_out=16'h9ff;
17'h43ed:	data_out=16'h8a00;
17'h43ee:	data_out=16'h6b1;
17'h43ef:	data_out=16'h1b9;
17'h43f0:	data_out=16'h69a;
17'h43f1:	data_out=16'h9f8;
17'h43f2:	data_out=16'h8a00;
17'h43f3:	data_out=16'h86f5;
17'h43f4:	data_out=16'h58d;
17'h43f5:	data_out=16'h8a00;
17'h43f6:	data_out=16'h8a00;
17'h43f7:	data_out=16'h9f7;
17'h43f8:	data_out=16'h8285;
17'h43f9:	data_out=16'h9fa;
17'h43fa:	data_out=16'h8a00;
17'h43fb:	data_out=16'h58a;
17'h43fc:	data_out=16'h9ff;
17'h43fd:	data_out=16'h80a9;
17'h43fe:	data_out=16'h854f;
17'h43ff:	data_out=16'h9f0;
17'h4400:	data_out=16'h89fb;
17'h4401:	data_out=16'h8a00;
17'h4402:	data_out=16'h9fc;
17'h4403:	data_out=16'h8a00;
17'h4404:	data_out=16'h302;
17'h4405:	data_out=16'h8294;
17'h4406:	data_out=16'h14a;
17'h4407:	data_out=16'ha00;
17'h4408:	data_out=16'h995;
17'h4409:	data_out=16'h8b8;
17'h440a:	data_out=16'h89ff;
17'h440b:	data_out=16'h8a00;
17'h440c:	data_out=16'h9fe;
17'h440d:	data_out=16'h3bc;
17'h440e:	data_out=16'h63e;
17'h440f:	data_out=16'h9f9;
17'h4410:	data_out=16'h83d7;
17'h4411:	data_out=16'h8957;
17'h4412:	data_out=16'h82e3;
17'h4413:	data_out=16'h87f5;
17'h4414:	data_out=16'h8a00;
17'h4415:	data_out=16'h7e9;
17'h4416:	data_out=16'h6fc;
17'h4417:	data_out=16'h8a00;
17'h4418:	data_out=16'h9ff;
17'h4419:	data_out=16'h4aa;
17'h441a:	data_out=16'h2a9;
17'h441b:	data_out=16'h89fe;
17'h441c:	data_out=16'h8a00;
17'h441d:	data_out=16'h8a00;
17'h441e:	data_out=16'h89c3;
17'h441f:	data_out=16'h9eb;
17'h4420:	data_out=16'h8a00;
17'h4421:	data_out=16'h619;
17'h4422:	data_out=16'h86f8;
17'h4423:	data_out=16'ha00;
17'h4424:	data_out=16'ha00;
17'h4425:	data_out=16'ha00;
17'h4426:	data_out=16'h83f5;
17'h4427:	data_out=16'h8a00;
17'h4428:	data_out=16'h5b9;
17'h4429:	data_out=16'h882a;
17'h442a:	data_out=16'h9f7;
17'h442b:	data_out=16'h8a00;
17'h442c:	data_out=16'h60b;
17'h442d:	data_out=16'h8a00;
17'h442e:	data_out=16'h9eb;
17'h442f:	data_out=16'h8a00;
17'h4430:	data_out=16'h81cb;
17'h4431:	data_out=16'h8a00;
17'h4432:	data_out=16'h82d6;
17'h4433:	data_out=16'h8a00;
17'h4434:	data_out=16'h8a00;
17'h4435:	data_out=16'h406;
17'h4436:	data_out=16'h7f7;
17'h4437:	data_out=16'h9fa;
17'h4438:	data_out=16'h8a00;
17'h4439:	data_out=16'h8a00;
17'h443a:	data_out=16'h653;
17'h443b:	data_out=16'h8547;
17'h443c:	data_out=16'h8a00;
17'h443d:	data_out=16'h878c;
17'h443e:	data_out=16'h5b5;
17'h443f:	data_out=16'h8282;
17'h4440:	data_out=16'h932;
17'h4441:	data_out=16'h4a7;
17'h4442:	data_out=16'h92b;
17'h4443:	data_out=16'h114;
17'h4444:	data_out=16'h8a00;
17'h4445:	data_out=16'h7fa;
17'h4446:	data_out=16'h8a00;
17'h4447:	data_out=16'h8bd;
17'h4448:	data_out=16'h20f;
17'h4449:	data_out=16'h9ab;
17'h444a:	data_out=16'h86f;
17'h444b:	data_out=16'h79e;
17'h444c:	data_out=16'ha00;
17'h444d:	data_out=16'h87ef;
17'h444e:	data_out=16'h9ef;
17'h444f:	data_out=16'ha00;
17'h4450:	data_out=16'h82c;
17'h4451:	data_out=16'h9f7;
17'h4452:	data_out=16'ha00;
17'h4453:	data_out=16'h8a00;
17'h4454:	data_out=16'h8a00;
17'h4455:	data_out=16'h9ac;
17'h4456:	data_out=16'h9f9;
17'h4457:	data_out=16'h9fb;
17'h4458:	data_out=16'h9f5;
17'h4459:	data_out=16'h9da;
17'h445a:	data_out=16'h8a00;
17'h445b:	data_out=16'h88e8;
17'h445c:	data_out=16'h8a00;
17'h445d:	data_out=16'h4f5;
17'h445e:	data_out=16'h8a00;
17'h445f:	data_out=16'h6d2;
17'h4460:	data_out=16'h894c;
17'h4461:	data_out=16'h89fc;
17'h4462:	data_out=16'h8a00;
17'h4463:	data_out=16'h8a00;
17'h4464:	data_out=16'h8a00;
17'h4465:	data_out=16'hb2;
17'h4466:	data_out=16'h49;
17'h4467:	data_out=16'h8a00;
17'h4468:	data_out=16'h5f5;
17'h4469:	data_out=16'h9cb;
17'h446a:	data_out=16'h660;
17'h446b:	data_out=16'h802c;
17'h446c:	data_out=16'h86d8;
17'h446d:	data_out=16'h8a00;
17'h446e:	data_out=16'h660;
17'h446f:	data_out=16'h89ff;
17'h4470:	data_out=16'h64e;
17'h4471:	data_out=16'h9f8;
17'h4472:	data_out=16'h8927;
17'h4473:	data_out=16'h84d4;
17'h4474:	data_out=16'h8164;
17'h4475:	data_out=16'h8a00;
17'h4476:	data_out=16'h8a00;
17'h4477:	data_out=16'ha00;
17'h4478:	data_out=16'h8222;
17'h4479:	data_out=16'h9fc;
17'h447a:	data_out=16'h8a00;
17'h447b:	data_out=16'h5b5;
17'h447c:	data_out=16'h9ff;
17'h447d:	data_out=16'h373;
17'h447e:	data_out=16'h87ce;
17'h447f:	data_out=16'h9ff;
17'h4480:	data_out=16'h8a00;
17'h4481:	data_out=16'h88d7;
17'h4482:	data_out=16'h3be;
17'h4483:	data_out=16'h86b0;
17'h4484:	data_out=16'h2d8;
17'h4485:	data_out=16'h80ec;
17'h4486:	data_out=16'hd5;
17'h4487:	data_out=16'h30d;
17'h4488:	data_out=16'h82a4;
17'h4489:	data_out=16'h8092;
17'h448a:	data_out=16'h8798;
17'h448b:	data_out=16'h8a00;
17'h448c:	data_out=16'h4e1;
17'h448d:	data_out=16'h83e8;
17'h448e:	data_out=16'h1b0;
17'h448f:	data_out=16'h2cd;
17'h4490:	data_out=16'h83ad;
17'h4491:	data_out=16'h8167;
17'h4492:	data_out=16'h82bd;
17'h4493:	data_out=16'h84d0;
17'h4494:	data_out=16'h8769;
17'h4495:	data_out=16'h80af;
17'h4496:	data_out=16'h840b;
17'h4497:	data_out=16'h89a4;
17'h4498:	data_out=16'h359;
17'h4499:	data_out=16'h538;
17'h449a:	data_out=16'h299;
17'h449b:	data_out=16'h89fe;
17'h449c:	data_out=16'h863f;
17'h449d:	data_out=16'h8a00;
17'h449e:	data_out=16'h870a;
17'h449f:	data_out=16'h5da;
17'h44a0:	data_out=16'h8a00;
17'h44a1:	data_out=16'h19d;
17'h44a2:	data_out=16'h81c4;
17'h44a3:	data_out=16'h3a2;
17'h44a4:	data_out=16'h3a2;
17'h44a5:	data_out=16'h31e;
17'h44a6:	data_out=16'h88b2;
17'h44a7:	data_out=16'h8a00;
17'h44a8:	data_out=16'h189;
17'h44a9:	data_out=16'h85a4;
17'h44aa:	data_out=16'h81fa;
17'h44ab:	data_out=16'h8a00;
17'h44ac:	data_out=16'h83aa;
17'h44ad:	data_out=16'h893d;
17'h44ae:	data_out=16'h179;
17'h44af:	data_out=16'h89d6;
17'h44b0:	data_out=16'h43;
17'h44b1:	data_out=16'h8a00;
17'h44b2:	data_out=16'h37;
17'h44b3:	data_out=16'h86c8;
17'h44b4:	data_out=16'h8624;
17'h44b5:	data_out=16'h9a;
17'h44b6:	data_out=16'h838f;
17'h44b7:	data_out=16'h36e;
17'h44b8:	data_out=16'h826b;
17'h44b9:	data_out=16'h86b6;
17'h44ba:	data_out=16'h1d;
17'h44bb:	data_out=16'h84be;
17'h44bc:	data_out=16'h84c1;
17'h44bd:	data_out=16'h8591;
17'h44be:	data_out=16'h17b;
17'h44bf:	data_out=16'h8073;
17'h44c0:	data_out=16'h558;
17'h44c1:	data_out=16'h31;
17'h44c2:	data_out=16'h2d2;
17'h44c3:	data_out=16'h19e;
17'h44c4:	data_out=16'h8864;
17'h44c5:	data_out=16'h8014;
17'h44c6:	data_out=16'h86c1;
17'h44c7:	data_out=16'h5f;
17'h44c8:	data_out=16'h8d;
17'h44c9:	data_out=16'h2c0;
17'h44ca:	data_out=16'h538;
17'h44cb:	data_out=16'h25c;
17'h44cc:	data_out=16'h76f;
17'h44cd:	data_out=16'h81f0;
17'h44ce:	data_out=16'h8066;
17'h44cf:	data_out=16'h60d;
17'h44d0:	data_out=16'h426;
17'h44d1:	data_out=16'h80be;
17'h44d2:	data_out=16'h422;
17'h44d3:	data_out=16'h8a00;
17'h44d4:	data_out=16'h87db;
17'h44d5:	data_out=16'h8170;
17'h44d6:	data_out=16'h275;
17'h44d7:	data_out=16'h40a;
17'h44d8:	data_out=16'hbe;
17'h44d9:	data_out=16'h4da;
17'h44da:	data_out=16'h8a00;
17'h44db:	data_out=16'h82fa;
17'h44dc:	data_out=16'h88f9;
17'h44dd:	data_out=16'h8183;
17'h44de:	data_out=16'h8953;
17'h44df:	data_out=16'h218;
17'h44e0:	data_out=16'h86d5;
17'h44e1:	data_out=16'h85a5;
17'h44e2:	data_out=16'h8a00;
17'h44e3:	data_out=16'h86fd;
17'h44e4:	data_out=16'h897b;
17'h44e5:	data_out=16'h8150;
17'h44e6:	data_out=16'hb5;
17'h44e7:	data_out=16'h84e7;
17'h44e8:	data_out=16'h19c;
17'h44e9:	data_out=16'h82f4;
17'h44ea:	data_out=16'h1bb;
17'h44eb:	data_out=16'h8053;
17'h44ec:	data_out=16'h8a00;
17'h44ed:	data_out=16'h86f2;
17'h44ee:	data_out=16'h1c7;
17'h44ef:	data_out=16'h83bb;
17'h44f0:	data_out=16'h1af;
17'h44f1:	data_out=16'h675;
17'h44f2:	data_out=16'h821b;
17'h44f3:	data_out=16'h8184;
17'h44f4:	data_out=16'h64;
17'h44f5:	data_out=16'h8841;
17'h44f6:	data_out=16'h8a00;
17'h44f7:	data_out=16'h480;
17'h44f8:	data_out=16'hd7;
17'h44f9:	data_out=16'h24b;
17'h44fa:	data_out=16'h874a;
17'h44fb:	data_out=16'h182;
17'h44fc:	data_out=16'h354;
17'h44fd:	data_out=16'h198;
17'h44fe:	data_out=16'h842c;
17'h44ff:	data_out=16'h8c7;
17'h4500:	data_out=16'h82bf;
17'h4501:	data_out=16'h8081;
17'h4502:	data_out=16'h8051;
17'h4503:	data_out=16'h80b0;
17'h4504:	data_out=16'h8033;
17'h4505:	data_out=16'h803d;
17'h4506:	data_out=16'h10d;
17'h4507:	data_out=16'h804d;
17'h4508:	data_out=16'h8320;
17'h4509:	data_out=16'h822d;
17'h450a:	data_out=16'h809d;
17'h450b:	data_out=16'h81c0;
17'h450c:	data_out=16'h81b6;
17'h450d:	data_out=16'h8116;
17'h450e:	data_out=16'h80;
17'h450f:	data_out=16'h8064;
17'h4510:	data_out=16'h8169;
17'h4511:	data_out=16'h8090;
17'h4512:	data_out=16'h808a;
17'h4513:	data_out=16'h1b;
17'h4514:	data_out=16'h8142;
17'h4515:	data_out=16'h807c;
17'h4516:	data_out=16'h8171;
17'h4517:	data_out=16'h8100;
17'h4518:	data_out=16'h8024;
17'h4519:	data_out=16'h172;
17'h451a:	data_out=16'h27;
17'h451b:	data_out=16'h817b;
17'h451c:	data_out=16'h80b0;
17'h451d:	data_out=16'h8263;
17'h451e:	data_out=16'h817d;
17'h451f:	data_out=16'h80ab;
17'h4520:	data_out=16'h8309;
17'h4521:	data_out=16'h7b;
17'h4522:	data_out=16'h8076;
17'h4523:	data_out=16'hb5;
17'h4524:	data_out=16'hc0;
17'h4525:	data_out=16'h806f;
17'h4526:	data_out=16'h8267;
17'h4527:	data_out=16'h8335;
17'h4528:	data_out=16'h7b;
17'h4529:	data_out=16'h95;
17'h452a:	data_out=16'h8151;
17'h452b:	data_out=16'h8337;
17'h452c:	data_out=16'h817f;
17'h452d:	data_out=16'h11c;
17'h452e:	data_out=16'h80c5;
17'h452f:	data_out=16'h815f;
17'h4530:	data_out=16'h21;
17'h4531:	data_out=16'h81dc;
17'h4532:	data_out=16'h57;
17'h4533:	data_out=16'h819a;
17'h4534:	data_out=16'h8009;
17'h4535:	data_out=16'h81d4;
17'h4536:	data_out=16'h81a6;
17'h4537:	data_out=16'h8007;
17'h4538:	data_out=16'h265;
17'h4539:	data_out=16'h81b6;
17'h453a:	data_out=16'h804a;
17'h453b:	data_out=16'h82de;
17'h453c:	data_out=16'h80e0;
17'h453d:	data_out=16'h8254;
17'h453e:	data_out=16'h7c;
17'h453f:	data_out=16'h3b;
17'h4540:	data_out=16'h17b;
17'h4541:	data_out=16'h81b1;
17'h4542:	data_out=16'hb9;
17'h4543:	data_out=16'h171;
17'h4544:	data_out=16'h8262;
17'h4545:	data_out=16'h80a0;
17'h4546:	data_out=16'hd6;
17'h4547:	data_out=16'h32;
17'h4548:	data_out=16'h806f;
17'h4549:	data_out=16'h804e;
17'h454a:	data_out=16'h8025;
17'h454b:	data_out=16'h71;
17'h454c:	data_out=16'h1be;
17'h454d:	data_out=16'h8061;
17'h454e:	data_out=16'h80a4;
17'h454f:	data_out=16'h12e;
17'h4550:	data_out=16'hf1;
17'h4551:	data_out=16'h8139;
17'h4552:	data_out=16'hb1;
17'h4553:	data_out=16'h82c6;
17'h4554:	data_out=16'h816a;
17'h4555:	data_out=16'h8184;
17'h4556:	data_out=16'h8059;
17'h4557:	data_out=16'h11f;
17'h4558:	data_out=16'h81c0;
17'h4559:	data_out=16'h15e;
17'h455a:	data_out=16'h80b6;
17'h455b:	data_out=16'hcd;
17'h455c:	data_out=16'h8156;
17'h455d:	data_out=16'h80b6;
17'h455e:	data_out=16'h815d;
17'h455f:	data_out=16'h3f;
17'h4560:	data_out=16'h11;
17'h4561:	data_out=16'h8059;
17'h4562:	data_out=16'h8106;
17'h4563:	data_out=16'h8172;
17'h4564:	data_out=16'h80cb;
17'h4565:	data_out=16'h8030;
17'h4566:	data_out=16'h800f;
17'h4567:	data_out=16'h23;
17'h4568:	data_out=16'h78;
17'h4569:	data_out=16'h8264;
17'h456a:	data_out=16'h96;
17'h456b:	data_out=16'h8102;
17'h456c:	data_out=16'h8196;
17'h456d:	data_out=16'h819a;
17'h456e:	data_out=16'h8d;
17'h456f:	data_out=16'h802e;
17'h4570:	data_out=16'h82;
17'h4571:	data_out=16'h80ca;
17'h4572:	data_out=16'hbc;
17'h4573:	data_out=16'h99;
17'h4574:	data_out=16'h36;
17'h4575:	data_out=16'h120;
17'h4576:	data_out=16'h82cf;
17'h4577:	data_out=16'h8025;
17'h4578:	data_out=16'h156;
17'h4579:	data_out=16'h80da;
17'h457a:	data_out=16'h8183;
17'h457b:	data_out=16'h7b;
17'h457c:	data_out=16'h1e;
17'h457d:	data_out=16'h10a;
17'h457e:	data_out=16'h8174;
17'h457f:	data_out=16'ha;
17'h4580:	data_out=16'h813e;
17'h4581:	data_out=16'h810a;
17'h4582:	data_out=16'h813d;
17'h4583:	data_out=16'h80ba;
17'h4584:	data_out=16'h56;
17'h4585:	data_out=16'h802a;
17'h4586:	data_out=16'h8006;
17'h4587:	data_out=16'h35;
17'h4588:	data_out=16'h81ce;
17'h4589:	data_out=16'h8082;
17'h458a:	data_out=16'h8095;
17'h458b:	data_out=16'h80cd;
17'h458c:	data_out=16'h175;
17'h458d:	data_out=16'h80a3;
17'h458e:	data_out=16'h8025;
17'h458f:	data_out=16'h813a;
17'h4590:	data_out=16'h8088;
17'h4591:	data_out=16'h18;
17'h4592:	data_out=16'h80e7;
17'h4593:	data_out=16'h8045;
17'h4594:	data_out=16'h8177;
17'h4595:	data_out=16'h806a;
17'h4596:	data_out=16'h80cd;
17'h4597:	data_out=16'h814c;
17'h4598:	data_out=16'h8069;
17'h4599:	data_out=16'h1e1;
17'h459a:	data_out=16'hb4;
17'h459b:	data_out=16'h80ff;
17'h459c:	data_out=16'h80f0;
17'h459d:	data_out=16'h8148;
17'h459e:	data_out=16'h818d;
17'h459f:	data_out=16'h80d4;
17'h45a0:	data_out=16'h817a;
17'h45a1:	data_out=16'h8022;
17'h45a2:	data_out=16'h30;
17'h45a3:	data_out=16'h802a;
17'h45a4:	data_out=16'h801e;
17'h45a5:	data_out=16'ha2;
17'h45a6:	data_out=16'h817a;
17'h45a7:	data_out=16'h819a;
17'h45a8:	data_out=16'h8029;
17'h45a9:	data_out=16'h807e;
17'h45aa:	data_out=16'h8174;
17'h45ab:	data_out=16'h8146;
17'h45ac:	data_out=16'h80ba;
17'h45ad:	data_out=16'hb0;
17'h45ae:	data_out=16'h8150;
17'h45af:	data_out=16'h80db;
17'h45b0:	data_out=16'hb1;
17'h45b1:	data_out=16'h8050;
17'h45b2:	data_out=16'hb9;
17'h45b3:	data_out=16'h8186;
17'h45b4:	data_out=16'h8035;
17'h45b5:	data_out=16'h6f;
17'h45b6:	data_out=16'h81a7;
17'h45b7:	data_out=16'h8133;
17'h45b8:	data_out=16'h8014;
17'h45b9:	data_out=16'h8189;
17'h45ba:	data_out=16'h80a4;
17'h45bb:	data_out=16'h8084;
17'h45bc:	data_out=16'h8157;
17'h45bd:	data_out=16'h8141;
17'h45be:	data_out=16'h8023;
17'h45bf:	data_out=16'h4e;
17'h45c0:	data_out=16'h48;
17'h45c1:	data_out=16'h814b;
17'h45c2:	data_out=16'h1a4;
17'h45c3:	data_out=16'h36;
17'h45c4:	data_out=16'h80bb;
17'h45c5:	data_out=16'h80b4;
17'h45c6:	data_out=16'h80c5;
17'h45c7:	data_out=16'h8075;
17'h45c8:	data_out=16'h8097;
17'h45c9:	data_out=16'h9a;
17'h45ca:	data_out=16'ha8;
17'h45cb:	data_out=16'h1df;
17'h45cc:	data_out=16'h14d;
17'h45cd:	data_out=16'h45;
17'h45ce:	data_out=16'h80b0;
17'h45cf:	data_out=16'h120;
17'h45d0:	data_out=16'ha;
17'h45d1:	data_out=16'h8131;
17'h45d2:	data_out=16'h8028;
17'h45d3:	data_out=16'h816f;
17'h45d4:	data_out=16'h813c;
17'h45d5:	data_out=16'h819f;
17'h45d6:	data_out=16'h80ff;
17'h45d7:	data_out=16'h80ce;
17'h45d8:	data_out=16'h8193;
17'h45d9:	data_out=16'h1b;
17'h45da:	data_out=16'h813a;
17'h45db:	data_out=16'h80aa;
17'h45dc:	data_out=16'h80a9;
17'h45dd:	data_out=16'h80a6;
17'h45de:	data_out=16'h8088;
17'h45df:	data_out=16'h806d;
17'h45e0:	data_out=16'h80db;
17'h45e1:	data_out=16'h8070;
17'h45e2:	data_out=16'h8153;
17'h45e3:	data_out=16'h817e;
17'h45e4:	data_out=16'h807c;
17'h45e5:	data_out=16'h119;
17'h45e6:	data_out=16'h182;
17'h45e7:	data_out=16'h80d8;
17'h45e8:	data_out=16'h802b;
17'h45e9:	data_out=16'h81b4;
17'h45ea:	data_out=16'h802f;
17'h45eb:	data_out=16'h8011;
17'h45ec:	data_out=16'h810c;
17'h45ed:	data_out=16'h8191;
17'h45ee:	data_out=16'h8021;
17'h45ef:	data_out=16'h22;
17'h45f0:	data_out=16'h801f;
17'h45f1:	data_out=16'h8189;
17'h45f2:	data_out=16'h8006;
17'h45f3:	data_out=16'h4;
17'h45f4:	data_out=16'haa;
17'h45f5:	data_out=16'h8088;
17'h45f6:	data_out=16'h8137;
17'h45f7:	data_out=16'h7c;
17'h45f8:	data_out=16'hb4;
17'h45f9:	data_out=16'h81af;
17'h45fa:	data_out=16'h8184;
17'h45fb:	data_out=16'h8028;
17'h45fc:	data_out=16'h809c;
17'h45fd:	data_out=16'h802e;
17'h45fe:	data_out=16'h80a1;
17'h45ff:	data_out=16'h2d;
17'h4600:	data_out=16'h3;
17'h4601:	data_out=16'h0;
17'h4602:	data_out=16'h0;
17'h4603:	data_out=16'h8004;
17'h4604:	data_out=16'h0;
17'h4605:	data_out=16'h8005;
17'h4606:	data_out=16'h0;
17'h4607:	data_out=16'h3;
17'h4608:	data_out=16'h3;
17'h4609:	data_out=16'h2;
17'h460a:	data_out=16'h5;
17'h460b:	data_out=16'h9;
17'h460c:	data_out=16'h3;
17'h460d:	data_out=16'h2;
17'h460e:	data_out=16'h8004;
17'h460f:	data_out=16'h2;
17'h4610:	data_out=16'h8;
17'h4611:	data_out=16'h8002;
17'h4612:	data_out=16'h8006;
17'h4613:	data_out=16'h8005;
17'h4614:	data_out=16'h9;
17'h4615:	data_out=16'h8009;
17'h4616:	data_out=16'h8002;
17'h4617:	data_out=16'h8004;
17'h4618:	data_out=16'h6;
17'h4619:	data_out=16'h8001;
17'h461a:	data_out=16'h3;
17'h461b:	data_out=16'h8003;
17'h461c:	data_out=16'h7;
17'h461d:	data_out=16'h8008;
17'h461e:	data_out=16'h4;
17'h461f:	data_out=16'h2;
17'h4620:	data_out=16'h2;
17'h4621:	data_out=16'h8005;
17'h4622:	data_out=16'h7;
17'h4623:	data_out=16'h8007;
17'h4624:	data_out=16'h8001;
17'h4625:	data_out=16'h8002;
17'h4626:	data_out=16'h5;
17'h4627:	data_out=16'h8007;
17'h4628:	data_out=16'h9;
17'h4629:	data_out=16'h1;
17'h462a:	data_out=16'h8008;
17'h462b:	data_out=16'h3;
17'h462c:	data_out=16'h8006;
17'h462d:	data_out=16'h8003;
17'h462e:	data_out=16'h8004;
17'h462f:	data_out=16'h8007;
17'h4630:	data_out=16'h5;
17'h4631:	data_out=16'h8001;
17'h4632:	data_out=16'h8002;
17'h4633:	data_out=16'h4;
17'h4634:	data_out=16'h8000;
17'h4635:	data_out=16'h5;
17'h4636:	data_out=16'h8009;
17'h4637:	data_out=16'h8003;
17'h4638:	data_out=16'h8005;
17'h4639:	data_out=16'h3;
17'h463a:	data_out=16'h3;
17'h463b:	data_out=16'h8007;
17'h463c:	data_out=16'h5;
17'h463d:	data_out=16'h8002;
17'h463e:	data_out=16'h4;
17'h463f:	data_out=16'h8003;
17'h4640:	data_out=16'h2;
17'h4641:	data_out=16'h2;
17'h4642:	data_out=16'h8001;
17'h4643:	data_out=16'h8008;
17'h4644:	data_out=16'h9;
17'h4645:	data_out=16'h8005;
17'h4646:	data_out=16'h8006;
17'h4647:	data_out=16'h9;
17'h4648:	data_out=16'h5;
17'h4649:	data_out=16'h8005;
17'h464a:	data_out=16'h3;
17'h464b:	data_out=16'h8;
17'h464c:	data_out=16'h1;
17'h464d:	data_out=16'h8;
17'h464e:	data_out=16'h8008;
17'h464f:	data_out=16'h8003;
17'h4650:	data_out=16'h8002;
17'h4651:	data_out=16'h8001;
17'h4652:	data_out=16'h8008;
17'h4653:	data_out=16'h7;
17'h4654:	data_out=16'h8005;
17'h4655:	data_out=16'h8007;
17'h4656:	data_out=16'h8005;
17'h4657:	data_out=16'h8002;
17'h4658:	data_out=16'h5;
17'h4659:	data_out=16'h7;
17'h465a:	data_out=16'h0;
17'h465b:	data_out=16'h0;
17'h465c:	data_out=16'h8005;
17'h465d:	data_out=16'h8005;
17'h465e:	data_out=16'h7;
17'h465f:	data_out=16'h6;
17'h4660:	data_out=16'h6;
17'h4661:	data_out=16'h8004;
17'h4662:	data_out=16'h7;
17'h4663:	data_out=16'h5;
17'h4664:	data_out=16'h0;
17'h4665:	data_out=16'h8008;
17'h4666:	data_out=16'h5;
17'h4667:	data_out=16'h8004;
17'h4668:	data_out=16'h8004;
17'h4669:	data_out=16'h8001;
17'h466a:	data_out=16'h8004;
17'h466b:	data_out=16'h7;
17'h466c:	data_out=16'h8003;
17'h466d:	data_out=16'h8003;
17'h466e:	data_out=16'h8006;
17'h466f:	data_out=16'h5;
17'h4670:	data_out=16'h5;
17'h4671:	data_out=16'h8004;
17'h4672:	data_out=16'h3;
17'h4673:	data_out=16'h9;
17'h4674:	data_out=16'h8002;
17'h4675:	data_out=16'h7;
17'h4676:	data_out=16'h8002;
17'h4677:	data_out=16'h8007;
17'h4678:	data_out=16'h4;
17'h4679:	data_out=16'h8;
17'h467a:	data_out=16'h3;
17'h467b:	data_out=16'h8;
17'h467c:	data_out=16'h8006;
17'h467d:	data_out=16'h0;
17'h467e:	data_out=16'h5;
17'h467f:	data_out=16'h9;
17'h4680:	data_out=16'h6;
17'h4681:	data_out=16'h3;
17'h4682:	data_out=16'h5;
17'h4683:	data_out=16'h8003;
17'h4684:	data_out=16'h4;
17'h4685:	data_out=16'h1;
17'h4686:	data_out=16'h2;
17'h4687:	data_out=16'h8009;
17'h4688:	data_out=16'h8;
17'h4689:	data_out=16'h7;
17'h468a:	data_out=16'h7;
17'h468b:	data_out=16'h8003;
17'h468c:	data_out=16'h8005;
17'h468d:	data_out=16'h8008;
17'h468e:	data_out=16'h8007;
17'h468f:	data_out=16'h8008;
17'h4690:	data_out=16'h8003;
17'h4691:	data_out=16'h5;
17'h4692:	data_out=16'h8009;
17'h4693:	data_out=16'h4;
17'h4694:	data_out=16'h2;
17'h4695:	data_out=16'h8001;
17'h4696:	data_out=16'h6;
17'h4697:	data_out=16'h8003;
17'h4698:	data_out=16'h8002;
17'h4699:	data_out=16'h0;
17'h469a:	data_out=16'h8004;
17'h469b:	data_out=16'h1;
17'h469c:	data_out=16'h8009;
17'h469d:	data_out=16'h8007;
17'h469e:	data_out=16'h0;
17'h469f:	data_out=16'h6;
17'h46a0:	data_out=16'h5;
17'h46a1:	data_out=16'h8004;
17'h46a2:	data_out=16'h8006;
17'h46a3:	data_out=16'h0;
17'h46a4:	data_out=16'h6;
17'h46a5:	data_out=16'h6;
17'h46a6:	data_out=16'h1;
17'h46a7:	data_out=16'h5;
17'h46a8:	data_out=16'h4;
17'h46a9:	data_out=16'h8001;
17'h46aa:	data_out=16'h8007;
17'h46ab:	data_out=16'h8;
17'h46ac:	data_out=16'h0;
17'h46ad:	data_out=16'h8005;
17'h46ae:	data_out=16'h9;
17'h46af:	data_out=16'h6;
17'h46b0:	data_out=16'h8;
17'h46b1:	data_out=16'h8009;
17'h46b2:	data_out=16'h1;
17'h46b3:	data_out=16'h1;
17'h46b4:	data_out=16'h8001;
17'h46b5:	data_out=16'h8002;
17'h46b6:	data_out=16'h7;
17'h46b7:	data_out=16'h6;
17'h46b8:	data_out=16'h8;
17'h46b9:	data_out=16'h8005;
17'h46ba:	data_out=16'h8002;
17'h46bb:	data_out=16'h8;
17'h46bc:	data_out=16'h8004;
17'h46bd:	data_out=16'h7;
17'h46be:	data_out=16'h6;
17'h46bf:	data_out=16'h8007;
17'h46c0:	data_out=16'h8006;
17'h46c1:	data_out=16'h9;
17'h46c2:	data_out=16'h2;
17'h46c3:	data_out=16'h9;
17'h46c4:	data_out=16'h6;
17'h46c5:	data_out=16'h8006;
17'h46c6:	data_out=16'h5;
17'h46c7:	data_out=16'h0;
17'h46c8:	data_out=16'h2;
17'h46c9:	data_out=16'h7;
17'h46ca:	data_out=16'h8001;
17'h46cb:	data_out=16'h8007;
17'h46cc:	data_out=16'h8008;
17'h46cd:	data_out=16'h8001;
17'h46ce:	data_out=16'h8;
17'h46cf:	data_out=16'h8009;
17'h46d0:	data_out=16'h8000;
17'h46d1:	data_out=16'h0;
17'h46d2:	data_out=16'h2;
17'h46d3:	data_out=16'h8;
17'h46d4:	data_out=16'h8;
17'h46d5:	data_out=16'h0;
17'h46d6:	data_out=16'h5;
17'h46d7:	data_out=16'h7;
17'h46d8:	data_out=16'h4;
17'h46d9:	data_out=16'h8006;
17'h46da:	data_out=16'h6;
17'h46db:	data_out=16'h8009;
17'h46dc:	data_out=16'h8009;
17'h46dd:	data_out=16'h3;
17'h46de:	data_out=16'h8007;
17'h46df:	data_out=16'h8006;
17'h46e0:	data_out=16'h2;
17'h46e1:	data_out=16'h4;
17'h46e2:	data_out=16'h8006;
17'h46e3:	data_out=16'h8001;
17'h46e4:	data_out=16'h7;
17'h46e5:	data_out=16'h8;
17'h46e6:	data_out=16'h8;
17'h46e7:	data_out=16'h8000;
17'h46e8:	data_out=16'h6;
17'h46e9:	data_out=16'h8002;
17'h46ea:	data_out=16'h2;
17'h46eb:	data_out=16'h7;
17'h46ec:	data_out=16'h7;
17'h46ed:	data_out=16'h1;
17'h46ee:	data_out=16'h8;
17'h46ef:	data_out=16'h8003;
17'h46f0:	data_out=16'h8008;
17'h46f1:	data_out=16'h0;
17'h46f2:	data_out=16'h8004;
17'h46f3:	data_out=16'h8009;
17'h46f4:	data_out=16'h8009;
17'h46f5:	data_out=16'h8008;
17'h46f6:	data_out=16'h7;
17'h46f7:	data_out=16'h4;
17'h46f8:	data_out=16'h8005;
17'h46f9:	data_out=16'h4;
17'h46fa:	data_out=16'h5;
17'h46fb:	data_out=16'h8004;
17'h46fc:	data_out=16'h8003;
17'h46fd:	data_out=16'h7;
17'h46fe:	data_out=16'h8001;
17'h46ff:	data_out=16'h9;
17'h4700:	data_out=16'h12;
17'h4701:	data_out=16'h6a;
17'h4702:	data_out=16'h38;
17'h4703:	data_out=16'h6e;
17'h4704:	data_out=16'h4d;
17'h4705:	data_out=16'h8a;
17'h4706:	data_out=16'h5e;
17'h4707:	data_out=16'h62;
17'h4708:	data_out=16'ha;
17'h4709:	data_out=16'h2a;
17'h470a:	data_out=16'h2e;
17'h470b:	data_out=16'h76;
17'h470c:	data_out=16'h1c;
17'h470d:	data_out=16'h5b;
17'h470e:	data_out=16'h15;
17'h470f:	data_out=16'h5d;
17'h4710:	data_out=16'h5a;
17'h4711:	data_out=16'h51;
17'h4712:	data_out=16'h7a;
17'h4713:	data_out=16'h84;
17'h4714:	data_out=16'hb8;
17'h4715:	data_out=16'h46;
17'h4716:	data_out=16'h69;
17'h4717:	data_out=16'hbd;
17'h4718:	data_out=16'h1c;
17'h4719:	data_out=16'h14;
17'h471a:	data_out=16'h50;
17'h471b:	data_out=16'h85;
17'h471c:	data_out=16'h95;
17'h471d:	data_out=16'h64;
17'h471e:	data_out=16'h7e;
17'h471f:	data_out=16'h7c;
17'h4720:	data_out=16'hb4;
17'h4721:	data_out=16'h1f;
17'h4722:	data_out=16'h87;
17'h4723:	data_out=16'h801c;
17'h4724:	data_out=16'h8011;
17'h4725:	data_out=16'h4c;
17'h4726:	data_out=16'hc;
17'h4727:	data_out=16'h6f;
17'h4728:	data_out=16'h26;
17'h4729:	data_out=16'h60;
17'h472a:	data_out=16'h44;
17'h472b:	data_out=16'h32;
17'h472c:	data_out=16'h5a;
17'h472d:	data_out=16'h34;
17'h472e:	data_out=16'h68;
17'h472f:	data_out=16'hac;
17'h4730:	data_out=16'hd4;
17'h4731:	data_out=16'h2a;
17'h4732:	data_out=16'hde;
17'h4733:	data_out=16'hbb;
17'h4734:	data_out=16'h30;
17'h4735:	data_out=16'h42;
17'h4736:	data_out=16'h46;
17'h4737:	data_out=16'h50;
17'h4738:	data_out=16'h53;
17'h4739:	data_out=16'h78;
17'h473a:	data_out=16'h43;
17'h473b:	data_out=16'h1e;
17'h473c:	data_out=16'h61;
17'h473d:	data_out=16'h5f;
17'h473e:	data_out=16'h1c;
17'h473f:	data_out=16'h76;
17'h4740:	data_out=16'h80;
17'h4741:	data_out=16'h58;
17'h4742:	data_out=16'h8002;
17'h4743:	data_out=16'h5e;
17'h4744:	data_out=16'h49;
17'h4745:	data_out=16'h48;
17'h4746:	data_out=16'h71;
17'h4747:	data_out=16'h31;
17'h4748:	data_out=16'h6f;
17'h4749:	data_out=16'h58;
17'h474a:	data_out=16'h25;
17'h474b:	data_out=16'h8001;
17'h474c:	data_out=16'h2d;
17'h474d:	data_out=16'h92;
17'h474e:	data_out=16'h55;
17'h474f:	data_out=16'h39;
17'h4750:	data_out=16'h5b;
17'h4751:	data_out=16'h57;
17'h4752:	data_out=16'hc;
17'h4753:	data_out=16'hb2;
17'h4754:	data_out=16'hc3;
17'h4755:	data_out=16'h3b;
17'h4756:	data_out=16'hb8;
17'h4757:	data_out=16'h60;
17'h4758:	data_out=16'h33;
17'h4759:	data_out=16'h7d;
17'h475a:	data_out=16'h60;
17'h475b:	data_out=16'h70;
17'h475c:	data_out=16'h4c;
17'h475d:	data_out=16'h68;
17'h475e:	data_out=16'hce;
17'h475f:	data_out=16'h38;
17'h4760:	data_out=16'h18;
17'h4761:	data_out=16'h83;
17'h4762:	data_out=16'h6c;
17'h4763:	data_out=16'hba;
17'h4764:	data_out=16'h54;
17'h4765:	data_out=16'h41;
17'h4766:	data_out=16'h28;
17'h4767:	data_out=16'h76;
17'h4768:	data_out=16'h25;
17'h4769:	data_out=16'h29;
17'h476a:	data_out=16'h22;
17'h476b:	data_out=16'h6c;
17'h476c:	data_out=16'h32;
17'h476d:	data_out=16'hb5;
17'h476e:	data_out=16'h1d;
17'h476f:	data_out=16'ha0;
17'h4770:	data_out=16'h16;
17'h4771:	data_out=16'h3a;
17'h4772:	data_out=16'h93;
17'h4773:	data_out=16'ha4;
17'h4774:	data_out=16'hce;
17'h4775:	data_out=16'h47;
17'h4776:	data_out=16'h29;
17'h4777:	data_out=16'h61;
17'h4778:	data_out=16'h4f;
17'h4779:	data_out=16'h59;
17'h477a:	data_out=16'hb5;
17'h477b:	data_out=16'h2b;
17'h477c:	data_out=16'h3b;
17'h477d:	data_out=16'h84;
17'h477e:	data_out=16'h45;
17'h477f:	data_out=16'h61;
17'h4780:	data_out=16'h8164;
17'h4781:	data_out=16'h12b;
17'h4782:	data_out=16'h82af;
17'h4783:	data_out=16'h8047;
17'h4784:	data_out=16'h8083;
17'h4785:	data_out=16'h3b6;
17'h4786:	data_out=16'h1c3;
17'h4787:	data_out=16'h8142;
17'h4788:	data_out=16'h82a2;
17'h4789:	data_out=16'h83b8;
17'h478a:	data_out=16'h81ee;
17'h478b:	data_out=16'h2f2;
17'h478c:	data_out=16'h82e0;
17'h478d:	data_out=16'h6;
17'h478e:	data_out=16'h808b;
17'h478f:	data_out=16'h821b;
17'h4790:	data_out=16'h841d;
17'h4791:	data_out=16'h34;
17'h4792:	data_out=16'h8178;
17'h4793:	data_out=16'h8189;
17'h4794:	data_out=16'h2b5;
17'h4795:	data_out=16'h8102;
17'h4796:	data_out=16'h8117;
17'h4797:	data_out=16'h2ab;
17'h4798:	data_out=16'h817b;
17'h4799:	data_out=16'h51;
17'h479a:	data_out=16'h8008;
17'h479b:	data_out=16'h486;
17'h479c:	data_out=16'h419;
17'h479d:	data_out=16'h106;
17'h479e:	data_out=16'h1e0;
17'h479f:	data_out=16'h156;
17'h47a0:	data_out=16'h463;
17'h47a1:	data_out=16'h8082;
17'h47a2:	data_out=16'h8273;
17'h47a3:	data_out=16'h8576;
17'h47a4:	data_out=16'h8577;
17'h47a5:	data_out=16'h8360;
17'h47a6:	data_out=16'h84f2;
17'h47a7:	data_out=16'h2d5;
17'h47a8:	data_out=16'h806f;
17'h47a9:	data_out=16'h8133;
17'h47aa:	data_out=16'h8587;
17'h47ab:	data_out=16'h350;
17'h47ac:	data_out=16'h8089;
17'h47ad:	data_out=16'h8649;
17'h47ae:	data_out=16'h83a6;
17'h47af:	data_out=16'h1cd;
17'h47b0:	data_out=16'h8191;
17'h47b1:	data_out=16'h3ed;
17'h47b2:	data_out=16'h819b;
17'h47b3:	data_out=16'h2f1;
17'h47b4:	data_out=16'h125;
17'h47b5:	data_out=16'h80eb;
17'h47b6:	data_out=16'h81a2;
17'h47b7:	data_out=16'h823e;
17'h47b8:	data_out=16'h3d2;
17'h47b9:	data_out=16'h301;
17'h47ba:	data_out=16'h8533;
17'h47bb:	data_out=16'h9f;
17'h47bc:	data_out=16'h80f4;
17'h47bd:	data_out=16'h77;
17'h47be:	data_out=16'h806d;
17'h47bf:	data_out=16'h225;
17'h47c0:	data_out=16'h84ac;
17'h47c1:	data_out=16'ha7;
17'h47c2:	data_out=16'h876c;
17'h47c3:	data_out=16'h2bb;
17'h47c4:	data_out=16'hf9;
17'h47c5:	data_out=16'h80e1;
17'h47c6:	data_out=16'h83;
17'h47c7:	data_out=16'h84b7;
17'h47c8:	data_out=16'h81e4;
17'h47c9:	data_out=16'h8340;
17'h47ca:	data_out=16'h82b6;
17'h47cb:	data_out=16'h84ea;
17'h47cc:	data_out=16'h85ef;
17'h47cd:	data_out=16'h8239;
17'h47ce:	data_out=16'h8365;
17'h47cf:	data_out=16'h85ae;
17'h47d0:	data_out=16'h8200;
17'h47d1:	data_out=16'h5f;
17'h47d2:	data_out=16'h86a6;
17'h47d3:	data_out=16'h6c4;
17'h47d4:	data_out=16'h173;
17'h47d5:	data_out=16'h3c;
17'h47d6:	data_out=16'h8405;
17'h47d7:	data_out=16'h855a;
17'h47d8:	data_out=16'h81c6;
17'h47d9:	data_out=16'h8554;
17'h47da:	data_out=16'h4af;
17'h47db:	data_out=16'h4d7;
17'h47dc:	data_out=16'h358;
17'h47dd:	data_out=16'h8350;
17'h47de:	data_out=16'h14f;
17'h47df:	data_out=16'h809c;
17'h47e0:	data_out=16'h8653;
17'h47e1:	data_out=16'h2b5;
17'h47e2:	data_out=16'h3cc;
17'h47e3:	data_out=16'h2e8;
17'h47e4:	data_out=16'h10d;
17'h47e5:	data_out=16'h8056;
17'h47e6:	data_out=16'h2b;
17'h47e7:	data_out=16'h82ac;
17'h47e8:	data_out=16'h8082;
17'h47e9:	data_out=16'h835e;
17'h47ea:	data_out=16'h80a0;
17'h47eb:	data_out=16'h2ad;
17'h47ec:	data_out=16'h85ab;
17'h47ed:	data_out=16'h319;
17'h47ee:	data_out=16'h80a2;
17'h47ef:	data_out=16'hb;
17'h47f0:	data_out=16'h8092;
17'h47f1:	data_out=16'h822f;
17'h47f2:	data_out=16'h8166;
17'h47f3:	data_out=16'h134;
17'h47f4:	data_out=16'h819e;
17'h47f5:	data_out=16'h60b;
17'h47f6:	data_out=16'h81;
17'h47f7:	data_out=16'h8579;
17'h47f8:	data_out=16'h2b3;
17'h47f9:	data_out=16'h849f;
17'h47fa:	data_out=16'h2c4;
17'h47fb:	data_out=16'h8065;
17'h47fc:	data_out=16'h15;
17'h47fd:	data_out=16'h408;
17'h47fe:	data_out=16'h82c5;
17'h47ff:	data_out=16'h831a;
17'h4800:	data_out=16'h8a00;
17'h4801:	data_out=16'h8a00;
17'h4802:	data_out=16'h8780;
17'h4803:	data_out=16'h84d5;
17'h4804:	data_out=16'h467;
17'h4805:	data_out=16'h7f3;
17'h4806:	data_out=16'h84a;
17'h4807:	data_out=16'h1a2;
17'h4808:	data_out=16'h89fb;
17'h4809:	data_out=16'h87a7;
17'h480a:	data_out=16'h8a00;
17'h480b:	data_out=16'ha00;
17'h480c:	data_out=16'h28c;
17'h480d:	data_out=16'h1e9;
17'h480e:	data_out=16'h8265;
17'h480f:	data_out=16'h86b6;
17'h4810:	data_out=16'h87ec;
17'h4811:	data_out=16'h37d;
17'h4812:	data_out=16'h107;
17'h4813:	data_out=16'h8370;
17'h4814:	data_out=16'h207;
17'h4815:	data_out=16'h868a;
17'h4816:	data_out=16'h89ec;
17'h4817:	data_out=16'h463;
17'h4818:	data_out=16'h8443;
17'h4819:	data_out=16'h6f4;
17'h481a:	data_out=16'h666;
17'h481b:	data_out=16'h9ad;
17'h481c:	data_out=16'h8194;
17'h481d:	data_out=16'h867c;
17'h481e:	data_out=16'h8b;
17'h481f:	data_out=16'h26d;
17'h4820:	data_out=16'h451;
17'h4821:	data_out=16'h8203;
17'h4822:	data_out=16'h826f;
17'h4823:	data_out=16'h8a00;
17'h4824:	data_out=16'h8a00;
17'h4825:	data_out=16'h841e;
17'h4826:	data_out=16'h8a00;
17'h4827:	data_out=16'h80b4;
17'h4828:	data_out=16'h8157;
17'h4829:	data_out=16'h83c3;
17'h482a:	data_out=16'h8a00;
17'h482b:	data_out=16'h7de;
17'h482c:	data_out=16'h8842;
17'h482d:	data_out=16'h8a00;
17'h482e:	data_out=16'h8547;
17'h482f:	data_out=16'h25a;
17'h4830:	data_out=16'h130;
17'h4831:	data_out=16'h57d;
17'h4832:	data_out=16'he9;
17'h4833:	data_out=16'h287;
17'h4834:	data_out=16'h8608;
17'h4835:	data_out=16'h2f1;
17'h4836:	data_out=16'h8a00;
17'h4837:	data_out=16'h86ac;
17'h4838:	data_out=16'h465;
17'h4839:	data_out=16'h27b;
17'h483a:	data_out=16'h8828;
17'h483b:	data_out=16'h8337;
17'h483c:	data_out=16'h89bc;
17'h483d:	data_out=16'h88eb;
17'h483e:	data_out=16'h813e;
17'h483f:	data_out=16'h7e0;
17'h4840:	data_out=16'h8340;
17'h4841:	data_out=16'h81df;
17'h4842:	data_out=16'h8925;
17'h4843:	data_out=16'h9a8;
17'h4844:	data_out=16'h8115;
17'h4845:	data_out=16'h86bb;
17'h4846:	data_out=16'h8524;
17'h4847:	data_out=16'h8701;
17'h4848:	data_out=16'h5d1;
17'h4849:	data_out=16'h83ca;
17'h484a:	data_out=16'h358;
17'h484b:	data_out=16'hcc;
17'h484c:	data_out=16'h84c8;
17'h484d:	data_out=16'h81ce;
17'h484e:	data_out=16'h85cc;
17'h484f:	data_out=16'h851e;
17'h4850:	data_out=16'h8088;
17'h4851:	data_out=16'h848a;
17'h4852:	data_out=16'h8a00;
17'h4853:	data_out=16'ha00;
17'h4854:	data_out=16'h848e;
17'h4855:	data_out=16'h8943;
17'h4856:	data_out=16'h8a00;
17'h4857:	data_out=16'h8a00;
17'h4858:	data_out=16'h89fa;
17'h4859:	data_out=16'h8962;
17'h485a:	data_out=16'h9fa;
17'h485b:	data_out=16'h8243;
17'h485c:	data_out=16'h72e;
17'h485d:	data_out=16'h8a00;
17'h485e:	data_out=16'h1db;
17'h485f:	data_out=16'h829b;
17'h4860:	data_out=16'h8a00;
17'h4861:	data_out=16'h829c;
17'h4862:	data_out=16'h90c;
17'h4863:	data_out=16'h3ab;
17'h4864:	data_out=16'h80;
17'h4865:	data_out=16'h6dd;
17'h4866:	data_out=16'h8d4;
17'h4867:	data_out=16'h80f8;
17'h4868:	data_out=16'h81bb;
17'h4869:	data_out=16'h8a00;
17'h486a:	data_out=16'h82de;
17'h486b:	data_out=16'h590;
17'h486c:	data_out=16'h8a00;
17'h486d:	data_out=16'h333;
17'h486e:	data_out=16'h82dc;
17'h486f:	data_out=16'h3dc;
17'h4870:	data_out=16'h828a;
17'h4871:	data_out=16'h8247;
17'h4872:	data_out=16'h874d;
17'h4873:	data_out=16'h80c0;
17'h4874:	data_out=16'h112;
17'h4875:	data_out=16'h795;
17'h4876:	data_out=16'h4dc;
17'h4877:	data_out=16'h87cf;
17'h4878:	data_out=16'h9ff;
17'h4879:	data_out=16'h896a;
17'h487a:	data_out=16'h2eb;
17'h487b:	data_out=16'h8130;
17'h487c:	data_out=16'h8230;
17'h487d:	data_out=16'ha00;
17'h487e:	data_out=16'h86e7;
17'h487f:	data_out=16'h85b7;
17'h4880:	data_out=16'h8a00;
17'h4881:	data_out=16'h8a00;
17'h4882:	data_out=16'h88d9;
17'h4883:	data_out=16'h170;
17'h4884:	data_out=16'h92;
17'h4885:	data_out=16'h9ea;
17'h4886:	data_out=16'ha00;
17'h4887:	data_out=16'h81bb;
17'h4888:	data_out=16'h891e;
17'h4889:	data_out=16'h89fc;
17'h488a:	data_out=16'h8a00;
17'h488b:	data_out=16'h9fd;
17'h488c:	data_out=16'h6c7;
17'h488d:	data_out=16'h9ce;
17'h488e:	data_out=16'h8520;
17'h488f:	data_out=16'h86b9;
17'h4890:	data_out=16'h89ff;
17'h4891:	data_out=16'h816b;
17'h4892:	data_out=16'h3fe;
17'h4893:	data_out=16'h492;
17'h4894:	data_out=16'h9fb;
17'h4895:	data_out=16'h88b2;
17'h4896:	data_out=16'h8a00;
17'h4897:	data_out=16'h9f6;
17'h4898:	data_out=16'h846f;
17'h4899:	data_out=16'ha00;
17'h489a:	data_out=16'h4a4;
17'h489b:	data_out=16'h9f5;
17'h489c:	data_out=16'h332;
17'h489d:	data_out=16'h8614;
17'h489e:	data_out=16'h9c1;
17'h489f:	data_out=16'h43d;
17'h48a0:	data_out=16'h9f5;
17'h48a1:	data_out=16'h8499;
17'h48a2:	data_out=16'h8791;
17'h48a3:	data_out=16'h8a00;
17'h48a4:	data_out=16'h8a00;
17'h48a5:	data_out=16'h8a00;
17'h48a6:	data_out=16'h8a00;
17'h48a7:	data_out=16'h710;
17'h48a8:	data_out=16'h829f;
17'h48a9:	data_out=16'h1f2;
17'h48aa:	data_out=16'h89fe;
17'h48ab:	data_out=16'h9ff;
17'h48ac:	data_out=16'h896e;
17'h48ad:	data_out=16'h8a00;
17'h48ae:	data_out=16'h8180;
17'h48af:	data_out=16'h9f8;
17'h48b0:	data_out=16'h84c8;
17'h48b1:	data_out=16'h8d5;
17'h48b2:	data_out=16'h8618;
17'h48b3:	data_out=16'ha00;
17'h48b4:	data_out=16'h8a00;
17'h48b5:	data_out=16'h3d4;
17'h48b6:	data_out=16'h87a6;
17'h48b7:	data_out=16'h8880;
17'h48b8:	data_out=16'h752;
17'h48b9:	data_out=16'ha00;
17'h48ba:	data_out=16'h89ff;
17'h48bb:	data_out=16'h8680;
17'h48bc:	data_out=16'h89fe;
17'h48bd:	data_out=16'h89ff;
17'h48be:	data_out=16'h827f;
17'h48bf:	data_out=16'h9e8;
17'h48c0:	data_out=16'h8a00;
17'h48c1:	data_out=16'h4c1;
17'h48c2:	data_out=16'h8a00;
17'h48c3:	data_out=16'ha00;
17'h48c4:	data_out=16'h236;
17'h48c5:	data_out=16'h88f5;
17'h48c6:	data_out=16'h8a00;
17'h48c7:	data_out=16'h89f9;
17'h48c8:	data_out=16'h9ff;
17'h48c9:	data_out=16'h8a00;
17'h48ca:	data_out=16'h600;
17'h48cb:	data_out=16'h1d1;
17'h48cc:	data_out=16'h8a00;
17'h48cd:	data_out=16'h85f7;
17'h48ce:	data_out=16'h8424;
17'h48cf:	data_out=16'h8a00;
17'h48d0:	data_out=16'h885d;
17'h48d1:	data_out=16'h8014;
17'h48d2:	data_out=16'h8a00;
17'h48d3:	data_out=16'ha00;
17'h48d4:	data_out=16'h2e0;
17'h48d5:	data_out=16'h87f1;
17'h48d6:	data_out=16'h8a00;
17'h48d7:	data_out=16'h8a00;
17'h48d8:	data_out=16'h896e;
17'h48d9:	data_out=16'h8a00;
17'h48da:	data_out=16'ha00;
17'h48db:	data_out=16'h816a;
17'h48dc:	data_out=16'h9f7;
17'h48dd:	data_out=16'h8a00;
17'h48de:	data_out=16'h9d9;
17'h48df:	data_out=16'h818d;
17'h48e0:	data_out=16'h8a00;
17'h48e1:	data_out=16'h810b;
17'h48e2:	data_out=16'h9ea;
17'h48e3:	data_out=16'ha00;
17'h48e4:	data_out=16'h83ea;
17'h48e5:	data_out=16'h538;
17'h48e6:	data_out=16'ha00;
17'h48e7:	data_out=16'h3d;
17'h48e8:	data_out=16'h83db;
17'h48e9:	data_out=16'h89fc;
17'h48ea:	data_out=16'h8598;
17'h48eb:	data_out=16'h51e;
17'h48ec:	data_out=16'h8a00;
17'h48ed:	data_out=16'ha00;
17'h48ee:	data_out=16'h8597;
17'h48ef:	data_out=16'h430;
17'h48f0:	data_out=16'h8553;
17'h48f1:	data_out=16'h566;
17'h48f2:	data_out=16'h8a00;
17'h48f3:	data_out=16'h859e;
17'h48f4:	data_out=16'h84b3;
17'h48f5:	data_out=16'h9e3;
17'h48f6:	data_out=16'h9fb;
17'h48f7:	data_out=16'h89ff;
17'h48f8:	data_out=16'h9fc;
17'h48f9:	data_out=16'h84fb;
17'h48fa:	data_out=16'ha00;
17'h48fb:	data_out=16'h824c;
17'h48fc:	data_out=16'h58;
17'h48fd:	data_out=16'ha00;
17'h48fe:	data_out=16'h89ff;
17'h48ff:	data_out=16'h89e0;
17'h4900:	data_out=16'h8a00;
17'h4901:	data_out=16'h86cd;
17'h4902:	data_out=16'h854b;
17'h4903:	data_out=16'h87a0;
17'h4904:	data_out=16'h9bc;
17'h4905:	data_out=16'h9f6;
17'h4906:	data_out=16'h85b;
17'h4907:	data_out=16'ha00;
17'h4908:	data_out=16'h86dc;
17'h4909:	data_out=16'h89f9;
17'h490a:	data_out=16'h8a00;
17'h490b:	data_out=16'ha00;
17'h490c:	data_out=16'ha00;
17'h490d:	data_out=16'h7c8;
17'h490e:	data_out=16'h814f;
17'h490f:	data_out=16'h802d;
17'h4910:	data_out=16'h89fe;
17'h4911:	data_out=16'h62e;
17'h4912:	data_out=16'h9fd;
17'h4913:	data_out=16'h8270;
17'h4914:	data_out=16'h9fd;
17'h4915:	data_out=16'h87e3;
17'h4916:	data_out=16'h8a00;
17'h4917:	data_out=16'h9f9;
17'h4918:	data_out=16'h8357;
17'h4919:	data_out=16'ha00;
17'h491a:	data_out=16'ha00;
17'h491b:	data_out=16'h9da;
17'h491c:	data_out=16'h129;
17'h491d:	data_out=16'h167;
17'h491e:	data_out=16'h9e5;
17'h491f:	data_out=16'ha00;
17'h4920:	data_out=16'h9e7;
17'h4921:	data_out=16'h80ac;
17'h4922:	data_out=16'h1de;
17'h4923:	data_out=16'h89fe;
17'h4924:	data_out=16'h89fe;
17'h4925:	data_out=16'h89ff;
17'h4926:	data_out=16'h8a00;
17'h4927:	data_out=16'h9fb;
17'h4928:	data_out=16'h43;
17'h4929:	data_out=16'h9b;
17'h492a:	data_out=16'h84f2;
17'h492b:	data_out=16'ha00;
17'h492c:	data_out=16'h89ff;
17'h492d:	data_out=16'h8a00;
17'h492e:	data_out=16'h6da;
17'h492f:	data_out=16'h9f7;
17'h4930:	data_out=16'h3b5;
17'h4931:	data_out=16'h959;
17'h4932:	data_out=16'h14c;
17'h4933:	data_out=16'ha00;
17'h4934:	data_out=16'h863d;
17'h4935:	data_out=16'h739;
17'h4936:	data_out=16'h8511;
17'h4937:	data_out=16'h852f;
17'h4938:	data_out=16'h9ff;
17'h4939:	data_out=16'h9ff;
17'h493a:	data_out=16'h833b;
17'h493b:	data_out=16'hb9;
17'h493c:	data_out=16'h89f5;
17'h493d:	data_out=16'h898c;
17'h493e:	data_out=16'h49;
17'h493f:	data_out=16'h9f4;
17'h4940:	data_out=16'h891b;
17'h4941:	data_out=16'h53;
17'h4942:	data_out=16'h89ff;
17'h4943:	data_out=16'h93b;
17'h4944:	data_out=16'h613;
17'h4945:	data_out=16'h8818;
17'h4946:	data_out=16'h89a3;
17'h4947:	data_out=16'h86c4;
17'h4948:	data_out=16'h9f9;
17'h4949:	data_out=16'h89ff;
17'h494a:	data_out=16'ha00;
17'h494b:	data_out=16'h1b0;
17'h494c:	data_out=16'h8a00;
17'h494d:	data_out=16'h369;
17'h494e:	data_out=16'h7d4;
17'h494f:	data_out=16'h8a00;
17'h4950:	data_out=16'h80c4;
17'h4951:	data_out=16'h8185;
17'h4952:	data_out=16'h89ff;
17'h4953:	data_out=16'ha00;
17'h4954:	data_out=16'h915;
17'h4955:	data_out=16'h890f;
17'h4956:	data_out=16'h89ff;
17'h4957:	data_out=16'h8a00;
17'h4958:	data_out=16'h89f3;
17'h4959:	data_out=16'h8a00;
17'h495a:	data_out=16'ha00;
17'h495b:	data_out=16'h511;
17'h495c:	data_out=16'h9f3;
17'h495d:	data_out=16'h895a;
17'h495e:	data_out=16'h9d4;
17'h495f:	data_out=16'h38a;
17'h4960:	data_out=16'h8a00;
17'h4961:	data_out=16'h2f0;
17'h4962:	data_out=16'h9e5;
17'h4963:	data_out=16'ha00;
17'h4964:	data_out=16'h847b;
17'h4965:	data_out=16'h45a;
17'h4966:	data_out=16'ha00;
17'h4967:	data_out=16'h897;
17'h4968:	data_out=16'h8037;
17'h4969:	data_out=16'h89fb;
17'h496a:	data_out=16'h82c7;
17'h496b:	data_out=16'h9c1;
17'h496c:	data_out=16'h8a00;
17'h496d:	data_out=16'ha00;
17'h496e:	data_out=16'h8297;
17'h496f:	data_out=16'h1a8;
17'h4970:	data_out=16'h8199;
17'h4971:	data_out=16'h9fd;
17'h4972:	data_out=16'h8a00;
17'h4973:	data_out=16'h8982;
17'h4974:	data_out=16'h3f8;
17'h4975:	data_out=16'h8029;
17'h4976:	data_out=16'h9fe;
17'h4977:	data_out=16'h89fa;
17'h4978:	data_out=16'ha00;
17'h4979:	data_out=16'h494;
17'h497a:	data_out=16'ha00;
17'h497b:	data_out=16'h4a;
17'h497c:	data_out=16'h39f;
17'h497d:	data_out=16'ha00;
17'h497e:	data_out=16'h89ff;
17'h497f:	data_out=16'h8630;
17'h4980:	data_out=16'h89fe;
17'h4981:	data_out=16'h8416;
17'h4982:	data_out=16'h83b9;
17'h4983:	data_out=16'h89fd;
17'h4984:	data_out=16'ha00;
17'h4985:	data_out=16'h9f2;
17'h4986:	data_out=16'he0;
17'h4987:	data_out=16'ha00;
17'h4988:	data_out=16'h87eb;
17'h4989:	data_out=16'h892c;
17'h498a:	data_out=16'h88e6;
17'h498b:	data_out=16'h2c9;
17'h498c:	data_out=16'h9fd;
17'h498d:	data_out=16'h89eb;
17'h498e:	data_out=16'h487;
17'h498f:	data_out=16'h349;
17'h4990:	data_out=16'h89fe;
17'h4991:	data_out=16'h1f7;
17'h4992:	data_out=16'h9f0;
17'h4993:	data_out=16'h89e9;
17'h4994:	data_out=16'h9e8;
17'h4995:	data_out=16'h89ae;
17'h4996:	data_out=16'h89f5;
17'h4997:	data_out=16'h84e;
17'h4998:	data_out=16'h828f;
17'h4999:	data_out=16'h9fd;
17'h499a:	data_out=16'ha00;
17'h499b:	data_out=16'h92c;
17'h499c:	data_out=16'h8735;
17'h499d:	data_out=16'h182;
17'h499e:	data_out=16'h9e7;
17'h499f:	data_out=16'h9ff;
17'h49a0:	data_out=16'h9d4;
17'h49a1:	data_out=16'h4e4;
17'h49a2:	data_out=16'h9eb;
17'h49a3:	data_out=16'h89fa;
17'h49a4:	data_out=16'h89fa;
17'h49a5:	data_out=16'h89fe;
17'h49a6:	data_out=16'h8a00;
17'h49a7:	data_out=16'h9eb;
17'h49a8:	data_out=16'h570;
17'h49a9:	data_out=16'h13f;
17'h49aa:	data_out=16'h80cc;
17'h49ab:	data_out=16'ha00;
17'h49ac:	data_out=16'h89f7;
17'h49ad:	data_out=16'h861a;
17'h49ae:	data_out=16'ha00;
17'h49af:	data_out=16'h9f6;
17'h49b0:	data_out=16'h9ee;
17'h49b1:	data_out=16'h5c5;
17'h49b2:	data_out=16'ha00;
17'h49b3:	data_out=16'h9fb;
17'h49b4:	data_out=16'h896a;
17'h49b5:	data_out=16'h585;
17'h49b6:	data_out=16'h84e9;
17'h49b7:	data_out=16'h8403;
17'h49b8:	data_out=16'h9fc;
17'h49b9:	data_out=16'h9f1;
17'h49ba:	data_out=16'h6d2;
17'h49bb:	data_out=16'h48a;
17'h49bc:	data_out=16'h89eb;
17'h49bd:	data_out=16'h8988;
17'h49be:	data_out=16'h573;
17'h49bf:	data_out=16'h9be;
17'h49c0:	data_out=16'h8245;
17'h49c1:	data_out=16'h89e0;
17'h49c2:	data_out=16'h89fd;
17'h49c3:	data_out=16'h464;
17'h49c4:	data_out=16'h8248;
17'h49c5:	data_out=16'h89fc;
17'h49c6:	data_out=16'h807f;
17'h49c7:	data_out=16'h8406;
17'h49c8:	data_out=16'h9e2;
17'h49c9:	data_out=16'h89fe;
17'h49ca:	data_out=16'ha00;
17'h49cb:	data_out=16'h8856;
17'h49cc:	data_out=16'h89ff;
17'h49cd:	data_out=16'h9f1;
17'h49ce:	data_out=16'ha00;
17'h49cf:	data_out=16'h89fe;
17'h49d0:	data_out=16'h848;
17'h49d1:	data_out=16'h89f0;
17'h49d2:	data_out=16'h89e3;
17'h49d3:	data_out=16'ha00;
17'h49d4:	data_out=16'h9fd;
17'h49d5:	data_out=16'h89dc;
17'h49d6:	data_out=16'h89f9;
17'h49d7:	data_out=16'h89f4;
17'h49d8:	data_out=16'h89eb;
17'h49d9:	data_out=16'h88d4;
17'h49da:	data_out=16'h9ed;
17'h49db:	data_out=16'h9ef;
17'h49dc:	data_out=16'h9e4;
17'h49dd:	data_out=16'h8511;
17'h49de:	data_out=16'h9d7;
17'h49df:	data_out=16'h854;
17'h49e0:	data_out=16'h89ff;
17'h49e1:	data_out=16'h823c;
17'h49e2:	data_out=16'h22c;
17'h49e3:	data_out=16'h9fe;
17'h49e4:	data_out=16'h89fa;
17'h49e5:	data_out=16'h18d;
17'h49e6:	data_out=16'ha00;
17'h49e7:	data_out=16'h9f9;
17'h49e8:	data_out=16'h51f;
17'h49e9:	data_out=16'h89ea;
17'h49ea:	data_out=16'h43a;
17'h49eb:	data_out=16'h99b;
17'h49ec:	data_out=16'h89f4;
17'h49ed:	data_out=16'h9fe;
17'h49ee:	data_out=16'h43b;
17'h49ef:	data_out=16'h470;
17'h49f0:	data_out=16'h465;
17'h49f1:	data_out=16'ha00;
17'h49f2:	data_out=16'h8a00;
17'h49f3:	data_out=16'h87b1;
17'h49f4:	data_out=16'h9dc;
17'h49f5:	data_out=16'h8837;
17'h49f6:	data_out=16'h9fe;
17'h49f7:	data_out=16'h89c5;
17'h49f8:	data_out=16'ha00;
17'h49f9:	data_out=16'h99c;
17'h49fa:	data_out=16'h9f9;
17'h49fb:	data_out=16'h572;
17'h49fc:	data_out=16'h7d5;
17'h49fd:	data_out=16'ha00;
17'h49fe:	data_out=16'h8a00;
17'h49ff:	data_out=16'h8a4;
17'h4a00:	data_out=16'h89e6;
17'h4a01:	data_out=16'h17;
17'h4a02:	data_out=16'h8809;
17'h4a03:	data_out=16'h89f2;
17'h4a04:	data_out=16'ha00;
17'h4a05:	data_out=16'h9e5;
17'h4a06:	data_out=16'h89b7;
17'h4a07:	data_out=16'ha00;
17'h4a08:	data_out=16'h8890;
17'h4a09:	data_out=16'h8900;
17'h4a0a:	data_out=16'h81e8;
17'h4a0b:	data_out=16'h8867;
17'h4a0c:	data_out=16'h800c;
17'h4a0d:	data_out=16'h89f2;
17'h4a0e:	data_out=16'h53f;
17'h4a0f:	data_out=16'h83a5;
17'h4a10:	data_out=16'h89ed;
17'h4a11:	data_out=16'h9c1;
17'h4a12:	data_out=16'h48a;
17'h4a13:	data_out=16'h89f0;
17'h4a14:	data_out=16'h897d;
17'h4a15:	data_out=16'h87d5;
17'h4a16:	data_out=16'h89ee;
17'h4a17:	data_out=16'h8977;
17'h4a18:	data_out=16'h86ee;
17'h4a19:	data_out=16'ha00;
17'h4a1a:	data_out=16'ha00;
17'h4a1b:	data_out=16'h8056;
17'h4a1c:	data_out=16'h882e;
17'h4a1d:	data_out=16'h929;
17'h4a1e:	data_out=16'h824b;
17'h4a1f:	data_out=16'h9fe;
17'h4a20:	data_out=16'h9da;
17'h4a21:	data_out=16'h588;
17'h4a22:	data_out=16'h9d2;
17'h4a23:	data_out=16'h89ed;
17'h4a24:	data_out=16'h89ed;
17'h4a25:	data_out=16'h89f2;
17'h4a26:	data_out=16'h8a00;
17'h4a27:	data_out=16'h9fd;
17'h4a28:	data_out=16'h613;
17'h4a29:	data_out=16'h82b5;
17'h4a2a:	data_out=16'h83d3;
17'h4a2b:	data_out=16'ha00;
17'h4a2c:	data_out=16'h89f0;
17'h4a2d:	data_out=16'h853f;
17'h4a2e:	data_out=16'h9e8;
17'h4a2f:	data_out=16'h9f5;
17'h4a30:	data_out=16'h9f1;
17'h4a31:	data_out=16'h71a;
17'h4a32:	data_out=16'ha00;
17'h4a33:	data_out=16'h8223;
17'h4a34:	data_out=16'h8137;
17'h4a35:	data_out=16'h865;
17'h4a36:	data_out=16'h8607;
17'h4a37:	data_out=16'h87c6;
17'h4a38:	data_out=16'h9ff;
17'h4a39:	data_out=16'h94;
17'h4a3a:	data_out=16'h907;
17'h4a3b:	data_out=16'h9fe;
17'h4a3c:	data_out=16'h89f5;
17'h4a3d:	data_out=16'h937;
17'h4a3e:	data_out=16'h616;
17'h4a3f:	data_out=16'h9e5;
17'h4a40:	data_out=16'ha00;
17'h4a41:	data_out=16'h89d4;
17'h4a42:	data_out=16'h89e0;
17'h4a43:	data_out=16'h4ed;
17'h4a44:	data_out=16'h826f;
17'h4a45:	data_out=16'h88cc;
17'h4a46:	data_out=16'h873b;
17'h4a47:	data_out=16'h8475;
17'h4a48:	data_out=16'h94f;
17'h4a49:	data_out=16'h89fe;
17'h4a4a:	data_out=16'ha00;
17'h4a4b:	data_out=16'h89f7;
17'h4a4c:	data_out=16'h89ff;
17'h4a4d:	data_out=16'ha00;
17'h4a4e:	data_out=16'ha00;
17'h4a4f:	data_out=16'h89fe;
17'h4a50:	data_out=16'h7ca;
17'h4a51:	data_out=16'h89f9;
17'h4a52:	data_out=16'h8808;
17'h4a53:	data_out=16'ha00;
17'h4a54:	data_out=16'h9ff;
17'h4a55:	data_out=16'h89ee;
17'h4a56:	data_out=16'h89f5;
17'h4a57:	data_out=16'h8648;
17'h4a58:	data_out=16'h89f0;
17'h4a59:	data_out=16'h9f1;
17'h4a5a:	data_out=16'h89db;
17'h4a5b:	data_out=16'h9f5;
17'h4a5c:	data_out=16'h98c;
17'h4a5d:	data_out=16'h81e1;
17'h4a5e:	data_out=16'h9cc;
17'h4a5f:	data_out=16'ha00;
17'h4a60:	data_out=16'h89d3;
17'h4a61:	data_out=16'h8141;
17'h4a62:	data_out=16'h895c;
17'h4a63:	data_out=16'h16c;
17'h4a64:	data_out=16'h89eb;
17'h4a65:	data_out=16'h9e8;
17'h4a66:	data_out=16'ha00;
17'h4a67:	data_out=16'ha00;
17'h4a68:	data_out=16'h5bd;
17'h4a69:	data_out=16'h89e1;
17'h4a6a:	data_out=16'h51c;
17'h4a6b:	data_out=16'h9fa;
17'h4a6c:	data_out=16'h89c5;
17'h4a6d:	data_out=16'hfb;
17'h4a6e:	data_out=16'h51c;
17'h4a6f:	data_out=16'ha00;
17'h4a70:	data_out=16'h52a;
17'h4a71:	data_out=16'h9fe;
17'h4a72:	data_out=16'h8043;
17'h4a73:	data_out=16'h373;
17'h4a74:	data_out=16'h9d3;
17'h4a75:	data_out=16'h89ef;
17'h4a76:	data_out=16'ha00;
17'h4a77:	data_out=16'h89e6;
17'h4a78:	data_out=16'ha00;
17'h4a79:	data_out=16'h4a0;
17'h4a7a:	data_out=16'h824a;
17'h4a7b:	data_out=16'h614;
17'h4a7c:	data_out=16'h9e3;
17'h4a7d:	data_out=16'ha00;
17'h4a7e:	data_out=16'h8a00;
17'h4a7f:	data_out=16'h854;
17'h4a80:	data_out=16'h892e;
17'h4a81:	data_out=16'h9f9;
17'h4a82:	data_out=16'h865e;
17'h4a83:	data_out=16'h89eb;
17'h4a84:	data_out=16'h9ff;
17'h4a85:	data_out=16'h9e4;
17'h4a86:	data_out=16'h89f6;
17'h4a87:	data_out=16'h9fd;
17'h4a88:	data_out=16'h8899;
17'h4a89:	data_out=16'h89f8;
17'h4a8a:	data_out=16'h9ec;
17'h4a8b:	data_out=16'h89a8;
17'h4a8c:	data_out=16'h822b;
17'h4a8d:	data_out=16'h89f3;
17'h4a8e:	data_out=16'h6a2;
17'h4a8f:	data_out=16'h8213;
17'h4a90:	data_out=16'h89f6;
17'h4a91:	data_out=16'h2a1;
17'h4a92:	data_out=16'h8903;
17'h4a93:	data_out=16'h89e9;
17'h4a94:	data_out=16'h89cf;
17'h4a95:	data_out=16'h250;
17'h4a96:	data_out=16'h89ae;
17'h4a97:	data_out=16'h89c3;
17'h4a98:	data_out=16'h83f4;
17'h4a99:	data_out=16'ha00;
17'h4a9a:	data_out=16'ha00;
17'h4a9b:	data_out=16'h89e8;
17'h4a9c:	data_out=16'h89ef;
17'h4a9d:	data_out=16'h9f6;
17'h4a9e:	data_out=16'h889f;
17'h4a9f:	data_out=16'h91a;
17'h4aa0:	data_out=16'h9ce;
17'h4aa1:	data_out=16'h6b8;
17'h4aa2:	data_out=16'h828c;
17'h4aa3:	data_out=16'h8966;
17'h4aa4:	data_out=16'h8969;
17'h4aa5:	data_out=16'h89da;
17'h4aa6:	data_out=16'h89d9;
17'h4aa7:	data_out=16'h9db;
17'h4aa8:	data_out=16'h70b;
17'h4aa9:	data_out=16'h36f;
17'h4aaa:	data_out=16'h823d;
17'h4aab:	data_out=16'ha00;
17'h4aac:	data_out=16'h898c;
17'h4aad:	data_out=16'h8933;
17'h4aae:	data_out=16'h2fe;
17'h4aaf:	data_out=16'h9fc;
17'h4ab0:	data_out=16'h9e8;
17'h4ab1:	data_out=16'h6a0;
17'h4ab2:	data_out=16'h9e7;
17'h4ab3:	data_out=16'h88b4;
17'h4ab4:	data_out=16'h83dc;
17'h4ab5:	data_out=16'h83f;
17'h4ab6:	data_out=16'h8413;
17'h4ab7:	data_out=16'h87ed;
17'h4ab8:	data_out=16'h9d0;
17'h4ab9:	data_out=16'h8982;
17'h4aba:	data_out=16'h865;
17'h4abb:	data_out=16'h9f5;
17'h4abc:	data_out=16'h89d6;
17'h4abd:	data_out=16'h984;
17'h4abe:	data_out=16'h70d;
17'h4abf:	data_out=16'h9e5;
17'h4ac0:	data_out=16'ha00;
17'h4ac1:	data_out=16'h89d8;
17'h4ac2:	data_out=16'h89f7;
17'h4ac3:	data_out=16'he5;
17'h4ac4:	data_out=16'h191;
17'h4ac5:	data_out=16'h166;
17'h4ac6:	data_out=16'h89e1;
17'h4ac7:	data_out=16'h83f7;
17'h4ac8:	data_out=16'h589;
17'h4ac9:	data_out=16'h89ef;
17'h4aca:	data_out=16'ha00;
17'h4acb:	data_out=16'h89ef;
17'h4acc:	data_out=16'h89fa;
17'h4acd:	data_out=16'h847;
17'h4ace:	data_out=16'ha00;
17'h4acf:	data_out=16'h89f1;
17'h4ad0:	data_out=16'h374;
17'h4ad1:	data_out=16'h89f8;
17'h4ad2:	data_out=16'h8338;
17'h4ad3:	data_out=16'ha00;
17'h4ad4:	data_out=16'ha00;
17'h4ad5:	data_out=16'h89c9;
17'h4ad6:	data_out=16'h89f2;
17'h4ad7:	data_out=16'h33;
17'h4ad8:	data_out=16'h89f6;
17'h4ad9:	data_out=16'h9ab;
17'h4ada:	data_out=16'h89df;
17'h4adb:	data_out=16'h9f2;
17'h4adc:	data_out=16'h742;
17'h4add:	data_out=16'h479;
17'h4ade:	data_out=16'h9d3;
17'h4adf:	data_out=16'ha00;
17'h4ae0:	data_out=16'h8980;
17'h4ae1:	data_out=16'h180;
17'h4ae2:	data_out=16'h89b6;
17'h4ae3:	data_out=16'h879e;
17'h4ae4:	data_out=16'h89e5;
17'h4ae5:	data_out=16'h5b8;
17'h4ae6:	data_out=16'ha00;
17'h4ae7:	data_out=16'ha00;
17'h4ae8:	data_out=16'h6cb;
17'h4ae9:	data_out=16'h89e2;
17'h4aea:	data_out=16'h6aa;
17'h4aeb:	data_out=16'h9f7;
17'h4aec:	data_out=16'h85ee;
17'h4aed:	data_out=16'h87c4;
17'h4aee:	data_out=16'h6a9;
17'h4aef:	data_out=16'h9ff;
17'h4af0:	data_out=16'h69e;
17'h4af1:	data_out=16'h9ff;
17'h4af2:	data_out=16'h759;
17'h4af3:	data_out=16'h7e2;
17'h4af4:	data_out=16'h9bf;
17'h4af5:	data_out=16'h89f8;
17'h4af6:	data_out=16'ha00;
17'h4af7:	data_out=16'h89e6;
17'h4af8:	data_out=16'ha00;
17'h4af9:	data_out=16'h80a;
17'h4afa:	data_out=16'h88c5;
17'h4afb:	data_out=16'h70c;
17'h4afc:	data_out=16'ha00;
17'h4afd:	data_out=16'ha00;
17'h4afe:	data_out=16'h8a00;
17'h4aff:	data_out=16'h929;
17'h4b00:	data_out=16'h991;
17'h4b01:	data_out=16'ha00;
17'h4b02:	data_out=16'h89b9;
17'h4b03:	data_out=16'h89bb;
17'h4b04:	data_out=16'h9eb;
17'h4b05:	data_out=16'h9e6;
17'h4b06:	data_out=16'h89f3;
17'h4b07:	data_out=16'h3e2;
17'h4b08:	data_out=16'h89cb;
17'h4b09:	data_out=16'h89ff;
17'h4b0a:	data_out=16'h9f4;
17'h4b0b:	data_out=16'h897b;
17'h4b0c:	data_out=16'h8997;
17'h4b0d:	data_out=16'h8a00;
17'h4b0e:	data_out=16'h3f0;
17'h4b0f:	data_out=16'h8989;
17'h4b10:	data_out=16'h89ed;
17'h4b11:	data_out=16'h52a;
17'h4b12:	data_out=16'h89e6;
17'h4b13:	data_out=16'h89cf;
17'h4b14:	data_out=16'h8931;
17'h4b15:	data_out=16'h9f4;
17'h4b16:	data_out=16'h88b7;
17'h4b17:	data_out=16'h890c;
17'h4b18:	data_out=16'h8746;
17'h4b19:	data_out=16'ha00;
17'h4b1a:	data_out=16'h9fc;
17'h4b1b:	data_out=16'h89e0;
17'h4b1c:	data_out=16'h8693;
17'h4b1d:	data_out=16'h9fb;
17'h4b1e:	data_out=16'h8941;
17'h4b1f:	data_out=16'h4a7;
17'h4b20:	data_out=16'h9da;
17'h4b21:	data_out=16'h3d2;
17'h4b22:	data_out=16'h89de;
17'h4b23:	data_out=16'h89ef;
17'h4b24:	data_out=16'h89f0;
17'h4b25:	data_out=16'h89eb;
17'h4b26:	data_out=16'h89e2;
17'h4b27:	data_out=16'h9a3;
17'h4b28:	data_out=16'h401;
17'h4b29:	data_out=16'h9f6;
17'h4b2a:	data_out=16'h889f;
17'h4b2b:	data_out=16'ha00;
17'h4b2c:	data_out=16'h8430;
17'h4b2d:	data_out=16'h8964;
17'h4b2e:	data_out=16'h8837;
17'h4b2f:	data_out=16'ha00;
17'h4b30:	data_out=16'h9d0;
17'h4b31:	data_out=16'h9f7;
17'h4b32:	data_out=16'h9d3;
17'h4b33:	data_out=16'h8981;
17'h4b34:	data_out=16'ha00;
17'h4b35:	data_out=16'h9bd;
17'h4b36:	data_out=16'h8882;
17'h4b37:	data_out=16'h8987;
17'h4b38:	data_out=16'h2da;
17'h4b39:	data_out=16'h89c9;
17'h4b3a:	data_out=16'h89f5;
17'h4b3b:	data_out=16'h9f4;
17'h4b3c:	data_out=16'h892d;
17'h4b3d:	data_out=16'h9c5;
17'h4b3e:	data_out=16'h401;
17'h4b3f:	data_out=16'h9e6;
17'h4b40:	data_out=16'h9e7;
17'h4b41:	data_out=16'h89ce;
17'h4b42:	data_out=16'h89ee;
17'h4b43:	data_out=16'ha00;
17'h4b44:	data_out=16'h889;
17'h4b45:	data_out=16'h9f4;
17'h4b46:	data_out=16'h89d4;
17'h4b47:	data_out=16'h89ed;
17'h4b48:	data_out=16'h89f6;
17'h4b49:	data_out=16'h89fd;
17'h4b4a:	data_out=16'ha00;
17'h4b4b:	data_out=16'h89f6;
17'h4b4c:	data_out=16'h8a00;
17'h4b4d:	data_out=16'h89d7;
17'h4b4e:	data_out=16'ha00;
17'h4b4f:	data_out=16'h8a00;
17'h4b50:	data_out=16'h37b;
17'h4b51:	data_out=16'h89f9;
17'h4b52:	data_out=16'h89c2;
17'h4b53:	data_out=16'h9e4;
17'h4b54:	data_out=16'h9e8;
17'h4b55:	data_out=16'h8971;
17'h4b56:	data_out=16'h89fc;
17'h4b57:	data_out=16'h821a;
17'h4b58:	data_out=16'h89ef;
17'h4b59:	data_out=16'h9ba;
17'h4b5a:	data_out=16'h89d1;
17'h4b5b:	data_out=16'h9e4;
17'h4b5c:	data_out=16'h396;
17'h4b5d:	data_out=16'h8410;
17'h4b5e:	data_out=16'h5b;
17'h4b5f:	data_out=16'h85e1;
17'h4b60:	data_out=16'h898c;
17'h4b61:	data_out=16'h9d7;
17'h4b62:	data_out=16'h893d;
17'h4b63:	data_out=16'h88eb;
17'h4b64:	data_out=16'h8814;
17'h4b65:	data_out=16'h244;
17'h4b66:	data_out=16'ha00;
17'h4b67:	data_out=16'ha00;
17'h4b68:	data_out=16'h3d0;
17'h4b69:	data_out=16'h89ed;
17'h4b6a:	data_out=16'h40e;
17'h4b6b:	data_out=16'h9e5;
17'h4b6c:	data_out=16'h813d;
17'h4b6d:	data_out=16'h88fd;
17'h4b6e:	data_out=16'h40b;
17'h4b6f:	data_out=16'ha00;
17'h4b70:	data_out=16'h3f4;
17'h4b71:	data_out=16'h8850;
17'h4b72:	data_out=16'h9d1;
17'h4b73:	data_out=16'h9f3;
17'h4b74:	data_out=16'h971;
17'h4b75:	data_out=16'h89ec;
17'h4b76:	data_out=16'ha00;
17'h4b77:	data_out=16'h89f9;
17'h4b78:	data_out=16'ha00;
17'h4b79:	data_out=16'h509;
17'h4b7a:	data_out=16'h8901;
17'h4b7b:	data_out=16'h3fd;
17'h4b7c:	data_out=16'h21a;
17'h4b7d:	data_out=16'h9f3;
17'h4b7e:	data_out=16'h8a00;
17'h4b7f:	data_out=16'h9ac;
17'h4b80:	data_out=16'h9c2;
17'h4b81:	data_out=16'ha00;
17'h4b82:	data_out=16'h89ad;
17'h4b83:	data_out=16'h8966;
17'h4b84:	data_out=16'h9de;
17'h4b85:	data_out=16'h624;
17'h4b86:	data_out=16'h8a00;
17'h4b87:	data_out=16'h89f3;
17'h4b88:	data_out=16'h89c4;
17'h4b89:	data_out=16'h8a00;
17'h4b8a:	data_out=16'h9f2;
17'h4b8b:	data_out=16'h88d4;
17'h4b8c:	data_out=16'h89e3;
17'h4b8d:	data_out=16'h8a00;
17'h4b8e:	data_out=16'h5b8;
17'h4b8f:	data_out=16'h89a2;
17'h4b90:	data_out=16'h89e2;
17'h4b91:	data_out=16'h872;
17'h4b92:	data_out=16'h89ec;
17'h4b93:	data_out=16'h89b0;
17'h4b94:	data_out=16'h88ef;
17'h4b95:	data_out=16'h9f5;
17'h4b96:	data_out=16'h894a;
17'h4b97:	data_out=16'h890d;
17'h4b98:	data_out=16'h89fd;
17'h4b99:	data_out=16'ha00;
17'h4b9a:	data_out=16'h9fe;
17'h4b9b:	data_out=16'h89d8;
17'h4b9c:	data_out=16'h84d5;
17'h4b9d:	data_out=16'h9ec;
17'h4b9e:	data_out=16'h894f;
17'h4b9f:	data_out=16'h8545;
17'h4ba0:	data_out=16'h9c8;
17'h4ba1:	data_out=16'h4ef;
17'h4ba2:	data_out=16'h8998;
17'h4ba3:	data_out=16'h89e3;
17'h4ba4:	data_out=16'h89e4;
17'h4ba5:	data_out=16'h89b1;
17'h4ba6:	data_out=16'h8958;
17'h4ba7:	data_out=16'h7fd;
17'h4ba8:	data_out=16'h469;
17'h4ba9:	data_out=16'ha00;
17'h4baa:	data_out=16'h895a;
17'h4bab:	data_out=16'ha00;
17'h4bac:	data_out=16'h8910;
17'h4bad:	data_out=16'h88f9;
17'h4bae:	data_out=16'h88cd;
17'h4baf:	data_out=16'h8891;
17'h4bb0:	data_out=16'h9d4;
17'h4bb1:	data_out=16'h9f5;
17'h4bb2:	data_out=16'h9cf;
17'h4bb3:	data_out=16'h8984;
17'h4bb4:	data_out=16'ha00;
17'h4bb5:	data_out=16'h9a8;
17'h4bb6:	data_out=16'h8949;
17'h4bb7:	data_out=16'h8983;
17'h4bb8:	data_out=16'h8601;
17'h4bb9:	data_out=16'h89a4;
17'h4bba:	data_out=16'h89f0;
17'h4bbb:	data_out=16'h720;
17'h4bbc:	data_out=16'h8735;
17'h4bbd:	data_out=16'h9b9;
17'h4bbe:	data_out=16'h465;
17'h4bbf:	data_out=16'h658;
17'h4bc0:	data_out=16'h9e4;
17'h4bc1:	data_out=16'h8978;
17'h4bc2:	data_out=16'h8a00;
17'h4bc3:	data_out=16'h7c0;
17'h4bc4:	data_out=16'h8e0;
17'h4bc5:	data_out=16'h9f4;
17'h4bc6:	data_out=16'h358;
17'h4bc7:	data_out=16'h89eb;
17'h4bc8:	data_out=16'h8a00;
17'h4bc9:	data_out=16'h89d5;
17'h4bca:	data_out=16'h89cb;
17'h4bcb:	data_out=16'h8a00;
17'h4bcc:	data_out=16'h89fc;
17'h4bcd:	data_out=16'h89b9;
17'h4bce:	data_out=16'h528;
17'h4bcf:	data_out=16'h8a00;
17'h4bd0:	data_out=16'h8918;
17'h4bd1:	data_out=16'h89c3;
17'h4bd2:	data_out=16'h85b2;
17'h4bd3:	data_out=16'h88ea;
17'h4bd4:	data_out=16'h9cd;
17'h4bd5:	data_out=16'h8947;
17'h4bd6:	data_out=16'h86b1;
17'h4bd7:	data_out=16'h5a9;
17'h4bd8:	data_out=16'h89e3;
17'h4bd9:	data_out=16'h9c0;
17'h4bda:	data_out=16'h89d6;
17'h4bdb:	data_out=16'h9e7;
17'h4bdc:	data_out=16'h824a;
17'h4bdd:	data_out=16'h877d;
17'h4bde:	data_out=16'h88f3;
17'h4bdf:	data_out=16'h898b;
17'h4be0:	data_out=16'h88f2;
17'h4be1:	data_out=16'h9d6;
17'h4be2:	data_out=16'h88ab;
17'h4be3:	data_out=16'h8971;
17'h4be4:	data_out=16'h9eb;
17'h4be5:	data_out=16'h9fc;
17'h4be6:	data_out=16'ha00;
17'h4be7:	data_out=16'ha00;
17'h4be8:	data_out=16'h49b;
17'h4be9:	data_out=16'h89e3;
17'h4bea:	data_out=16'h646;
17'h4beb:	data_out=16'h9d7;
17'h4bec:	data_out=16'h9ee;
17'h4bed:	data_out=16'h8974;
17'h4bee:	data_out=16'h641;
17'h4bef:	data_out=16'ha00;
17'h4bf0:	data_out=16'h5ee;
17'h4bf1:	data_out=16'h8977;
17'h4bf2:	data_out=16'h9db;
17'h4bf3:	data_out=16'ha00;
17'h4bf4:	data_out=16'h94c;
17'h4bf5:	data_out=16'h89e7;
17'h4bf6:	data_out=16'ha00;
17'h4bf7:	data_out=16'h89fe;
17'h4bf8:	data_out=16'ha00;
17'h4bf9:	data_out=16'h3d3;
17'h4bfa:	data_out=16'h8938;
17'h4bfb:	data_out=16'h45e;
17'h4bfc:	data_out=16'h87c3;
17'h4bfd:	data_out=16'h543;
17'h4bfe:	data_out=16'h89f5;
17'h4bff:	data_out=16'h888c;
17'h4c00:	data_out=16'h993;
17'h4c01:	data_out=16'h9f7;
17'h4c02:	data_out=16'h89b0;
17'h4c03:	data_out=16'h894e;
17'h4c04:	data_out=16'h9bf;
17'h4c05:	data_out=16'h3d6;
17'h4c06:	data_out=16'h89f6;
17'h4c07:	data_out=16'h8a00;
17'h4c08:	data_out=16'h89d9;
17'h4c09:	data_out=16'h89f7;
17'h4c0a:	data_out=16'h9ed;
17'h4c0b:	data_out=16'h37;
17'h4c0c:	data_out=16'h89f9;
17'h4c0d:	data_out=16'h8a00;
17'h4c0e:	data_out=16'h22f;
17'h4c0f:	data_out=16'h89b3;
17'h4c10:	data_out=16'h895e;
17'h4c11:	data_out=16'h81c;
17'h4c12:	data_out=16'h89fc;
17'h4c13:	data_out=16'h8980;
17'h4c14:	data_out=16'h88cb;
17'h4c15:	data_out=16'h38a;
17'h4c16:	data_out=16'h899d;
17'h4c17:	data_out=16'h8927;
17'h4c18:	data_out=16'h89ff;
17'h4c19:	data_out=16'ha00;
17'h4c1a:	data_out=16'h9f1;
17'h4c1b:	data_out=16'h89ca;
17'h4c1c:	data_out=16'h89a2;
17'h4c1d:	data_out=16'h9ec;
17'h4c1e:	data_out=16'h8960;
17'h4c1f:	data_out=16'h85d0;
17'h4c20:	data_out=16'h9a8;
17'h4c21:	data_out=16'h15a;
17'h4c22:	data_out=16'h8904;
17'h4c23:	data_out=16'h89d8;
17'h4c24:	data_out=16'h89da;
17'h4c25:	data_out=16'h8961;
17'h4c26:	data_out=16'h8947;
17'h4c27:	data_out=16'h661;
17'h4c28:	data_out=16'hf2;
17'h4c29:	data_out=16'ha00;
17'h4c2a:	data_out=16'h8958;
17'h4c2b:	data_out=16'ha00;
17'h4c2c:	data_out=16'h8970;
17'h4c2d:	data_out=16'h8710;
17'h4c2e:	data_out=16'h88a5;
17'h4c2f:	data_out=16'h8957;
17'h4c30:	data_out=16'h9db;
17'h4c31:	data_out=16'h9d3;
17'h4c32:	data_out=16'h9e3;
17'h4c33:	data_out=16'h8985;
17'h4c34:	data_out=16'ha00;
17'h4c35:	data_out=16'h81a;
17'h4c36:	data_out=16'h8986;
17'h4c37:	data_out=16'h8983;
17'h4c38:	data_out=16'h89ed;
17'h4c39:	data_out=16'h89ab;
17'h4c3a:	data_out=16'h89da;
17'h4c3b:	data_out=16'h3bd;
17'h4c3c:	data_out=16'h862a;
17'h4c3d:	data_out=16'h98c;
17'h4c3e:	data_out=16'hef;
17'h4c3f:	data_out=16'h41e;
17'h4c40:	data_out=16'h9d8;
17'h4c41:	data_out=16'h8959;
17'h4c42:	data_out=16'h8a00;
17'h4c43:	data_out=16'ha00;
17'h4c44:	data_out=16'h709;
17'h4c45:	data_out=16'h275;
17'h4c46:	data_out=16'h703;
17'h4c47:	data_out=16'h89e1;
17'h4c48:	data_out=16'h89fd;
17'h4c49:	data_out=16'h896a;
17'h4c4a:	data_out=16'h89c1;
17'h4c4b:	data_out=16'h8a00;
17'h4c4c:	data_out=16'h89ea;
17'h4c4d:	data_out=16'h8906;
17'h4c4e:	data_out=16'h8185;
17'h4c4f:	data_out=16'h89f0;
17'h4c50:	data_out=16'h8872;
17'h4c51:	data_out=16'h89fa;
17'h4c52:	data_out=16'h81b4;
17'h4c53:	data_out=16'h89d6;
17'h4c54:	data_out=16'h192;
17'h4c55:	data_out=16'h892f;
17'h4c56:	data_out=16'h890b;
17'h4c57:	data_out=16'h8233;
17'h4c58:	data_out=16'h89fd;
17'h4c59:	data_out=16'h9c0;
17'h4c5a:	data_out=16'h89e9;
17'h4c5b:	data_out=16'h9df;
17'h4c5c:	data_out=16'h89fd;
17'h4c5d:	data_out=16'h881b;
17'h4c5e:	data_out=16'h8906;
17'h4c5f:	data_out=16'h89e4;
17'h4c60:	data_out=16'h88f8;
17'h4c61:	data_out=16'h9cb;
17'h4c62:	data_out=16'h87e6;
17'h4c63:	data_out=16'h8979;
17'h4c64:	data_out=16'h9e2;
17'h4c65:	data_out=16'ha00;
17'h4c66:	data_out=16'ha00;
17'h4c67:	data_out=16'ha00;
17'h4c68:	data_out=16'h10b;
17'h4c69:	data_out=16'h89f8;
17'h4c6a:	data_out=16'h2bd;
17'h4c6b:	data_out=16'h9b8;
17'h4c6c:	data_out=16'h84ac;
17'h4c6d:	data_out=16'h8979;
17'h4c6e:	data_out=16'h2ba;
17'h4c6f:	data_out=16'ha00;
17'h4c70:	data_out=16'h26c;
17'h4c71:	data_out=16'h8990;
17'h4c72:	data_out=16'h9df;
17'h4c73:	data_out=16'ha00;
17'h4c74:	data_out=16'h8ed;
17'h4c75:	data_out=16'h89ff;
17'h4c76:	data_out=16'ha00;
17'h4c77:	data_out=16'h89f1;
17'h4c78:	data_out=16'ha00;
17'h4c79:	data_out=16'h156;
17'h4c7a:	data_out=16'h894e;
17'h4c7b:	data_out=16'he8;
17'h4c7c:	data_out=16'h89fe;
17'h4c7d:	data_out=16'h80a6;
17'h4c7e:	data_out=16'h89e0;
17'h4c7f:	data_out=16'h88c7;
17'h4c80:	data_out=16'h859;
17'h4c81:	data_out=16'ha00;
17'h4c82:	data_out=16'h89b2;
17'h4c83:	data_out=16'h886c;
17'h4c84:	data_out=16'h9cd;
17'h4c85:	data_out=16'ha00;
17'h4c86:	data_out=16'h89f2;
17'h4c87:	data_out=16'h8a00;
17'h4c88:	data_out=16'h89cb;
17'h4c89:	data_out=16'h89f4;
17'h4c8a:	data_out=16'ha00;
17'h4c8b:	data_out=16'h9f5;
17'h4c8c:	data_out=16'h89fb;
17'h4c8d:	data_out=16'h8a00;
17'h4c8e:	data_out=16'h8875;
17'h4c8f:	data_out=16'h89a7;
17'h4c90:	data_out=16'h8911;
17'h4c91:	data_out=16'h951;
17'h4c92:	data_out=16'h89ff;
17'h4c93:	data_out=16'h8815;
17'h4c94:	data_out=16'h86da;
17'h4c95:	data_out=16'h80e0;
17'h4c96:	data_out=16'h88f8;
17'h4c97:	data_out=16'h87a2;
17'h4c98:	data_out=16'h8a00;
17'h4c99:	data_out=16'ha00;
17'h4c9a:	data_out=16'ha00;
17'h4c9b:	data_out=16'h8953;
17'h4c9c:	data_out=16'h8925;
17'h4c9d:	data_out=16'h9ed;
17'h4c9e:	data_out=16'h886c;
17'h4c9f:	data_out=16'h8542;
17'h4ca0:	data_out=16'h915;
17'h4ca1:	data_out=16'h89a5;
17'h4ca2:	data_out=16'h8967;
17'h4ca3:	data_out=16'h89ed;
17'h4ca4:	data_out=16'h89ed;
17'h4ca5:	data_out=16'h8950;
17'h4ca6:	data_out=16'h87e7;
17'h4ca7:	data_out=16'h811;
17'h4ca8:	data_out=16'h89a9;
17'h4ca9:	data_out=16'ha00;
17'h4caa:	data_out=16'h8876;
17'h4cab:	data_out=16'ha00;
17'h4cac:	data_out=16'h88a3;
17'h4cad:	data_out=16'h8561;
17'h4cae:	data_out=16'h87d6;
17'h4caf:	data_out=16'h891d;
17'h4cb0:	data_out=16'h9ba;
17'h4cb1:	data_out=16'h9e9;
17'h4cb2:	data_out=16'ha00;
17'h4cb3:	data_out=16'h8924;
17'h4cb4:	data_out=16'ha00;
17'h4cb5:	data_out=16'h9ad;
17'h4cb6:	data_out=16'h88ec;
17'h4cb7:	data_out=16'h8903;
17'h4cb8:	data_out=16'h89f5;
17'h4cb9:	data_out=16'h898a;
17'h4cba:	data_out=16'h89db;
17'h4cbb:	data_out=16'h619;
17'h4cbc:	data_out=16'h81a0;
17'h4cbd:	data_out=16'h8a4;
17'h4cbe:	data_out=16'h89a8;
17'h4cbf:	data_out=16'ha00;
17'h4cc0:	data_out=16'ha00;
17'h4cc1:	data_out=16'h88bf;
17'h4cc2:	data_out=16'h8a00;
17'h4cc3:	data_out=16'ha00;
17'h4cc4:	data_out=16'h9c9;
17'h4cc5:	data_out=16'h8102;
17'h4cc6:	data_out=16'h8eb;
17'h4cc7:	data_out=16'h89e6;
17'h4cc8:	data_out=16'h89fb;
17'h4cc9:	data_out=16'h894b;
17'h4cca:	data_out=16'h8996;
17'h4ccb:	data_out=16'h8a00;
17'h4ccc:	data_out=16'h89ff;
17'h4ccd:	data_out=16'h89bb;
17'h4cce:	data_out=16'h8729;
17'h4ccf:	data_out=16'h89f6;
17'h4cd0:	data_out=16'h88ba;
17'h4cd1:	data_out=16'h89fc;
17'h4cd2:	data_out=16'h375;
17'h4cd3:	data_out=16'h897c;
17'h4cd4:	data_out=16'h87ee;
17'h4cd5:	data_out=16'h87cb;
17'h4cd6:	data_out=16'h80da;
17'h4cd7:	data_out=16'h83a9;
17'h4cd8:	data_out=16'h89f2;
17'h4cd9:	data_out=16'h9e2;
17'h4cda:	data_out=16'h89e1;
17'h4cdb:	data_out=16'h9ec;
17'h4cdc:	data_out=16'h89ad;
17'h4cdd:	data_out=16'h886a;
17'h4cde:	data_out=16'h8869;
17'h4cdf:	data_out=16'h89e3;
17'h4ce0:	data_out=16'h8556;
17'h4ce1:	data_out=16'h9f5;
17'h4ce2:	data_out=16'h8501;
17'h4ce3:	data_out=16'h88f0;
17'h4ce4:	data_out=16'h9c7;
17'h4ce5:	data_out=16'ha00;
17'h4ce6:	data_out=16'ha00;
17'h4ce7:	data_out=16'ha00;
17'h4ce8:	data_out=16'h89b4;
17'h4ce9:	data_out=16'h8a00;
17'h4cea:	data_out=16'h87ba;
17'h4ceb:	data_out=16'h9af;
17'h4cec:	data_out=16'h8334;
17'h4ced:	data_out=16'h88f6;
17'h4cee:	data_out=16'h87be;
17'h4cef:	data_out=16'ha00;
17'h4cf0:	data_out=16'h8821;
17'h4cf1:	data_out=16'h8978;
17'h4cf2:	data_out=16'h9fc;
17'h4cf3:	data_out=16'ha00;
17'h4cf4:	data_out=16'h840;
17'h4cf5:	data_out=16'h89de;
17'h4cf6:	data_out=16'ha00;
17'h4cf7:	data_out=16'h89f4;
17'h4cf8:	data_out=16'ha00;
17'h4cf9:	data_out=16'h8536;
17'h4cfa:	data_out=16'h8824;
17'h4cfb:	data_out=16'h89a8;
17'h4cfc:	data_out=16'h89fd;
17'h4cfd:	data_out=16'h8427;
17'h4cfe:	data_out=16'h89d6;
17'h4cff:	data_out=16'h89f4;
17'h4d00:	data_out=16'h895c;
17'h4d01:	data_out=16'h9ff;
17'h4d02:	data_out=16'h897e;
17'h4d03:	data_out=16'h8888;
17'h4d04:	data_out=16'h9ee;
17'h4d05:	data_out=16'ha00;
17'h4d06:	data_out=16'h89be;
17'h4d07:	data_out=16'h89f9;
17'h4d08:	data_out=16'h89dc;
17'h4d09:	data_out=16'h897d;
17'h4d0a:	data_out=16'ha00;
17'h4d0b:	data_out=16'h8434;
17'h4d0c:	data_out=16'h89da;
17'h4d0d:	data_out=16'h8a00;
17'h4d0e:	data_out=16'h875a;
17'h4d0f:	data_out=16'h894a;
17'h4d10:	data_out=16'h88de;
17'h4d11:	data_out=16'h740;
17'h4d12:	data_out=16'h8a00;
17'h4d13:	data_out=16'h85a0;
17'h4d14:	data_out=16'h8682;
17'h4d15:	data_out=16'h88b2;
17'h4d16:	data_out=16'h88a9;
17'h4d17:	data_out=16'h86fa;
17'h4d18:	data_out=16'h8a00;
17'h4d19:	data_out=16'ha00;
17'h4d1a:	data_out=16'ha00;
17'h4d1b:	data_out=16'h8905;
17'h4d1c:	data_out=16'h899f;
17'h4d1d:	data_out=16'h9d7;
17'h4d1e:	data_out=16'h8837;
17'h4d1f:	data_out=16'h801f;
17'h4d20:	data_out=16'h8784;
17'h4d21:	data_out=16'h8860;
17'h4d22:	data_out=16'h8982;
17'h4d23:	data_out=16'h89de;
17'h4d24:	data_out=16'h89de;
17'h4d25:	data_out=16'h88c6;
17'h4d26:	data_out=16'h888f;
17'h4d27:	data_out=16'h8372;
17'h4d28:	data_out=16'h88a7;
17'h4d29:	data_out=16'ha00;
17'h4d2a:	data_out=16'h87ce;
17'h4d2b:	data_out=16'h9ee;
17'h4d2c:	data_out=16'h888c;
17'h4d2d:	data_out=16'h89d1;
17'h4d2e:	data_out=16'h8671;
17'h4d2f:	data_out=16'h8942;
17'h4d30:	data_out=16'h9f1;
17'h4d31:	data_out=16'h9ff;
17'h4d32:	data_out=16'ha00;
17'h4d33:	data_out=16'h893a;
17'h4d34:	data_out=16'h9ee;
17'h4d35:	data_out=16'h39;
17'h4d36:	data_out=16'h890e;
17'h4d37:	data_out=16'h8870;
17'h4d38:	data_out=16'h89fb;
17'h4d39:	data_out=16'h898a;
17'h4d3a:	data_out=16'h8987;
17'h4d3b:	data_out=16'h644;
17'h4d3c:	data_out=16'h1d8;
17'h4d3d:	data_out=16'h85e5;
17'h4d3e:	data_out=16'h88a1;
17'h4d3f:	data_out=16'ha00;
17'h4d40:	data_out=16'ha00;
17'h4d41:	data_out=16'h89c6;
17'h4d42:	data_out=16'h8a00;
17'h4d43:	data_out=16'ha00;
17'h4d44:	data_out=16'h9e6;
17'h4d45:	data_out=16'h88a1;
17'h4d46:	data_out=16'h8954;
17'h4d47:	data_out=16'h89de;
17'h4d48:	data_out=16'h89df;
17'h4d49:	data_out=16'h8910;
17'h4d4a:	data_out=16'h8950;
17'h4d4b:	data_out=16'h8a00;
17'h4d4c:	data_out=16'h89f8;
17'h4d4d:	data_out=16'h89b1;
17'h4d4e:	data_out=16'h8982;
17'h4d4f:	data_out=16'h89ee;
17'h4d50:	data_out=16'h8882;
17'h4d51:	data_out=16'h89bd;
17'h4d52:	data_out=16'h4ee;
17'h4d53:	data_out=16'h8909;
17'h4d54:	data_out=16'h88ad;
17'h4d55:	data_out=16'h85ef;
17'h4d56:	data_out=16'h87ff;
17'h4d57:	data_out=16'h8528;
17'h4d58:	data_out=16'h89f2;
17'h4d59:	data_out=16'ha00;
17'h4d5a:	data_out=16'h89be;
17'h4d5b:	data_out=16'h9f5;
17'h4d5c:	data_out=16'h8971;
17'h4d5d:	data_out=16'h88ad;
17'h4d5e:	data_out=16'h87f3;
17'h4d5f:	data_out=16'h89dd;
17'h4d60:	data_out=16'h87ed;
17'h4d61:	data_out=16'ha00;
17'h4d62:	data_out=16'h8341;
17'h4d63:	data_out=16'h88eb;
17'h4d64:	data_out=16'h994;
17'h4d65:	data_out=16'ha00;
17'h4d66:	data_out=16'ha00;
17'h4d67:	data_out=16'ha00;
17'h4d68:	data_out=16'h88ac;
17'h4d69:	data_out=16'h89fe;
17'h4d6a:	data_out=16'h86b2;
17'h4d6b:	data_out=16'h8fc;
17'h4d6c:	data_out=16'h883b;
17'h4d6d:	data_out=16'h88fb;
17'h4d6e:	data_out=16'h86b3;
17'h4d6f:	data_out=16'ha00;
17'h4d70:	data_out=16'h8708;
17'h4d71:	data_out=16'h88e0;
17'h4d72:	data_out=16'ha00;
17'h4d73:	data_out=16'ha00;
17'h4d74:	data_out=16'h869;
17'h4d75:	data_out=16'h8965;
17'h4d76:	data_out=16'h9ea;
17'h4d77:	data_out=16'h89d1;
17'h4d78:	data_out=16'ha00;
17'h4d79:	data_out=16'h89f8;
17'h4d7a:	data_out=16'h8813;
17'h4d7b:	data_out=16'h88a3;
17'h4d7c:	data_out=16'h89fe;
17'h4d7d:	data_out=16'h8392;
17'h4d7e:	data_out=16'h89cd;
17'h4d7f:	data_out=16'h89e5;
17'h4d80:	data_out=16'h89ea;
17'h4d81:	data_out=16'h9fa;
17'h4d82:	data_out=16'h8999;
17'h4d83:	data_out=16'h898d;
17'h4d84:	data_out=16'h9fe;
17'h4d85:	data_out=16'ha00;
17'h4d86:	data_out=16'h89a7;
17'h4d87:	data_out=16'h89ed;
17'h4d88:	data_out=16'h89de;
17'h4d89:	data_out=16'h892e;
17'h4d8a:	data_out=16'ha00;
17'h4d8b:	data_out=16'h8839;
17'h4d8c:	data_out=16'h89eb;
17'h4d8d:	data_out=16'h8a00;
17'h4d8e:	data_out=16'h212;
17'h4d8f:	data_out=16'h8971;
17'h4d90:	data_out=16'h8963;
17'h4d91:	data_out=16'h951;
17'h4d92:	data_out=16'h8a00;
17'h4d93:	data_out=16'h839f;
17'h4d94:	data_out=16'h886f;
17'h4d95:	data_out=16'h898d;
17'h4d96:	data_out=16'h8929;
17'h4d97:	data_out=16'h888f;
17'h4d98:	data_out=16'h8a00;
17'h4d99:	data_out=16'ha00;
17'h4d9a:	data_out=16'ha00;
17'h4d9b:	data_out=16'h893b;
17'h4d9c:	data_out=16'h89db;
17'h4d9d:	data_out=16'h9df;
17'h4d9e:	data_out=16'h890f;
17'h4d9f:	data_out=16'h274;
17'h4da0:	data_out=16'h88d0;
17'h4da1:	data_out=16'h137;
17'h4da2:	data_out=16'h8977;
17'h4da3:	data_out=16'h964;
17'h4da4:	data_out=16'h924;
17'h4da5:	data_out=16'h880c;
17'h4da6:	data_out=16'h8984;
17'h4da7:	data_out=16'h80de;
17'h4da8:	data_out=16'h173;
17'h4da9:	data_out=16'h9e4;
17'h4daa:	data_out=16'h8861;
17'h4dab:	data_out=16'h9fe;
17'h4dac:	data_out=16'h8926;
17'h4dad:	data_out=16'h89fe;
17'h4dae:	data_out=16'h85ac;
17'h4daf:	data_out=16'h8944;
17'h4db0:	data_out=16'h9f7;
17'h4db1:	data_out=16'ha00;
17'h4db2:	data_out=16'ha00;
17'h4db3:	data_out=16'h8968;
17'h4db4:	data_out=16'h9f0;
17'h4db5:	data_out=16'h4ed;
17'h4db6:	data_out=16'h8966;
17'h4db7:	data_out=16'h88a2;
17'h4db8:	data_out=16'h89ba;
17'h4db9:	data_out=16'h89a3;
17'h4dba:	data_out=16'h896e;
17'h4dbb:	data_out=16'h9b4;
17'h4dbc:	data_out=16'h278;
17'h4dbd:	data_out=16'h88aa;
17'h4dbe:	data_out=16'h180;
17'h4dbf:	data_out=16'ha00;
17'h4dc0:	data_out=16'ha00;
17'h4dc1:	data_out=16'h89dd;
17'h4dc2:	data_out=16'h8a00;
17'h4dc3:	data_out=16'ha00;
17'h4dc4:	data_out=16'ha00;
17'h4dc5:	data_out=16'h8987;
17'h4dc6:	data_out=16'h89f9;
17'h4dc7:	data_out=16'h89d3;
17'h4dc8:	data_out=16'h89bd;
17'h4dc9:	data_out=16'h892f;
17'h4dca:	data_out=16'h8928;
17'h4dcb:	data_out=16'h8a00;
17'h4dcc:	data_out=16'h89ee;
17'h4dcd:	data_out=16'h89a3;
17'h4dce:	data_out=16'h89d7;
17'h4dcf:	data_out=16'h89df;
17'h4dd0:	data_out=16'h892b;
17'h4dd1:	data_out=16'h89d5;
17'h4dd2:	data_out=16'h74b;
17'h4dd3:	data_out=16'h88b4;
17'h4dd4:	data_out=16'h891e;
17'h4dd5:	data_out=16'h868b;
17'h4dd6:	data_out=16'h892b;
17'h4dd7:	data_out=16'h873c;
17'h4dd8:	data_out=16'h89ef;
17'h4dd9:	data_out=16'ha00;
17'h4dda:	data_out=16'h89b7;
17'h4ddb:	data_out=16'ha00;
17'h4ddc:	data_out=16'h895b;
17'h4ddd:	data_out=16'h8928;
17'h4dde:	data_out=16'h8839;
17'h4ddf:	data_out=16'h89e0;
17'h4de0:	data_out=16'h8943;
17'h4de1:	data_out=16'ha00;
17'h4de2:	data_out=16'h8356;
17'h4de3:	data_out=16'h893e;
17'h4de4:	data_out=16'h6f1;
17'h4de5:	data_out=16'ha00;
17'h4de6:	data_out=16'ha00;
17'h4de7:	data_out=16'ha00;
17'h4de8:	data_out=16'h108;
17'h4de9:	data_out=16'h8a00;
17'h4dea:	data_out=16'h2a0;
17'h4deb:	data_out=16'ha00;
17'h4dec:	data_out=16'h89db;
17'h4ded:	data_out=16'h8945;
17'h4dee:	data_out=16'h2a1;
17'h4def:	data_out=16'ha00;
17'h4df0:	data_out=16'h261;
17'h4df1:	data_out=16'h892c;
17'h4df2:	data_out=16'ha00;
17'h4df3:	data_out=16'ha00;
17'h4df4:	data_out=16'h98b;
17'h4df5:	data_out=16'h247;
17'h4df6:	data_out=16'h9e0;
17'h4df7:	data_out=16'h89af;
17'h4df8:	data_out=16'ha00;
17'h4df9:	data_out=16'h8a00;
17'h4dfa:	data_out=16'h88fe;
17'h4dfb:	data_out=16'h182;
17'h4dfc:	data_out=16'h8a00;
17'h4dfd:	data_out=16'h82be;
17'h4dfe:	data_out=16'h89ae;
17'h4dff:	data_out=16'h89d3;
17'h4e00:	data_out=16'h8a00;
17'h4e01:	data_out=16'h9fe;
17'h4e02:	data_out=16'h8939;
17'h4e03:	data_out=16'h89a8;
17'h4e04:	data_out=16'h9ff;
17'h4e05:	data_out=16'ha00;
17'h4e06:	data_out=16'h89ad;
17'h4e07:	data_out=16'h158;
17'h4e08:	data_out=16'h89ef;
17'h4e09:	data_out=16'h889c;
17'h4e0a:	data_out=16'ha00;
17'h4e0b:	data_out=16'h8989;
17'h4e0c:	data_out=16'h89f1;
17'h4e0d:	data_out=16'h8a00;
17'h4e0e:	data_out=16'h9ff;
17'h4e0f:	data_out=16'h8933;
17'h4e10:	data_out=16'h899a;
17'h4e11:	data_out=16'ha00;
17'h4e12:	data_out=16'h8a00;
17'h4e13:	data_out=16'h83ac;
17'h4e14:	data_out=16'h8957;
17'h4e15:	data_out=16'h89d8;
17'h4e16:	data_out=16'h89d3;
17'h4e17:	data_out=16'h894e;
17'h4e18:	data_out=16'h8a00;
17'h4e19:	data_out=16'ha00;
17'h4e1a:	data_out=16'ha00;
17'h4e1b:	data_out=16'h8956;
17'h4e1c:	data_out=16'h89fe;
17'h4e1d:	data_out=16'h9e8;
17'h4e1e:	data_out=16'h8959;
17'h4e1f:	data_out=16'h15f;
17'h4e20:	data_out=16'h85fd;
17'h4e21:	data_out=16'h9ff;
17'h4e22:	data_out=16'h86a0;
17'h4e23:	data_out=16'h9e6;
17'h4e24:	data_out=16'h9e4;
17'h4e25:	data_out=16'h12b;
17'h4e26:	data_out=16'h8916;
17'h4e27:	data_out=16'ha00;
17'h4e28:	data_out=16'h9ff;
17'h4e29:	data_out=16'h9e7;
17'h4e2a:	data_out=16'h8766;
17'h4e2b:	data_out=16'h9ff;
17'h4e2c:	data_out=16'h89d9;
17'h4e2d:	data_out=16'h89bf;
17'h4e2e:	data_out=16'h8269;
17'h4e2f:	data_out=16'h8975;
17'h4e30:	data_out=16'ha00;
17'h4e31:	data_out=16'ha00;
17'h4e32:	data_out=16'ha00;
17'h4e33:	data_out=16'h899f;
17'h4e34:	data_out=16'h9e2;
17'h4e35:	data_out=16'ha00;
17'h4e36:	data_out=16'h893f;
17'h4e37:	data_out=16'h8689;
17'h4e38:	data_out=16'h88f9;
17'h4e39:	data_out=16'h89d3;
17'h4e3a:	data_out=16'h891c;
17'h4e3b:	data_out=16'h9fe;
17'h4e3c:	data_out=16'h355;
17'h4e3d:	data_out=16'h85ad;
17'h4e3e:	data_out=16'h9ff;
17'h4e3f:	data_out=16'ha00;
17'h4e40:	data_out=16'ha00;
17'h4e41:	data_out=16'h8a00;
17'h4e42:	data_out=16'h8a00;
17'h4e43:	data_out=16'ha00;
17'h4e44:	data_out=16'ha00;
17'h4e45:	data_out=16'h89dc;
17'h4e46:	data_out=16'h89b0;
17'h4e47:	data_out=16'h89c4;
17'h4e48:	data_out=16'h89b4;
17'h4e49:	data_out=16'h1fb;
17'h4e4a:	data_out=16'h855c;
17'h4e4b:	data_out=16'h8a00;
17'h4e4c:	data_out=16'h8930;
17'h4e4d:	data_out=16'h8674;
17'h4e4e:	data_out=16'h89dc;
17'h4e4f:	data_out=16'h86fb;
17'h4e50:	data_out=16'h898e;
17'h4e51:	data_out=16'h89f3;
17'h4e52:	data_out=16'h9c8;
17'h4e53:	data_out=16'h86ee;
17'h4e54:	data_out=16'h88cd;
17'h4e55:	data_out=16'h8848;
17'h4e56:	data_out=16'h256;
17'h4e57:	data_out=16'h9ea;
17'h4e58:	data_out=16'h89f4;
17'h4e59:	data_out=16'ha00;
17'h4e5a:	data_out=16'h89d6;
17'h4e5b:	data_out=16'ha00;
17'h4e5c:	data_out=16'h8989;
17'h4e5d:	data_out=16'h87e2;
17'h4e5e:	data_out=16'h8840;
17'h4e5f:	data_out=16'h89db;
17'h4e60:	data_out=16'h88ea;
17'h4e61:	data_out=16'ha00;
17'h4e62:	data_out=16'h852e;
17'h4e63:	data_out=16'h897d;
17'h4e64:	data_out=16'h8000;
17'h4e65:	data_out=16'ha00;
17'h4e66:	data_out=16'ha00;
17'h4e67:	data_out=16'ha00;
17'h4e68:	data_out=16'h9ff;
17'h4e69:	data_out=16'h8a00;
17'h4e6a:	data_out=16'h9fe;
17'h4e6b:	data_out=16'ha00;
17'h4e6c:	data_out=16'h89f8;
17'h4e6d:	data_out=16'h8981;
17'h4e6e:	data_out=16'h9fe;
17'h4e6f:	data_out=16'ha00;
17'h4e70:	data_out=16'h9fe;
17'h4e71:	data_out=16'h88f5;
17'h4e72:	data_out=16'ha00;
17'h4e73:	data_out=16'ha00;
17'h4e74:	data_out=16'h9e2;
17'h4e75:	data_out=16'h9eb;
17'h4e76:	data_out=16'h9f7;
17'h4e77:	data_out=16'h8978;
17'h4e78:	data_out=16'ha00;
17'h4e79:	data_out=16'h8a00;
17'h4e7a:	data_out=16'h8965;
17'h4e7b:	data_out=16'h9ff;
17'h4e7c:	data_out=16'h8a00;
17'h4e7d:	data_out=16'h807a;
17'h4e7e:	data_out=16'h8988;
17'h4e7f:	data_out=16'h89e5;
17'h4e80:	data_out=16'h89f5;
17'h4e81:	data_out=16'h9ff;
17'h4e82:	data_out=16'h89b1;
17'h4e83:	data_out=16'h89ff;
17'h4e84:	data_out=16'h9ff;
17'h4e85:	data_out=16'ha00;
17'h4e86:	data_out=16'h89f1;
17'h4e87:	data_out=16'h9c2;
17'h4e88:	data_out=16'h8a00;
17'h4e89:	data_out=16'h23e;
17'h4e8a:	data_out=16'ha00;
17'h4e8b:	data_out=16'h899b;
17'h4e8c:	data_out=16'h80b8;
17'h4e8d:	data_out=16'h8a00;
17'h4e8e:	data_out=16'h9ff;
17'h4e8f:	data_out=16'h8996;
17'h4e90:	data_out=16'h89b3;
17'h4e91:	data_out=16'ha00;
17'h4e92:	data_out=16'h8a00;
17'h4e93:	data_out=16'h85b0;
17'h4e94:	data_out=16'h89ea;
17'h4e95:	data_out=16'h89e8;
17'h4e96:	data_out=16'h89e8;
17'h4e97:	data_out=16'h89ff;
17'h4e98:	data_out=16'h8a00;
17'h4e99:	data_out=16'ha00;
17'h4e9a:	data_out=16'ha00;
17'h4e9b:	data_out=16'h89c3;
17'h4e9c:	data_out=16'h8a00;
17'h4e9d:	data_out=16'ha00;
17'h4e9e:	data_out=16'h89cd;
17'h4e9f:	data_out=16'h85f4;
17'h4ea0:	data_out=16'h8858;
17'h4ea1:	data_out=16'h9ff;
17'h4ea2:	data_out=16'h495;
17'h4ea3:	data_out=16'ha00;
17'h4ea4:	data_out=16'ha00;
17'h4ea5:	data_out=16'ha00;
17'h4ea6:	data_out=16'h8760;
17'h4ea7:	data_out=16'ha00;
17'h4ea8:	data_out=16'h9ff;
17'h4ea9:	data_out=16'h822;
17'h4eaa:	data_out=16'h86f8;
17'h4eab:	data_out=16'h827;
17'h4eac:	data_out=16'h89ee;
17'h4ead:	data_out=16'h896c;
17'h4eae:	data_out=16'h8470;
17'h4eaf:	data_out=16'h89cd;
17'h4eb0:	data_out=16'ha00;
17'h4eb1:	data_out=16'ha00;
17'h4eb2:	data_out=16'ha00;
17'h4eb3:	data_out=16'h8a00;
17'h4eb4:	data_out=16'h9b9;
17'h4eb5:	data_out=16'ha00;
17'h4eb6:	data_out=16'h89b5;
17'h4eb7:	data_out=16'h3a4;
17'h4eb8:	data_out=16'h88aa;
17'h4eb9:	data_out=16'h8a00;
17'h4eba:	data_out=16'h8298;
17'h4ebb:	data_out=16'ha00;
17'h4ebc:	data_out=16'h8048;
17'h4ebd:	data_out=16'h8506;
17'h4ebe:	data_out=16'h9ff;
17'h4ebf:	data_out=16'ha00;
17'h4ec0:	data_out=16'ha00;
17'h4ec1:	data_out=16'h8a00;
17'h4ec2:	data_out=16'h89ff;
17'h4ec3:	data_out=16'ha00;
17'h4ec4:	data_out=16'ha00;
17'h4ec5:	data_out=16'h89e9;
17'h4ec6:	data_out=16'h8973;
17'h4ec7:	data_out=16'h89ca;
17'h4ec8:	data_out=16'h81a8;
17'h4ec9:	data_out=16'h9fb;
17'h4eca:	data_out=16'h8a3;
17'h4ecb:	data_out=16'h8a00;
17'h4ecc:	data_out=16'h9e4;
17'h4ecd:	data_out=16'h1ca;
17'h4ece:	data_out=16'h8a00;
17'h4ecf:	data_out=16'h9f3;
17'h4ed0:	data_out=16'h89de;
17'h4ed1:	data_out=16'h8a00;
17'h4ed2:	data_out=16'ha00;
17'h4ed3:	data_out=16'h88a8;
17'h4ed4:	data_out=16'h897f;
17'h4ed5:	data_out=16'h897b;
17'h4ed6:	data_out=16'h9da;
17'h4ed7:	data_out=16'h9f3;
17'h4ed8:	data_out=16'h8a00;
17'h4ed9:	data_out=16'ha00;
17'h4eda:	data_out=16'h8a00;
17'h4edb:	data_out=16'ha00;
17'h4edc:	data_out=16'h89eb;
17'h4edd:	data_out=16'h857f;
17'h4ede:	data_out=16'h88ef;
17'h4edf:	data_out=16'h89e7;
17'h4ee0:	data_out=16'h9a3;
17'h4ee1:	data_out=16'ha00;
17'h4ee2:	data_out=16'h886f;
17'h4ee3:	data_out=16'h8a00;
17'h4ee4:	data_out=16'h813f;
17'h4ee5:	data_out=16'ha00;
17'h4ee6:	data_out=16'ha00;
17'h4ee7:	data_out=16'h9f9;
17'h4ee8:	data_out=16'h9ff;
17'h4ee9:	data_out=16'h8a00;
17'h4eea:	data_out=16'h9ff;
17'h4eeb:	data_out=16'ha00;
17'h4eec:	data_out=16'h89e6;
17'h4eed:	data_out=16'h8a00;
17'h4eee:	data_out=16'h9ff;
17'h4eef:	data_out=16'ha00;
17'h4ef0:	data_out=16'h9ff;
17'h4ef1:	data_out=16'h898d;
17'h4ef2:	data_out=16'ha00;
17'h4ef3:	data_out=16'ha00;
17'h4ef4:	data_out=16'h9fd;
17'h4ef5:	data_out=16'h9ec;
17'h4ef6:	data_out=16'h9fc;
17'h4ef7:	data_out=16'h88d0;
17'h4ef8:	data_out=16'ha00;
17'h4ef9:	data_out=16'h8a00;
17'h4efa:	data_out=16'h89f7;
17'h4efb:	data_out=16'h9ff;
17'h4efc:	data_out=16'h8a00;
17'h4efd:	data_out=16'h807c;
17'h4efe:	data_out=16'h885b;
17'h4eff:	data_out=16'h89ed;
17'h4f00:	data_out=16'h89ef;
17'h4f01:	data_out=16'h9fd;
17'h4f02:	data_out=16'h89f1;
17'h4f03:	data_out=16'h89fc;
17'h4f04:	data_out=16'h9fe;
17'h4f05:	data_out=16'ha00;
17'h4f06:	data_out=16'h8259;
17'h4f07:	data_out=16'h9db;
17'h4f08:	data_out=16'h8a00;
17'h4f09:	data_out=16'h9d6;
17'h4f0a:	data_out=16'ha00;
17'h4f0b:	data_out=16'h89ee;
17'h4f0c:	data_out=16'h9ba;
17'h4f0d:	data_out=16'h8a00;
17'h4f0e:	data_out=16'h9fc;
17'h4f0f:	data_out=16'h89df;
17'h4f10:	data_out=16'h89be;
17'h4f11:	data_out=16'ha00;
17'h4f12:	data_out=16'h8a00;
17'h4f13:	data_out=16'h82ee;
17'h4f14:	data_out=16'h8a00;
17'h4f15:	data_out=16'h895e;
17'h4f16:	data_out=16'h89be;
17'h4f17:	data_out=16'h8a00;
17'h4f18:	data_out=16'h8a00;
17'h4f19:	data_out=16'ha00;
17'h4f1a:	data_out=16'ha00;
17'h4f1b:	data_out=16'h89f3;
17'h4f1c:	data_out=16'h8a00;
17'h4f1d:	data_out=16'h979;
17'h4f1e:	data_out=16'h89f8;
17'h4f1f:	data_out=16'h8289;
17'h4f20:	data_out=16'h8826;
17'h4f21:	data_out=16'h9fc;
17'h4f22:	data_out=16'h832c;
17'h4f23:	data_out=16'ha00;
17'h4f24:	data_out=16'ha00;
17'h4f25:	data_out=16'h9f1;
17'h4f26:	data_out=16'h88a6;
17'h4f27:	data_out=16'h9fb;
17'h4f28:	data_out=16'h9fb;
17'h4f29:	data_out=16'h8810;
17'h4f2a:	data_out=16'h88c8;
17'h4f2b:	data_out=16'h892f;
17'h4f2c:	data_out=16'h89c3;
17'h4f2d:	data_out=16'h89f9;
17'h4f2e:	data_out=16'h894c;
17'h4f2f:	data_out=16'h89db;
17'h4f30:	data_out=16'ha00;
17'h4f31:	data_out=16'ha00;
17'h4f32:	data_out=16'ha00;
17'h4f33:	data_out=16'h8a00;
17'h4f34:	data_out=16'h81de;
17'h4f35:	data_out=16'ha00;
17'h4f36:	data_out=16'h89e1;
17'h4f37:	data_out=16'h8691;
17'h4f38:	data_out=16'h89ed;
17'h4f39:	data_out=16'h8a00;
17'h4f3a:	data_out=16'h5c9;
17'h4f3b:	data_out=16'ha00;
17'h4f3c:	data_out=16'h878d;
17'h4f3d:	data_out=16'h874e;
17'h4f3e:	data_out=16'h9fb;
17'h4f3f:	data_out=16'ha00;
17'h4f40:	data_out=16'ha00;
17'h4f41:	data_out=16'h8a00;
17'h4f42:	data_out=16'h89fb;
17'h4f43:	data_out=16'ha00;
17'h4f44:	data_out=16'ha00;
17'h4f45:	data_out=16'h8965;
17'h4f46:	data_out=16'h89f4;
17'h4f47:	data_out=16'h89f1;
17'h4f48:	data_out=16'h66a;
17'h4f49:	data_out=16'h9ef;
17'h4f4a:	data_out=16'h9e4;
17'h4f4b:	data_out=16'h89ff;
17'h4f4c:	data_out=16'h9df;
17'h4f4d:	data_out=16'h8558;
17'h4f4e:	data_out=16'h8a00;
17'h4f4f:	data_out=16'h9e8;
17'h4f50:	data_out=16'h89d5;
17'h4f51:	data_out=16'h8a00;
17'h4f52:	data_out=16'ha00;
17'h4f53:	data_out=16'h88d7;
17'h4f54:	data_out=16'h89a1;
17'h4f55:	data_out=16'h89e0;
17'h4f56:	data_out=16'h5b6;
17'h4f57:	data_out=16'h31f;
17'h4f58:	data_out=16'h8a00;
17'h4f59:	data_out=16'ha00;
17'h4f5a:	data_out=16'h8a00;
17'h4f5b:	data_out=16'ha00;
17'h4f5c:	data_out=16'h89dc;
17'h4f5d:	data_out=16'h840d;
17'h4f5e:	data_out=16'h893b;
17'h4f5f:	data_out=16'h89ee;
17'h4f60:	data_out=16'h8599;
17'h4f61:	data_out=16'ha00;
17'h4f62:	data_out=16'h89b2;
17'h4f63:	data_out=16'h8a00;
17'h4f64:	data_out=16'h89e4;
17'h4f65:	data_out=16'ha00;
17'h4f66:	data_out=16'ha00;
17'h4f67:	data_out=16'h6bd;
17'h4f68:	data_out=16'h9fc;
17'h4f69:	data_out=16'h8a00;
17'h4f6a:	data_out=16'h9fc;
17'h4f6b:	data_out=16'ha00;
17'h4f6c:	data_out=16'h89e9;
17'h4f6d:	data_out=16'h8a00;
17'h4f6e:	data_out=16'h9fc;
17'h4f6f:	data_out=16'ha00;
17'h4f70:	data_out=16'h9fc;
17'h4f71:	data_out=16'h89d1;
17'h4f72:	data_out=16'ha00;
17'h4f73:	data_out=16'ha00;
17'h4f74:	data_out=16'ha00;
17'h4f75:	data_out=16'h9f7;
17'h4f76:	data_out=16'h85d3;
17'h4f77:	data_out=16'h859f;
17'h4f78:	data_out=16'h9fe;
17'h4f79:	data_out=16'h8a00;
17'h4f7a:	data_out=16'h8a00;
17'h4f7b:	data_out=16'h9fb;
17'h4f7c:	data_out=16'h8a00;
17'h4f7d:	data_out=16'h94b;
17'h4f7e:	data_out=16'h828a;
17'h4f7f:	data_out=16'h89ee;
17'h4f80:	data_out=16'h89f3;
17'h4f81:	data_out=16'h87e;
17'h4f82:	data_out=16'h890e;
17'h4f83:	data_out=16'h89f5;
17'h4f84:	data_out=16'h9fe;
17'h4f85:	data_out=16'ha00;
17'h4f86:	data_out=16'h74d;
17'h4f87:	data_out=16'h9fa;
17'h4f88:	data_out=16'h89f9;
17'h4f89:	data_out=16'h4fb;
17'h4f8a:	data_out=16'ha00;
17'h4f8b:	data_out=16'h89ff;
17'h4f8c:	data_out=16'h9df;
17'h4f8d:	data_out=16'h8a00;
17'h4f8e:	data_out=16'ha00;
17'h4f8f:	data_out=16'h88f9;
17'h4f90:	data_out=16'h89ee;
17'h4f91:	data_out=16'ha00;
17'h4f92:	data_out=16'h8a00;
17'h4f93:	data_out=16'h1f5;
17'h4f94:	data_out=16'h89e4;
17'h4f95:	data_out=16'h9d0;
17'h4f96:	data_out=16'ha00;
17'h4f97:	data_out=16'h89e9;
17'h4f98:	data_out=16'h89f9;
17'h4f99:	data_out=16'h9ff;
17'h4f9a:	data_out=16'ha00;
17'h4f9b:	data_out=16'h89a2;
17'h4f9c:	data_out=16'h8a00;
17'h4f9d:	data_out=16'h2fa;
17'h4f9e:	data_out=16'h89ca;
17'h4f9f:	data_out=16'h5e9;
17'h4fa0:	data_out=16'h8993;
17'h4fa1:	data_out=16'ha00;
17'h4fa2:	data_out=16'h899b;
17'h4fa3:	data_out=16'ha00;
17'h4fa4:	data_out=16'ha00;
17'h4fa5:	data_out=16'h9fa;
17'h4fa6:	data_out=16'h8912;
17'h4fa7:	data_out=16'h877d;
17'h4fa8:	data_out=16'ha00;
17'h4fa9:	data_out=16'h8054;
17'h4faa:	data_out=16'h87de;
17'h4fab:	data_out=16'h89fb;
17'h4fac:	data_out=16'ha00;
17'h4fad:	data_out=16'h89f6;
17'h4fae:	data_out=16'h8859;
17'h4faf:	data_out=16'h89c8;
17'h4fb0:	data_out=16'ha00;
17'h4fb1:	data_out=16'ha00;
17'h4fb2:	data_out=16'ha00;
17'h4fb3:	data_out=16'h8a00;
17'h4fb4:	data_out=16'h89cf;
17'h4fb5:	data_out=16'h9fe;
17'h4fb6:	data_out=16'h89bb;
17'h4fb7:	data_out=16'h84de;
17'h4fb8:	data_out=16'h8a00;
17'h4fb9:	data_out=16'h8a00;
17'h4fba:	data_out=16'h807e;
17'h4fbb:	data_out=16'ha00;
17'h4fbc:	data_out=16'h881a;
17'h4fbd:	data_out=16'h8805;
17'h4fbe:	data_out=16'ha00;
17'h4fbf:	data_out=16'ha00;
17'h4fc0:	data_out=16'ha00;
17'h4fc1:	data_out=16'h8a00;
17'h4fc2:	data_out=16'h89e0;
17'h4fc3:	data_out=16'ha00;
17'h4fc4:	data_out=16'ha00;
17'h4fc5:	data_out=16'h9fe;
17'h4fc6:	data_out=16'h89e8;
17'h4fc7:	data_out=16'h89ed;
17'h4fc8:	data_out=16'h4ed;
17'h4fc9:	data_out=16'h9fa;
17'h4fca:	data_out=16'h9ef;
17'h4fcb:	data_out=16'h89f1;
17'h4fcc:	data_out=16'h9f6;
17'h4fcd:	data_out=16'h898d;
17'h4fce:	data_out=16'h8a00;
17'h4fcf:	data_out=16'h9f1;
17'h4fd0:	data_out=16'h87cf;
17'h4fd1:	data_out=16'h852e;
17'h4fd2:	data_out=16'ha00;
17'h4fd3:	data_out=16'h8977;
17'h4fd4:	data_out=16'h89bc;
17'h4fd5:	data_out=16'h86a7;
17'h4fd6:	data_out=16'h80ee;
17'h4fd7:	data_out=16'h104;
17'h4fd8:	data_out=16'h89fe;
17'h4fd9:	data_out=16'ha00;
17'h4fda:	data_out=16'h8a00;
17'h4fdb:	data_out=16'h9f9;
17'h4fdc:	data_out=16'h89c9;
17'h4fdd:	data_out=16'h823d;
17'h4fde:	data_out=16'h8822;
17'h4fdf:	data_out=16'h89f2;
17'h4fe0:	data_out=16'h88d5;
17'h4fe1:	data_out=16'ha00;
17'h4fe2:	data_out=16'h89a5;
17'h4fe3:	data_out=16'h8a00;
17'h4fe4:	data_out=16'h8a00;
17'h4fe5:	data_out=16'ha00;
17'h4fe6:	data_out=16'ha00;
17'h4fe7:	data_out=16'h88b5;
17'h4fe8:	data_out=16'ha00;
17'h4fe9:	data_out=16'h8a00;
17'h4fea:	data_out=16'ha00;
17'h4feb:	data_out=16'ha00;
17'h4fec:	data_out=16'h89dc;
17'h4fed:	data_out=16'h8a00;
17'h4fee:	data_out=16'ha00;
17'h4fef:	data_out=16'ha00;
17'h4ff0:	data_out=16'ha00;
17'h4ff1:	data_out=16'h86ce;
17'h4ff2:	data_out=16'ha00;
17'h4ff3:	data_out=16'ha00;
17'h4ff4:	data_out=16'ha00;
17'h4ff5:	data_out=16'ha00;
17'h4ff6:	data_out=16'h89df;
17'h4ff7:	data_out=16'h85dc;
17'h4ff8:	data_out=16'ha00;
17'h4ff9:	data_out=16'h8a00;
17'h4ffa:	data_out=16'h89f8;
17'h4ffb:	data_out=16'ha00;
17'h4ffc:	data_out=16'h89fa;
17'h4ffd:	data_out=16'h9eb;
17'h4ffe:	data_out=16'h83a3;
17'h4fff:	data_out=16'h853b;
17'h5000:	data_out=16'h89d1;
17'h5001:	data_out=16'h409;
17'h5002:	data_out=16'h8933;
17'h5003:	data_out=16'h89dc;
17'h5004:	data_out=16'h9f7;
17'h5005:	data_out=16'ha00;
17'h5006:	data_out=16'h8143;
17'h5007:	data_out=16'ha00;
17'h5008:	data_out=16'h8a00;
17'h5009:	data_out=16'h868b;
17'h500a:	data_out=16'ha00;
17'h500b:	data_out=16'h8a00;
17'h500c:	data_out=16'h823e;
17'h500d:	data_out=16'h899c;
17'h500e:	data_out=16'ha00;
17'h500f:	data_out=16'h888b;
17'h5010:	data_out=16'h89f3;
17'h5011:	data_out=16'ha00;
17'h5012:	data_out=16'h89fe;
17'h5013:	data_out=16'h3fb;
17'h5014:	data_out=16'h89f4;
17'h5015:	data_out=16'ha00;
17'h5016:	data_out=16'ha00;
17'h5017:	data_out=16'h89ec;
17'h5018:	data_out=16'h89c9;
17'h5019:	data_out=16'h9cd;
17'h501a:	data_out=16'ha00;
17'h501b:	data_out=16'h89f2;
17'h501c:	data_out=16'h890c;
17'h501d:	data_out=16'h809e;
17'h501e:	data_out=16'h8981;
17'h501f:	data_out=16'h5dd;
17'h5020:	data_out=16'h8999;
17'h5021:	data_out=16'ha00;
17'h5022:	data_out=16'h89f9;
17'h5023:	data_out=16'ha00;
17'h5024:	data_out=16'ha00;
17'h5025:	data_out=16'h90d;
17'h5026:	data_out=16'h89af;
17'h5027:	data_out=16'h89c8;
17'h5028:	data_out=16'h9ff;
17'h5029:	data_out=16'h89c4;
17'h502a:	data_out=16'h88ad;
17'h502b:	data_out=16'h8a00;
17'h502c:	data_out=16'ha00;
17'h502d:	data_out=16'h89f4;
17'h502e:	data_out=16'h89d5;
17'h502f:	data_out=16'h89b2;
17'h5030:	data_out=16'ha00;
17'h5031:	data_out=16'ha00;
17'h5032:	data_out=16'ha00;
17'h5033:	data_out=16'h89ff;
17'h5034:	data_out=16'h89d6;
17'h5035:	data_out=16'h9f4;
17'h5036:	data_out=16'h89ef;
17'h5037:	data_out=16'h8905;
17'h5038:	data_out=16'h8a00;
17'h5039:	data_out=16'h8a00;
17'h503a:	data_out=16'h84ff;
17'h503b:	data_out=16'h9fe;
17'h503c:	data_out=16'h89e0;
17'h503d:	data_out=16'h9d8;
17'h503e:	data_out=16'h9ff;
17'h503f:	data_out=16'ha00;
17'h5040:	data_out=16'ha00;
17'h5041:	data_out=16'h8a00;
17'h5042:	data_out=16'h89ed;
17'h5043:	data_out=16'ha00;
17'h5044:	data_out=16'ha00;
17'h5045:	data_out=16'ha00;
17'h5046:	data_out=16'h8a00;
17'h5047:	data_out=16'h89d3;
17'h5048:	data_out=16'h89da;
17'h5049:	data_out=16'ha00;
17'h504a:	data_out=16'h1b2;
17'h504b:	data_out=16'h8a00;
17'h504c:	data_out=16'h5bd;
17'h504d:	data_out=16'h89f9;
17'h504e:	data_out=16'h8a00;
17'h504f:	data_out=16'h9e0;
17'h5050:	data_out=16'h83d7;
17'h5051:	data_out=16'h665;
17'h5052:	data_out=16'ha00;
17'h5053:	data_out=16'h89dc;
17'h5054:	data_out=16'h89fc;
17'h5055:	data_out=16'h86ff;
17'h5056:	data_out=16'h644;
17'h5057:	data_out=16'h4a7;
17'h5058:	data_out=16'h89f1;
17'h5059:	data_out=16'ha00;
17'h505a:	data_out=16'h8a00;
17'h505b:	data_out=16'h9c8;
17'h505c:	data_out=16'h89bc;
17'h505d:	data_out=16'h83fb;
17'h505e:	data_out=16'h889d;
17'h505f:	data_out=16'h89f5;
17'h5060:	data_out=16'h89bf;
17'h5061:	data_out=16'h9fd;
17'h5062:	data_out=16'h89f7;
17'h5063:	data_out=16'h8a00;
17'h5064:	data_out=16'h8a00;
17'h5065:	data_out=16'ha00;
17'h5066:	data_out=16'h9f6;
17'h5067:	data_out=16'h8985;
17'h5068:	data_out=16'h9ff;
17'h5069:	data_out=16'h8a00;
17'h506a:	data_out=16'ha00;
17'h506b:	data_out=16'ha00;
17'h506c:	data_out=16'h510;
17'h506d:	data_out=16'h8a00;
17'h506e:	data_out=16'ha00;
17'h506f:	data_out=16'ha00;
17'h5070:	data_out=16'ha00;
17'h5071:	data_out=16'he9;
17'h5072:	data_out=16'ha00;
17'h5073:	data_out=16'ha00;
17'h5074:	data_out=16'ha00;
17'h5075:	data_out=16'h9f8;
17'h5076:	data_out=16'h8a00;
17'h5077:	data_out=16'h8857;
17'h5078:	data_out=16'h9f6;
17'h5079:	data_out=16'h8a00;
17'h507a:	data_out=16'h89ff;
17'h507b:	data_out=16'h9ff;
17'h507c:	data_out=16'h87fc;
17'h507d:	data_out=16'h9e8;
17'h507e:	data_out=16'h89ff;
17'h507f:	data_out=16'h9ca;
17'h5080:	data_out=16'h9e2;
17'h5081:	data_out=16'h9fc;
17'h5082:	data_out=16'h89a3;
17'h5083:	data_out=16'h89d1;
17'h5084:	data_out=16'h9fe;
17'h5085:	data_out=16'h9fc;
17'h5086:	data_out=16'h8a00;
17'h5087:	data_out=16'ha00;
17'h5088:	data_out=16'h8a00;
17'h5089:	data_out=16'h89bd;
17'h508a:	data_out=16'ha00;
17'h508b:	data_out=16'h8a00;
17'h508c:	data_out=16'h89ff;
17'h508d:	data_out=16'h822c;
17'h508e:	data_out=16'ha00;
17'h508f:	data_out=16'h88d5;
17'h5090:	data_out=16'h89fd;
17'h5091:	data_out=16'ha00;
17'h5092:	data_out=16'h89fd;
17'h5093:	data_out=16'h6a9;
17'h5094:	data_out=16'h89f9;
17'h5095:	data_out=16'ha00;
17'h5096:	data_out=16'ha00;
17'h5097:	data_out=16'h89fa;
17'h5098:	data_out=16'h9fa;
17'h5099:	data_out=16'h917;
17'h509a:	data_out=16'h9f6;
17'h509b:	data_out=16'h8a00;
17'h509c:	data_out=16'h107;
17'h509d:	data_out=16'h5ae;
17'h509e:	data_out=16'h88ed;
17'h509f:	data_out=16'h23b;
17'h50a0:	data_out=16'h8448;
17'h50a1:	data_out=16'ha00;
17'h50a2:	data_out=16'h89ff;
17'h50a3:	data_out=16'ha00;
17'h50a4:	data_out=16'ha00;
17'h50a5:	data_out=16'h8086;
17'h50a6:	data_out=16'h89e8;
17'h50a7:	data_out=16'h896b;
17'h50a8:	data_out=16'h9ff;
17'h50a9:	data_out=16'h89e9;
17'h50aa:	data_out=16'h892b;
17'h50ab:	data_out=16'h8a00;
17'h50ac:	data_out=16'ha00;
17'h50ad:	data_out=16'h89f7;
17'h50ae:	data_out=16'h89fe;
17'h50af:	data_out=16'h8912;
17'h50b0:	data_out=16'h9fe;
17'h50b1:	data_out=16'ha00;
17'h50b2:	data_out=16'h9f1;
17'h50b3:	data_out=16'h89fe;
17'h50b4:	data_out=16'h84cb;
17'h50b5:	data_out=16'h920;
17'h50b6:	data_out=16'h89ff;
17'h50b7:	data_out=16'h89d7;
17'h50b8:	data_out=16'h8a00;
17'h50b9:	data_out=16'h89fd;
17'h50ba:	data_out=16'h8775;
17'h50bb:	data_out=16'h9ec;
17'h50bc:	data_out=16'h8a00;
17'h50bd:	data_out=16'h9f1;
17'h50be:	data_out=16'h9ff;
17'h50bf:	data_out=16'h9fb;
17'h50c0:	data_out=16'h9ff;
17'h50c1:	data_out=16'h8a00;
17'h50c2:	data_out=16'h8a00;
17'h50c3:	data_out=16'ha00;
17'h50c4:	data_out=16'h9f8;
17'h50c5:	data_out=16'ha00;
17'h50c6:	data_out=16'h8a00;
17'h50c7:	data_out=16'h89ee;
17'h50c8:	data_out=16'h89ec;
17'h50c9:	data_out=16'h3e2;
17'h50ca:	data_out=16'h87e6;
17'h50cb:	data_out=16'h8a00;
17'h50cc:	data_out=16'hf6;
17'h50cd:	data_out=16'h89ff;
17'h50ce:	data_out=16'h8a00;
17'h50cf:	data_out=16'h9c6;
17'h50d0:	data_out=16'h81a9;
17'h50d1:	data_out=16'h9ed;
17'h50d2:	data_out=16'h9fe;
17'h50d3:	data_out=16'h8a00;
17'h50d4:	data_out=16'h89ae;
17'h50d5:	data_out=16'h87c8;
17'h50d6:	data_out=16'h933;
17'h50d7:	data_out=16'ha00;
17'h50d8:	data_out=16'h89f8;
17'h50d9:	data_out=16'ha00;
17'h50da:	data_out=16'h8a00;
17'h50db:	data_out=16'h9ed;
17'h50dc:	data_out=16'h89d7;
17'h50dd:	data_out=16'h9f0;
17'h50de:	data_out=16'h8811;
17'h50df:	data_out=16'h8162;
17'h50e0:	data_out=16'h89ec;
17'h50e1:	data_out=16'h9f8;
17'h50e2:	data_out=16'h89fd;
17'h50e3:	data_out=16'h8a00;
17'h50e4:	data_out=16'h89ff;
17'h50e5:	data_out=16'ha00;
17'h50e6:	data_out=16'h210;
17'h50e7:	data_out=16'h89bb;
17'h50e8:	data_out=16'ha00;
17'h50e9:	data_out=16'h8a00;
17'h50ea:	data_out=16'ha00;
17'h50eb:	data_out=16'ha00;
17'h50ec:	data_out=16'ha00;
17'h50ed:	data_out=16'h8a00;
17'h50ee:	data_out=16'ha00;
17'h50ef:	data_out=16'h9f7;
17'h50f0:	data_out=16'ha00;
17'h50f1:	data_out=16'h912;
17'h50f2:	data_out=16'ha00;
17'h50f3:	data_out=16'ha00;
17'h50f4:	data_out=16'h9fe;
17'h50f5:	data_out=16'h9e8;
17'h50f6:	data_out=16'h89ff;
17'h50f7:	data_out=16'h89dd;
17'h50f8:	data_out=16'h9e3;
17'h50f9:	data_out=16'h8a00;
17'h50fa:	data_out=16'h89fd;
17'h50fb:	data_out=16'h9ff;
17'h50fc:	data_out=16'h9fb;
17'h50fd:	data_out=16'h802b;
17'h50fe:	data_out=16'h8a00;
17'h50ff:	data_out=16'h9ec;
17'h5100:	data_out=16'h9f7;
17'h5101:	data_out=16'h8020;
17'h5102:	data_out=16'h1c1;
17'h5103:	data_out=16'h89f4;
17'h5104:	data_out=16'ha00;
17'h5105:	data_out=16'h9ee;
17'h5106:	data_out=16'h82eb;
17'h5107:	data_out=16'ha00;
17'h5108:	data_out=16'h8a00;
17'h5109:	data_out=16'h89fa;
17'h510a:	data_out=16'ha00;
17'h510b:	data_out=16'h8a00;
17'h510c:	data_out=16'h413;
17'h510d:	data_out=16'h9f0;
17'h510e:	data_out=16'ha00;
17'h510f:	data_out=16'h9fa;
17'h5110:	data_out=16'h8a00;
17'h5111:	data_out=16'h9f8;
17'h5112:	data_out=16'h8902;
17'h5113:	data_out=16'h45f;
17'h5114:	data_out=16'h89ff;
17'h5115:	data_out=16'ha00;
17'h5116:	data_out=16'ha00;
17'h5117:	data_out=16'h8a00;
17'h5118:	data_out=16'ha00;
17'h5119:	data_out=16'h89f2;
17'h511a:	data_out=16'h9ee;
17'h511b:	data_out=16'h8a00;
17'h511c:	data_out=16'h2c3;
17'h511d:	data_out=16'h820e;
17'h511e:	data_out=16'h888a;
17'h511f:	data_out=16'h44e;
17'h5120:	data_out=16'h87ce;
17'h5121:	data_out=16'ha00;
17'h5122:	data_out=16'h8a00;
17'h5123:	data_out=16'ha00;
17'h5124:	data_out=16'ha00;
17'h5125:	data_out=16'h81b6;
17'h5126:	data_out=16'h8945;
17'h5127:	data_out=16'h89d5;
17'h5128:	data_out=16'ha00;
17'h5129:	data_out=16'h89f5;
17'h512a:	data_out=16'h9e7;
17'h512b:	data_out=16'h8a00;
17'h512c:	data_out=16'ha00;
17'h512d:	data_out=16'h89fe;
17'h512e:	data_out=16'h89ff;
17'h512f:	data_out=16'h89d0;
17'h5130:	data_out=16'h9bd;
17'h5131:	data_out=16'ha00;
17'h5132:	data_out=16'h9e4;
17'h5133:	data_out=16'h8a00;
17'h5134:	data_out=16'h85e1;
17'h5135:	data_out=16'h42f;
17'h5136:	data_out=16'h89f3;
17'h5137:	data_out=16'h8848;
17'h5138:	data_out=16'h8a00;
17'h5139:	data_out=16'h8a00;
17'h513a:	data_out=16'h6be;
17'h513b:	data_out=16'h6d6;
17'h513c:	data_out=16'h8a00;
17'h513d:	data_out=16'h9fe;
17'h513e:	data_out=16'ha00;
17'h513f:	data_out=16'h9ed;
17'h5140:	data_out=16'h9fa;
17'h5141:	data_out=16'h8a00;
17'h5142:	data_out=16'h89fc;
17'h5143:	data_out=16'h9ff;
17'h5144:	data_out=16'h9f9;
17'h5145:	data_out=16'ha00;
17'h5146:	data_out=16'h8a00;
17'h5147:	data_out=16'h6f5;
17'h5148:	data_out=16'h89ff;
17'h5149:	data_out=16'h21e;
17'h514a:	data_out=16'h16;
17'h514b:	data_out=16'h8a00;
17'h514c:	data_out=16'h9ff;
17'h514d:	data_out=16'h8a00;
17'h514e:	data_out=16'h811b;
17'h514f:	data_out=16'h9fa;
17'h5150:	data_out=16'h5d5;
17'h5151:	data_out=16'ha00;
17'h5152:	data_out=16'h9fe;
17'h5153:	data_out=16'h8a00;
17'h5154:	data_out=16'h89ec;
17'h5155:	data_out=16'h86b4;
17'h5156:	data_out=16'h9ea;
17'h5157:	data_out=16'ha00;
17'h5158:	data_out=16'h8844;
17'h5159:	data_out=16'ha00;
17'h515a:	data_out=16'h8a00;
17'h515b:	data_out=16'h9f4;
17'h515c:	data_out=16'h8a00;
17'h515d:	data_out=16'h9ec;
17'h515e:	data_out=16'h892e;
17'h515f:	data_out=16'h9fc;
17'h5160:	data_out=16'h880b;
17'h5161:	data_out=16'h9f4;
17'h5162:	data_out=16'h8a00;
17'h5163:	data_out=16'h8a00;
17'h5164:	data_out=16'h8a00;
17'h5165:	data_out=16'h298;
17'h5166:	data_out=16'h88be;
17'h5167:	data_out=16'h89f0;
17'h5168:	data_out=16'ha00;
17'h5169:	data_out=16'h89f8;
17'h516a:	data_out=16'ha00;
17'h516b:	data_out=16'ha00;
17'h516c:	data_out=16'ha00;
17'h516d:	data_out=16'h8a00;
17'h516e:	data_out=16'ha00;
17'h516f:	data_out=16'h9e5;
17'h5170:	data_out=16'ha00;
17'h5171:	data_out=16'ha00;
17'h5172:	data_out=16'ha00;
17'h5173:	data_out=16'h9ee;
17'h5174:	data_out=16'h9ec;
17'h5175:	data_out=16'h9db;
17'h5176:	data_out=16'h89ff;
17'h5177:	data_out=16'h8407;
17'h5178:	data_out=16'h84c;
17'h5179:	data_out=16'h89e9;
17'h517a:	data_out=16'h8a00;
17'h517b:	data_out=16'ha00;
17'h517c:	data_out=16'ha00;
17'h517d:	data_out=16'h80df;
17'h517e:	data_out=16'h8982;
17'h517f:	data_out=16'h9eb;
17'h5180:	data_out=16'h8a2;
17'h5181:	data_out=16'h89f4;
17'h5182:	data_out=16'h9fc;
17'h5183:	data_out=16'h85a9;
17'h5184:	data_out=16'ha00;
17'h5185:	data_out=16'h9f5;
17'h5186:	data_out=16'h9b2;
17'h5187:	data_out=16'ha00;
17'h5188:	data_out=16'h3cf;
17'h5189:	data_out=16'h924;
17'h518a:	data_out=16'ha00;
17'h518b:	data_out=16'h8a00;
17'h518c:	data_out=16'h9e3;
17'h518d:	data_out=16'ha00;
17'h518e:	data_out=16'ha00;
17'h518f:	data_out=16'h9fe;
17'h5190:	data_out=16'h89ff;
17'h5191:	data_out=16'h209;
17'h5192:	data_out=16'h1c0;
17'h5193:	data_out=16'ha00;
17'h5194:	data_out=16'h8a00;
17'h5195:	data_out=16'ha00;
17'h5196:	data_out=16'ha00;
17'h5197:	data_out=16'h8a00;
17'h5198:	data_out=16'ha00;
17'h5199:	data_out=16'h89fd;
17'h519a:	data_out=16'h9f4;
17'h519b:	data_out=16'h8a00;
17'h519c:	data_out=16'h89ff;
17'h519d:	data_out=16'h8a00;
17'h519e:	data_out=16'h87a8;
17'h519f:	data_out=16'h9d4;
17'h51a0:	data_out=16'h89ed;
17'h51a1:	data_out=16'ha00;
17'h51a2:	data_out=16'h87e9;
17'h51a3:	data_out=16'ha00;
17'h51a4:	data_out=16'ha00;
17'h51a5:	data_out=16'ha00;
17'h51a6:	data_out=16'h9fc;
17'h51a7:	data_out=16'h89f3;
17'h51a8:	data_out=16'ha00;
17'h51a9:	data_out=16'h88d3;
17'h51aa:	data_out=16'h9fc;
17'h51ab:	data_out=16'h8a00;
17'h51ac:	data_out=16'ha00;
17'h51ad:	data_out=16'h8a00;
17'h51ae:	data_out=16'h659;
17'h51af:	data_out=16'h89ff;
17'h51b0:	data_out=16'h9ff;
17'h51b1:	data_out=16'h8568;
17'h51b2:	data_out=16'h9f2;
17'h51b3:	data_out=16'h8a00;
17'h51b4:	data_out=16'h89f0;
17'h51b5:	data_out=16'h57b;
17'h51b6:	data_out=16'h5e0;
17'h51b7:	data_out=16'h9fa;
17'h51b8:	data_out=16'h8a00;
17'h51b9:	data_out=16'h8a00;
17'h51ba:	data_out=16'h9f9;
17'h51bb:	data_out=16'h546;
17'h51bc:	data_out=16'h8a00;
17'h51bd:	data_out=16'ha00;
17'h51be:	data_out=16'ha00;
17'h51bf:	data_out=16'h9f5;
17'h51c0:	data_out=16'h9ff;
17'h51c1:	data_out=16'h89ef;
17'h51c2:	data_out=16'h9f5;
17'h51c3:	data_out=16'h9f2;
17'h51c4:	data_out=16'h414;
17'h51c5:	data_out=16'ha00;
17'h51c6:	data_out=16'h8a00;
17'h51c7:	data_out=16'h9fd;
17'h51c8:	data_out=16'h329;
17'h51c9:	data_out=16'ha00;
17'h51ca:	data_out=16'h45a;
17'h51cb:	data_out=16'h3d3;
17'h51cc:	data_out=16'ha00;
17'h51cd:	data_out=16'h8a00;
17'h51ce:	data_out=16'h7ab;
17'h51cf:	data_out=16'ha00;
17'h51d0:	data_out=16'h656;
17'h51d1:	data_out=16'ha00;
17'h51d2:	data_out=16'ha00;
17'h51d3:	data_out=16'h8a00;
17'h51d4:	data_out=16'h89fb;
17'h51d5:	data_out=16'h97c;
17'h51d6:	data_out=16'h9fb;
17'h51d7:	data_out=16'h9ff;
17'h51d8:	data_out=16'h81a;
17'h51d9:	data_out=16'ha00;
17'h51da:	data_out=16'h8a00;
17'h51db:	data_out=16'h73e;
17'h51dc:	data_out=16'h8a00;
17'h51dd:	data_out=16'h9f4;
17'h51de:	data_out=16'h89f1;
17'h51df:	data_out=16'h9ff;
17'h51e0:	data_out=16'h9ec;
17'h51e1:	data_out=16'h9fc;
17'h51e2:	data_out=16'h8a00;
17'h51e3:	data_out=16'h8a00;
17'h51e4:	data_out=16'h8a00;
17'h51e5:	data_out=16'h251;
17'h51e6:	data_out=16'h89d8;
17'h51e7:	data_out=16'h8a00;
17'h51e8:	data_out=16'ha00;
17'h51e9:	data_out=16'h3f8;
17'h51ea:	data_out=16'ha00;
17'h51eb:	data_out=16'h9f8;
17'h51ec:	data_out=16'ha00;
17'h51ed:	data_out=16'h8a00;
17'h51ee:	data_out=16'ha00;
17'h51ef:	data_out=16'h9ed;
17'h51f0:	data_out=16'ha00;
17'h51f1:	data_out=16'ha00;
17'h51f2:	data_out=16'h9fc;
17'h51f3:	data_out=16'h9f3;
17'h51f4:	data_out=16'ha00;
17'h51f5:	data_out=16'h11e;
17'h51f6:	data_out=16'h8a00;
17'h51f7:	data_out=16'h9f7;
17'h51f8:	data_out=16'h5e2;
17'h51f9:	data_out=16'h532;
17'h51fa:	data_out=16'h8a00;
17'h51fb:	data_out=16'ha00;
17'h51fc:	data_out=16'ha00;
17'h51fd:	data_out=16'h763;
17'h51fe:	data_out=16'h8716;
17'h51ff:	data_out=16'h9ef;
17'h5200:	data_out=16'h83e8;
17'h5201:	data_out=16'h89f8;
17'h5202:	data_out=16'h9fa;
17'h5203:	data_out=16'h813;
17'h5204:	data_out=16'h952;
17'h5205:	data_out=16'h9ff;
17'h5206:	data_out=16'h9f6;
17'h5207:	data_out=16'ha00;
17'h5208:	data_out=16'h684;
17'h5209:	data_out=16'h9ee;
17'h520a:	data_out=16'h83c4;
17'h520b:	data_out=16'h8a00;
17'h520c:	data_out=16'ha00;
17'h520d:	data_out=16'ha00;
17'h520e:	data_out=16'ha00;
17'h520f:	data_out=16'h9fd;
17'h5210:	data_out=16'h83cf;
17'h5211:	data_out=16'h23a;
17'h5212:	data_out=16'h850;
17'h5213:	data_out=16'ha00;
17'h5214:	data_out=16'h89ff;
17'h5215:	data_out=16'ha00;
17'h5216:	data_out=16'ha00;
17'h5217:	data_out=16'h89fa;
17'h5218:	data_out=16'h9ff;
17'h5219:	data_out=16'h89f6;
17'h521a:	data_out=16'h9fe;
17'h521b:	data_out=16'h89fe;
17'h521c:	data_out=16'h2df;
17'h521d:	data_out=16'h8a00;
17'h521e:	data_out=16'h823e;
17'h521f:	data_out=16'h9f1;
17'h5220:	data_out=16'h89fc;
17'h5221:	data_out=16'ha00;
17'h5222:	data_out=16'h830f;
17'h5223:	data_out=16'ha00;
17'h5224:	data_out=16'ha00;
17'h5225:	data_out=16'ha00;
17'h5226:	data_out=16'h257;
17'h5227:	data_out=16'h89ff;
17'h5228:	data_out=16'ha00;
17'h5229:	data_out=16'h86c2;
17'h522a:	data_out=16'h9f8;
17'h522b:	data_out=16'h8a00;
17'h522c:	data_out=16'ha00;
17'h522d:	data_out=16'h8a00;
17'h522e:	data_out=16'h9f1;
17'h522f:	data_out=16'h89fc;
17'h5230:	data_out=16'h9fd;
17'h5231:	data_out=16'h89f3;
17'h5232:	data_out=16'h9f5;
17'h5233:	data_out=16'h8a00;
17'h5234:	data_out=16'h89fe;
17'h5235:	data_out=16'h517;
17'h5236:	data_out=16'h817;
17'h5237:	data_out=16'h9f9;
17'h5238:	data_out=16'h8a00;
17'h5239:	data_out=16'h8a00;
17'h523a:	data_out=16'h9f4;
17'h523b:	data_out=16'h67c;
17'h523c:	data_out=16'h8752;
17'h523d:	data_out=16'h9c3;
17'h523e:	data_out=16'ha00;
17'h523f:	data_out=16'h9ff;
17'h5240:	data_out=16'h9f8;
17'h5241:	data_out=16'h85;
17'h5242:	data_out=16'ha00;
17'h5243:	data_out=16'h9fd;
17'h5244:	data_out=16'h4;
17'h5245:	data_out=16'ha00;
17'h5246:	data_out=16'h8a00;
17'h5247:	data_out=16'h9d9;
17'h5248:	data_out=16'h9fd;
17'h5249:	data_out=16'ha00;
17'h524a:	data_out=16'h6a0;
17'h524b:	data_out=16'h9fe;
17'h524c:	data_out=16'ha00;
17'h524d:	data_out=16'h8503;
17'h524e:	data_out=16'h904;
17'h524f:	data_out=16'ha00;
17'h5250:	data_out=16'h9f5;
17'h5251:	data_out=16'h9fc;
17'h5252:	data_out=16'ha00;
17'h5253:	data_out=16'h8a00;
17'h5254:	data_out=16'h8a00;
17'h5255:	data_out=16'h9fd;
17'h5256:	data_out=16'h9b3;
17'h5257:	data_out=16'h9f8;
17'h5258:	data_out=16'h9eb;
17'h5259:	data_out=16'h9ff;
17'h525a:	data_out=16'h8a00;
17'h525b:	data_out=16'h711;
17'h525c:	data_out=16'h8a00;
17'h525d:	data_out=16'h9fa;
17'h525e:	data_out=16'h89f3;
17'h525f:	data_out=16'h9f8;
17'h5260:	data_out=16'h124;
17'h5261:	data_out=16'h9fd;
17'h5262:	data_out=16'h89fc;
17'h5263:	data_out=16'h8a00;
17'h5264:	data_out=16'h8a00;
17'h5265:	data_out=16'h191;
17'h5266:	data_out=16'h89f0;
17'h5267:	data_out=16'h8a00;
17'h5268:	data_out=16'ha00;
17'h5269:	data_out=16'h628;
17'h526a:	data_out=16'ha00;
17'h526b:	data_out=16'h9fd;
17'h526c:	data_out=16'h9fd;
17'h526d:	data_out=16'h8a00;
17'h526e:	data_out=16'ha00;
17'h526f:	data_out=16'ha00;
17'h5270:	data_out=16'ha00;
17'h5271:	data_out=16'ha00;
17'h5272:	data_out=16'h9fe;
17'h5273:	data_out=16'h9fd;
17'h5274:	data_out=16'ha00;
17'h5275:	data_out=16'h4d2;
17'h5276:	data_out=16'h8a00;
17'h5277:	data_out=16'h9fe;
17'h5278:	data_out=16'h9ea;
17'h5279:	data_out=16'h8e4;
17'h527a:	data_out=16'h8a00;
17'h527b:	data_out=16'ha00;
17'h527c:	data_out=16'h9ff;
17'h527d:	data_out=16'h9f5;
17'h527e:	data_out=16'h84bb;
17'h527f:	data_out=16'h9fb;
17'h5280:	data_out=16'h89ce;
17'h5281:	data_out=16'h801d;
17'h5282:	data_out=16'ha00;
17'h5283:	data_out=16'h83ea;
17'h5284:	data_out=16'h9c9;
17'h5285:	data_out=16'ha00;
17'h5286:	data_out=16'h293;
17'h5287:	data_out=16'ha00;
17'h5288:	data_out=16'h990;
17'h5289:	data_out=16'h4e;
17'h528a:	data_out=16'h8012;
17'h528b:	data_out=16'h8a00;
17'h528c:	data_out=16'h9f3;
17'h528d:	data_out=16'h81c4;
17'h528e:	data_out=16'h87a;
17'h528f:	data_out=16'ha00;
17'h5290:	data_out=16'h81e1;
17'h5291:	data_out=16'h91c;
17'h5292:	data_out=16'h13c;
17'h5293:	data_out=16'h822c;
17'h5294:	data_out=16'h85a8;
17'h5295:	data_out=16'h87d;
17'h5296:	data_out=16'h682;
17'h5297:	data_out=16'h89fd;
17'h5298:	data_out=16'h9fc;
17'h5299:	data_out=16'h332;
17'h529a:	data_out=16'ha00;
17'h529b:	data_out=16'h89f6;
17'h529c:	data_out=16'h944;
17'h529d:	data_out=16'h837f;
17'h529e:	data_out=16'h81f1;
17'h529f:	data_out=16'h936;
17'h52a0:	data_out=16'h88dd;
17'h52a1:	data_out=16'h85c;
17'h52a2:	data_out=16'h813e;
17'h52a3:	data_out=16'h9c9;
17'h52a4:	data_out=16'h9cb;
17'h52a5:	data_out=16'h678;
17'h52a6:	data_out=16'h815c;
17'h52a7:	data_out=16'h8671;
17'h52a8:	data_out=16'h835;
17'h52a9:	data_out=16'h85ee;
17'h52aa:	data_out=16'h9ff;
17'h52ab:	data_out=16'h8a00;
17'h52ac:	data_out=16'h5a3;
17'h52ad:	data_out=16'h89f3;
17'h52ae:	data_out=16'ha00;
17'h52af:	data_out=16'h8753;
17'h52b0:	data_out=16'ha00;
17'h52b1:	data_out=16'h89fd;
17'h52b2:	data_out=16'ha00;
17'h52b3:	data_out=16'h851f;
17'h52b4:	data_out=16'h82ee;
17'h52b5:	data_out=16'h84a;
17'h52b6:	data_out=16'h830;
17'h52b7:	data_out=16'ha00;
17'h52b8:	data_out=16'h998;
17'h52b9:	data_out=16'h840e;
17'h52ba:	data_out=16'h1af;
17'h52bb:	data_out=16'h2c;
17'h52bc:	data_out=16'h7c6;
17'h52bd:	data_out=16'h748;
17'h52be:	data_out=16'h834;
17'h52bf:	data_out=16'ha00;
17'h52c0:	data_out=16'ha00;
17'h52c1:	data_out=16'h881;
17'h52c2:	data_out=16'h8d1;
17'h52c3:	data_out=16'h257;
17'h52c4:	data_out=16'h853c;
17'h52c5:	data_out=16'h88e;
17'h52c6:	data_out=16'h803d;
17'h52c7:	data_out=16'h4c8;
17'h52c8:	data_out=16'h3df;
17'h52c9:	data_out=16'h659;
17'h52ca:	data_out=16'h8dc;
17'h52cb:	data_out=16'h4ba;
17'h52cc:	data_out=16'ha00;
17'h52cd:	data_out=16'h81a4;
17'h52ce:	data_out=16'h9ff;
17'h52cf:	data_out=16'ha00;
17'h52d0:	data_out=16'h842;
17'h52d1:	data_out=16'h9e7;
17'h52d2:	data_out=16'ha00;
17'h52d3:	data_out=16'h89f3;
17'h52d4:	data_out=16'hf7;
17'h52d5:	data_out=16'h9bc;
17'h52d6:	data_out=16'h9fd;
17'h52d7:	data_out=16'h9ff;
17'h52d8:	data_out=16'h9e4;
17'h52d9:	data_out=16'ha00;
17'h52da:	data_out=16'h89fe;
17'h52db:	data_out=16'h973;
17'h52dc:	data_out=16'h8875;
17'h52dd:	data_out=16'h9d7;
17'h52de:	data_out=16'h86b3;
17'h52df:	data_out=16'h6dd;
17'h52e0:	data_out=16'h302;
17'h52e1:	data_out=16'ha00;
17'h52e2:	data_out=16'h89f8;
17'h52e3:	data_out=16'h8549;
17'h52e4:	data_out=16'h8a00;
17'h52e5:	data_out=16'h83f2;
17'h52e6:	data_out=16'h8899;
17'h52e7:	data_out=16'h844b;
17'h52e8:	data_out=16'h846;
17'h52e9:	data_out=16'h950;
17'h52ea:	data_out=16'h895;
17'h52eb:	data_out=16'h9b4;
17'h52ec:	data_out=16'h80;
17'h52ed:	data_out=16'h851f;
17'h52ee:	data_out=16'h895;
17'h52ef:	data_out=16'h826;
17'h52f0:	data_out=16'h887;
17'h52f1:	data_out=16'ha00;
17'h52f2:	data_out=16'ha00;
17'h52f3:	data_out=16'ha00;
17'h52f4:	data_out=16'ha00;
17'h52f5:	data_out=16'h274;
17'h52f6:	data_out=16'h8a00;
17'h52f7:	data_out=16'ha00;
17'h52f8:	data_out=16'h580;
17'h52f9:	data_out=16'h9ff;
17'h52fa:	data_out=16'h850c;
17'h52fb:	data_out=16'h835;
17'h52fc:	data_out=16'h937;
17'h52fd:	data_out=16'h1c7;
17'h52fe:	data_out=16'h8322;
17'h52ff:	data_out=16'h9f8;
17'h5300:	data_out=16'h8121;
17'h5301:	data_out=16'h1ef;
17'h5302:	data_out=16'h422;
17'h5303:	data_out=16'h19b;
17'h5304:	data_out=16'h736;
17'h5305:	data_out=16'h675;
17'h5306:	data_out=16'h20d;
17'h5307:	data_out=16'h472;
17'h5308:	data_out=16'h160;
17'h5309:	data_out=16'h80b7;
17'h530a:	data_out=16'h24d;
17'h530b:	data_out=16'h85ba;
17'h530c:	data_out=16'h78c;
17'h530d:	data_out=16'h1e9;
17'h530e:	data_out=16'h22b;
17'h530f:	data_out=16'h405;
17'h5310:	data_out=16'h196;
17'h5311:	data_out=16'h51d;
17'h5312:	data_out=16'h812f;
17'h5313:	data_out=16'h1a6;
17'h5314:	data_out=16'h81d7;
17'h5315:	data_out=16'h30f;
17'h5316:	data_out=16'h35f;
17'h5317:	data_out=16'h82cc;
17'h5318:	data_out=16'h281;
17'h5319:	data_out=16'h200;
17'h531a:	data_out=16'h649;
17'h531b:	data_out=16'h8257;
17'h531c:	data_out=16'h477;
17'h531d:	data_out=16'h8021;
17'h531e:	data_out=16'h8106;
17'h531f:	data_out=16'h48d;
17'h5320:	data_out=16'h8002;
17'h5321:	data_out=16'h22b;
17'h5322:	data_out=16'h8001;
17'h5323:	data_out=16'h311;
17'h5324:	data_out=16'h312;
17'h5325:	data_out=16'h36f;
17'h5326:	data_out=16'h8256;
17'h5327:	data_out=16'h8085;
17'h5328:	data_out=16'h22b;
17'h5329:	data_out=16'h819f;
17'h532a:	data_out=16'h802b;
17'h532b:	data_out=16'h8910;
17'h532c:	data_out=16'h2db;
17'h532d:	data_out=16'h8197;
17'h532e:	data_out=16'h1e8;
17'h532f:	data_out=16'h1e4;
17'h5330:	data_out=16'h5d8;
17'h5331:	data_out=16'h8127;
17'h5332:	data_out=16'h5d5;
17'h5333:	data_out=16'h8204;
17'h5334:	data_out=16'h92;
17'h5335:	data_out=16'h830;
17'h5336:	data_out=16'h26b;
17'h5337:	data_out=16'h45d;
17'h5338:	data_out=16'h450;
17'h5339:	data_out=16'h81a3;
17'h533a:	data_out=16'h800f;
17'h533b:	data_out=16'hf6;
17'h533c:	data_out=16'hb9;
17'h533d:	data_out=16'h254;
17'h533e:	data_out=16'h22b;
17'h533f:	data_out=16'h67a;
17'h5340:	data_out=16'h774;
17'h5341:	data_out=16'h33e;
17'h5342:	data_out=16'h524;
17'h5343:	data_out=16'h202;
17'h5344:	data_out=16'h177;
17'h5345:	data_out=16'h31b;
17'h5346:	data_out=16'h8261;
17'h5347:	data_out=16'h155;
17'h5348:	data_out=16'h806e;
17'h5349:	data_out=16'h3ad;
17'h534a:	data_out=16'h6b2;
17'h534b:	data_out=16'h480;
17'h534c:	data_out=16'h52d;
17'h534d:	data_out=16'h8004;
17'h534e:	data_out=16'h20f;
17'h534f:	data_out=16'h473;
17'h5350:	data_out=16'h762;
17'h5351:	data_out=16'h49a;
17'h5352:	data_out=16'h372;
17'h5353:	data_out=16'h81ef;
17'h5354:	data_out=16'h299;
17'h5355:	data_out=16'h25b;
17'h5356:	data_out=16'h2b6;
17'h5357:	data_out=16'h37a;
17'h5358:	data_out=16'h36a;
17'h5359:	data_out=16'h797;
17'h535a:	data_out=16'h82c6;
17'h535b:	data_out=16'h942;
17'h535c:	data_out=16'h16a;
17'h535d:	data_out=16'h3a5;
17'h535e:	data_out=16'h1b5;
17'h535f:	data_out=16'h1e1;
17'h5360:	data_out=16'h811a;
17'h5361:	data_out=16'h5bc;
17'h5362:	data_out=16'h822d;
17'h5363:	data_out=16'h818a;
17'h5364:	data_out=16'h811c;
17'h5365:	data_out=16'h2a4;
17'h5366:	data_out=16'h1bf;
17'h5367:	data_out=16'h8231;
17'h5368:	data_out=16'h229;
17'h5369:	data_out=16'h256;
17'h536a:	data_out=16'h22d;
17'h536b:	data_out=16'h543;
17'h536c:	data_out=16'h1a0;
17'h536d:	data_out=16'h81e4;
17'h536e:	data_out=16'h22d;
17'h536f:	data_out=16'h324;
17'h5370:	data_out=16'h22c;
17'h5371:	data_out=16'h1cb;
17'h5372:	data_out=16'h568;
17'h5373:	data_out=16'h66e;
17'h5374:	data_out=16'h5e4;
17'h5375:	data_out=16'h21d;
17'h5376:	data_out=16'h8776;
17'h5377:	data_out=16'h6c0;
17'h5378:	data_out=16'h21d;
17'h5379:	data_out=16'h2e8;
17'h537a:	data_out=16'h81b0;
17'h537b:	data_out=16'h22b;
17'h537c:	data_out=16'h22b;
17'h537d:	data_out=16'h1f5;
17'h537e:	data_out=16'h811a;
17'h537f:	data_out=16'h873;
17'h5380:	data_out=16'h81c3;
17'h5381:	data_out=16'h815d;
17'h5382:	data_out=16'h812d;
17'h5383:	data_out=16'h8057;
17'h5384:	data_out=16'hf0;
17'h5385:	data_out=16'h75;
17'h5386:	data_out=16'h60;
17'h5387:	data_out=16'hdc;
17'h5388:	data_out=16'h821e;
17'h5389:	data_out=16'h8023;
17'h538a:	data_out=16'h8108;
17'h538b:	data_out=16'h80f9;
17'h538c:	data_out=16'h287;
17'h538d:	data_out=16'h800d;
17'h538e:	data_out=16'h8029;
17'h538f:	data_out=16'h80fd;
17'h5390:	data_out=16'h8034;
17'h5391:	data_out=16'h37;
17'h5392:	data_out=16'h80cd;
17'h5393:	data_out=16'h2a;
17'h5394:	data_out=16'h815b;
17'h5395:	data_out=16'h8044;
17'h5396:	data_out=16'h808c;
17'h5397:	data_out=16'h8144;
17'h5398:	data_out=16'h8035;
17'h5399:	data_out=16'h1dc;
17'h539a:	data_out=16'h167;
17'h539b:	data_out=16'h80e2;
17'h539c:	data_out=16'h80bf;
17'h539d:	data_out=16'h81ab;
17'h539e:	data_out=16'h816d;
17'h539f:	data_out=16'h8037;
17'h53a0:	data_out=16'h815d;
17'h53a1:	data_out=16'h8023;
17'h53a2:	data_out=16'h96;
17'h53a3:	data_out=16'h8042;
17'h53a4:	data_out=16'h803f;
17'h53a5:	data_out=16'h173;
17'h53a6:	data_out=16'h8225;
17'h53a7:	data_out=16'h8212;
17'h53a8:	data_out=16'h801d;
17'h53a9:	data_out=16'h807f;
17'h53aa:	data_out=16'h8170;
17'h53ab:	data_out=16'h8217;
17'h53ac:	data_out=16'h807c;
17'h53ad:	data_out=16'h5e;
17'h53ae:	data_out=16'h811a;
17'h53af:	data_out=16'h8084;
17'h53b0:	data_out=16'h112;
17'h53b1:	data_out=16'h8073;
17'h53b2:	data_out=16'h111;
17'h53b3:	data_out=16'h816e;
17'h53b4:	data_out=16'h8061;
17'h53b5:	data_out=16'h13a;
17'h53b6:	data_out=16'h81ad;
17'h53b7:	data_out=16'h811b;
17'h53b8:	data_out=16'h8039;
17'h53b9:	data_out=16'h8178;
17'h53ba:	data_out=16'h8057;
17'h53bb:	data_out=16'h807c;
17'h53bc:	data_out=16'h8199;
17'h53bd:	data_out=16'h8118;
17'h53be:	data_out=16'h8012;
17'h53bf:	data_out=16'h122;
17'h53c0:	data_out=16'h14b;
17'h53c1:	data_out=16'h8109;
17'h53c2:	data_out=16'h252;
17'h53c3:	data_out=16'hd4;
17'h53c4:	data_out=16'h8085;
17'h53c5:	data_out=16'h808d;
17'h53c6:	data_out=16'h816c;
17'h53c7:	data_out=16'h800e;
17'h53c8:	data_out=16'h8013;
17'h53c9:	data_out=16'h16a;
17'h53ca:	data_out=16'h193;
17'h53cb:	data_out=16'h2cb;
17'h53cc:	data_out=16'h224;
17'h53cd:	data_out=16'haa;
17'h53ce:	data_out=16'h8069;
17'h53cf:	data_out=16'h200;
17'h53d0:	data_out=16'hf3;
17'h53d1:	data_out=16'h811e;
17'h53d2:	data_out=16'h803a;
17'h53d3:	data_out=16'h819e;
17'h53d4:	data_out=16'h8124;
17'h53d5:	data_out=16'h8189;
17'h53d6:	data_out=16'h80cd;
17'h53d7:	data_out=16'h8091;
17'h53d8:	data_out=16'h81a9;
17'h53d9:	data_out=16'hc8;
17'h53da:	data_out=16'h8160;
17'h53db:	data_out=16'h8086;
17'h53dc:	data_out=16'h8097;
17'h53dd:	data_out=16'h8066;
17'h53de:	data_out=16'h801c;
17'h53df:	data_out=16'h803f;
17'h53e0:	data_out=16'h8151;
17'h53e1:	data_out=16'h802b;
17'h53e2:	data_out=16'h8159;
17'h53e3:	data_out=16'h815d;
17'h53e4:	data_out=16'h80c8;
17'h53e5:	data_out=16'h1b9;
17'h53e6:	data_out=16'h1df;
17'h53e7:	data_out=16'h80ad;
17'h53e8:	data_out=16'h8018;
17'h53e9:	data_out=16'h81f1;
17'h53ea:	data_out=16'h801b;
17'h53eb:	data_out=16'h9e;
17'h53ec:	data_out=16'h8154;
17'h53ed:	data_out=16'h817b;
17'h53ee:	data_out=16'h8027;
17'h53ef:	data_out=16'hb3;
17'h53f0:	data_out=16'h8020;
17'h53f1:	data_out=16'h8159;
17'h53f2:	data_out=16'h6b;
17'h53f3:	data_out=16'h60;
17'h53f4:	data_out=16'h11a;
17'h53f5:	data_out=16'h809f;
17'h53f6:	data_out=16'h81fc;
17'h53f7:	data_out=16'h1a0;
17'h53f8:	data_out=16'h140;
17'h53f9:	data_out=16'h8176;
17'h53fa:	data_out=16'h816a;
17'h53fb:	data_out=16'h8022;
17'h53fc:	data_out=16'h8099;
17'h53fd:	data_out=16'h70;
17'h53fe:	data_out=16'h8070;
17'h53ff:	data_out=16'h111;
17'h5400:	data_out=16'h8006;
17'h5401:	data_out=16'h5;
17'h5402:	data_out=16'h7;
17'h5403:	data_out=16'h9;
17'h5404:	data_out=16'h5;
17'h5405:	data_out=16'h8007;
17'h5406:	data_out=16'h4;
17'h5407:	data_out=16'h8001;
17'h5408:	data_out=16'h1;
17'h5409:	data_out=16'h4;
17'h540a:	data_out=16'h5;
17'h540b:	data_out=16'h8004;
17'h540c:	data_out=16'h6;
17'h540d:	data_out=16'h8007;
17'h540e:	data_out=16'h8;
17'h540f:	data_out=16'h8001;
17'h5410:	data_out=16'h8003;
17'h5411:	data_out=16'h8001;
17'h5412:	data_out=16'h4;
17'h5413:	data_out=16'h8008;
17'h5414:	data_out=16'h5;
17'h5415:	data_out=16'h2;
17'h5416:	data_out=16'h8008;
17'h5417:	data_out=16'h8007;
17'h5418:	data_out=16'h8006;
17'h5419:	data_out=16'h8007;
17'h541a:	data_out=16'h8007;
17'h541b:	data_out=16'h8004;
17'h541c:	data_out=16'h4;
17'h541d:	data_out=16'h4;
17'h541e:	data_out=16'h9;
17'h541f:	data_out=16'h7;
17'h5420:	data_out=16'h0;
17'h5421:	data_out=16'h7;
17'h5422:	data_out=16'h6;
17'h5423:	data_out=16'h8004;
17'h5424:	data_out=16'h8009;
17'h5425:	data_out=16'h1;
17'h5426:	data_out=16'h4;
17'h5427:	data_out=16'h1;
17'h5428:	data_out=16'h8005;
17'h5429:	data_out=16'h8000;
17'h542a:	data_out=16'h6;
17'h542b:	data_out=16'h8007;
17'h542c:	data_out=16'h1;
17'h542d:	data_out=16'h5;
17'h542e:	data_out=16'h1;
17'h542f:	data_out=16'h8;
17'h5430:	data_out=16'h8006;
17'h5431:	data_out=16'h8004;
17'h5432:	data_out=16'h9;
17'h5433:	data_out=16'h9;
17'h5434:	data_out=16'h7;
17'h5435:	data_out=16'h8008;
17'h5436:	data_out=16'h8008;
17'h5437:	data_out=16'h8008;
17'h5438:	data_out=16'h8006;
17'h5439:	data_out=16'h8006;
17'h543a:	data_out=16'h8002;
17'h543b:	data_out=16'h7;
17'h543c:	data_out=16'h8;
17'h543d:	data_out=16'h8003;
17'h543e:	data_out=16'h4;
17'h543f:	data_out=16'h8001;
17'h5440:	data_out=16'h8005;
17'h5441:	data_out=16'h2;
17'h5442:	data_out=16'h3;
17'h5443:	data_out=16'h8005;
17'h5444:	data_out=16'h8007;
17'h5445:	data_out=16'h8002;
17'h5446:	data_out=16'h5;
17'h5447:	data_out=16'h8002;
17'h5448:	data_out=16'h7;
17'h5449:	data_out=16'h2;
17'h544a:	data_out=16'h8000;
17'h544b:	data_out=16'h8001;
17'h544c:	data_out=16'h8003;
17'h544d:	data_out=16'h8008;
17'h544e:	data_out=16'h8003;
17'h544f:	data_out=16'h1;
17'h5450:	data_out=16'h8003;
17'h5451:	data_out=16'h8003;
17'h5452:	data_out=16'h0;
17'h5453:	data_out=16'h8005;
17'h5454:	data_out=16'h8002;
17'h5455:	data_out=16'h2;
17'h5456:	data_out=16'h8004;
17'h5457:	data_out=16'h1;
17'h5458:	data_out=16'h5;
17'h5459:	data_out=16'h3;
17'h545a:	data_out=16'h8001;
17'h545b:	data_out=16'h3;
17'h545c:	data_out=16'h8009;
17'h545d:	data_out=16'h8006;
17'h545e:	data_out=16'h8007;
17'h545f:	data_out=16'h8004;
17'h5460:	data_out=16'h5;
17'h5461:	data_out=16'h5;
17'h5462:	data_out=16'h0;
17'h5463:	data_out=16'h7;
17'h5464:	data_out=16'h8006;
17'h5465:	data_out=16'h8004;
17'h5466:	data_out=16'h8004;
17'h5467:	data_out=16'h8009;
17'h5468:	data_out=16'h7;
17'h5469:	data_out=16'h5;
17'h546a:	data_out=16'h8001;
17'h546b:	data_out=16'h8004;
17'h546c:	data_out=16'h5;
17'h546d:	data_out=16'h5;
17'h546e:	data_out=16'h6;
17'h546f:	data_out=16'h8007;
17'h5470:	data_out=16'h8007;
17'h5471:	data_out=16'h8003;
17'h5472:	data_out=16'h8003;
17'h5473:	data_out=16'h8000;
17'h5474:	data_out=16'h7;
17'h5475:	data_out=16'h3;
17'h5476:	data_out=16'h8009;
17'h5477:	data_out=16'h3;
17'h5478:	data_out=16'h8004;
17'h5479:	data_out=16'h8001;
17'h547a:	data_out=16'h8003;
17'h547b:	data_out=16'h8003;
17'h547c:	data_out=16'h3;
17'h547d:	data_out=16'h8001;
17'h547e:	data_out=16'h2;
17'h547f:	data_out=16'h8002;
17'h5480:	data_out=16'h8003;
17'h5481:	data_out=16'h8008;
17'h5482:	data_out=16'h8009;
17'h5483:	data_out=16'h8007;
17'h5484:	data_out=16'h8007;
17'h5485:	data_out=16'h5;
17'h5486:	data_out=16'h2;
17'h5487:	data_out=16'h8008;
17'h5488:	data_out=16'h8000;
17'h5489:	data_out=16'h8;
17'h548a:	data_out=16'h8003;
17'h548b:	data_out=16'h8003;
17'h548c:	data_out=16'h5;
17'h548d:	data_out=16'h8009;
17'h548e:	data_out=16'h8006;
17'h548f:	data_out=16'h3;
17'h5490:	data_out=16'h8004;
17'h5491:	data_out=16'h1;
17'h5492:	data_out=16'h8009;
17'h5493:	data_out=16'h8007;
17'h5494:	data_out=16'h8009;
17'h5495:	data_out=16'h8009;
17'h5496:	data_out=16'h800c;
17'h5497:	data_out=16'h8004;
17'h5498:	data_out=16'h0;
17'h5499:	data_out=16'h9;
17'h549a:	data_out=16'h2;
17'h549b:	data_out=16'h0;
17'h549c:	data_out=16'h8001;
17'h549d:	data_out=16'h8001;
17'h549e:	data_out=16'h7;
17'h549f:	data_out=16'h8004;
17'h54a0:	data_out=16'h8;
17'h54a1:	data_out=16'h8009;
17'h54a2:	data_out=16'h2;
17'h54a3:	data_out=16'h8001;
17'h54a4:	data_out=16'h8006;
17'h54a5:	data_out=16'h800a;
17'h54a6:	data_out=16'h8004;
17'h54a7:	data_out=16'hc;
17'h54a8:	data_out=16'h8008;
17'h54a9:	data_out=16'h8002;
17'h54aa:	data_out=16'h800f;
17'h54ab:	data_out=16'h10;
17'h54ac:	data_out=16'h800b;
17'h54ad:	data_out=16'h8010;
17'h54ae:	data_out=16'h8006;
17'h54af:	data_out=16'h9;
17'h54b0:	data_out=16'h1;
17'h54b1:	data_out=16'ha;
17'h54b2:	data_out=16'h8007;
17'h54b3:	data_out=16'h800a;
17'h54b4:	data_out=16'h8006;
17'h54b5:	data_out=16'h8;
17'h54b6:	data_out=16'h5;
17'h54b7:	data_out=16'h3;
17'h54b8:	data_out=16'h5;
17'h54b9:	data_out=16'h0;
17'h54ba:	data_out=16'h800e;
17'h54bb:	data_out=16'h8000;
17'h54bc:	data_out=16'h5;
17'h54bd:	data_out=16'h8007;
17'h54be:	data_out=16'h4;
17'h54bf:	data_out=16'h8000;
17'h54c0:	data_out=16'h8011;
17'h54c1:	data_out=16'h5;
17'h54c2:	data_out=16'h800a;
17'h54c3:	data_out=16'h9;
17'h54c4:	data_out=16'h1;
17'h54c5:	data_out=16'h8005;
17'h54c6:	data_out=16'h6;
17'h54c7:	data_out=16'h8003;
17'h54c8:	data_out=16'h8008;
17'h54c9:	data_out=16'h1;
17'h54ca:	data_out=16'h8004;
17'h54cb:	data_out=16'h8002;
17'h54cc:	data_out=16'h8011;
17'h54cd:	data_out=16'h8006;
17'h54ce:	data_out=16'h8007;
17'h54cf:	data_out=16'h8001;
17'h54d0:	data_out=16'h8011;
17'h54d1:	data_out=16'h7;
17'h54d2:	data_out=16'h8011;
17'h54d3:	data_out=16'h6;
17'h54d4:	data_out=16'h5;
17'h54d5:	data_out=16'h4;
17'h54d6:	data_out=16'h800d;
17'h54d7:	data_out=16'h8001;
17'h54d8:	data_out=16'h800b;
17'h54d9:	data_out=16'h8007;
17'h54da:	data_out=16'h8004;
17'h54db:	data_out=16'h2;
17'h54dc:	data_out=16'h9;
17'h54dd:	data_out=16'h800d;
17'h54de:	data_out=16'h2;
17'h54df:	data_out=16'h800d;
17'h54e0:	data_out=16'h8004;
17'h54e1:	data_out=16'h6;
17'h54e2:	data_out=16'hc;
17'h54e3:	data_out=16'h8003;
17'h54e4:	data_out=16'h8001;
17'h54e5:	data_out=16'h8001;
17'h54e6:	data_out=16'h3;
17'h54e7:	data_out=16'h8003;
17'h54e8:	data_out=16'h8001;
17'h54e9:	data_out=16'h8009;
17'h54ea:	data_out=16'h8004;
17'h54eb:	data_out=16'h1;
17'h54ec:	data_out=16'h800f;
17'h54ed:	data_out=16'h3;
17'h54ee:	data_out=16'h0;
17'h54ef:	data_out=16'h8001;
17'h54f0:	data_out=16'h2;
17'h54f1:	data_out=16'h8003;
17'h54f2:	data_out=16'h8011;
17'h54f3:	data_out=16'h8006;
17'h54f4:	data_out=16'h800a;
17'h54f5:	data_out=16'h2;
17'h54f6:	data_out=16'h3;
17'h54f7:	data_out=16'h800d;
17'h54f8:	data_out=16'h8005;
17'h54f9:	data_out=16'h8004;
17'h54fa:	data_out=16'h8005;
17'h54fb:	data_out=16'h6;
17'h54fc:	data_out=16'h6;
17'h54fd:	data_out=16'hd;
17'h54fe:	data_out=16'h7;
17'h54ff:	data_out=16'h800a;
17'h5500:	data_out=16'h80d8;
17'h5501:	data_out=16'h83;
17'h5502:	data_out=16'he0;
17'h5503:	data_out=16'h8071;
17'h5504:	data_out=16'h829a;
17'h5505:	data_out=16'h8068;
17'h5506:	data_out=16'h81d6;
17'h5507:	data_out=16'h826e;
17'h5508:	data_out=16'h801d;
17'h5509:	data_out=16'h81e0;
17'h550a:	data_out=16'h80b9;
17'h550b:	data_out=16'h8062;
17'h550c:	data_out=16'h8170;
17'h550d:	data_out=16'h811e;
17'h550e:	data_out=16'h80c0;
17'h550f:	data_out=16'h80f0;
17'h5510:	data_out=16'h8118;
17'h5511:	data_out=16'h8188;
17'h5512:	data_out=16'h77;
17'h5513:	data_out=16'h81d8;
17'h5514:	data_out=16'h16f;
17'h5515:	data_out=16'h81af;
17'h5516:	data_out=16'h824e;
17'h5517:	data_out=16'h171;
17'h5518:	data_out=16'h8116;
17'h5519:	data_out=16'h38;
17'h551a:	data_out=16'h82ab;
17'h551b:	data_out=16'h15e;
17'h551c:	data_out=16'h3b;
17'h551d:	data_out=16'h1e6;
17'h551e:	data_out=16'h1bc;
17'h551f:	data_out=16'h8209;
17'h5520:	data_out=16'h3df;
17'h5521:	data_out=16'h80c0;
17'h5522:	data_out=16'h225;
17'h5523:	data_out=16'h8329;
17'h5524:	data_out=16'h8328;
17'h5525:	data_out=16'h80f4;
17'h5526:	data_out=16'h8268;
17'h5527:	data_out=16'h2f3;
17'h5528:	data_out=16'h80b5;
17'h5529:	data_out=16'h2f;
17'h552a:	data_out=16'h81e5;
17'h552b:	data_out=16'h169;
17'h552c:	data_out=16'h81b4;
17'h552d:	data_out=16'h823e;
17'h552e:	data_out=16'h80ad;
17'h552f:	data_out=16'h263;
17'h5530:	data_out=16'h8336;
17'h5531:	data_out=16'hac;
17'h5532:	data_out=16'h8343;
17'h5533:	data_out=16'h1b4;
17'h5534:	data_out=16'h81db;
17'h5535:	data_out=16'h811b;
17'h5536:	data_out=16'h121;
17'h5537:	data_out=16'he0;
17'h5538:	data_out=16'h80ff;
17'h5539:	data_out=16'h100;
17'h553a:	data_out=16'h5f;
17'h553b:	data_out=16'h816c;
17'h553c:	data_out=16'h1b9;
17'h553d:	data_out=16'h80d9;
17'h553e:	data_out=16'h80ba;
17'h553f:	data_out=16'h8171;
17'h5540:	data_out=16'h8270;
17'h5541:	data_out=16'h197;
17'h5542:	data_out=16'h814f;
17'h5543:	data_out=16'h815e;
17'h5544:	data_out=16'h81a2;
17'h5545:	data_out=16'h81ba;
17'h5546:	data_out=16'h1de;
17'h5547:	data_out=16'h813a;
17'h5548:	data_out=16'h8023;
17'h5549:	data_out=16'h80f3;
17'h554a:	data_out=16'h8223;
17'h554b:	data_out=16'h80c0;
17'h554c:	data_out=16'h8227;
17'h554d:	data_out=16'h25c;
17'h554e:	data_out=16'h8173;
17'h554f:	data_out=16'h824f;
17'h5550:	data_out=16'h8198;
17'h5551:	data_out=16'h8293;
17'h5552:	data_out=16'h837e;
17'h5553:	data_out=16'h57e;
17'h5554:	data_out=16'h24e;
17'h5555:	data_out=16'h8052;
17'h5556:	data_out=16'h80db;
17'h5557:	data_out=16'h80e3;
17'h5558:	data_out=16'hbd;
17'h5559:	data_out=16'h81a7;
17'h555a:	data_out=16'h237;
17'h555b:	data_out=16'h80a7;
17'h555c:	data_out=16'h1fa;
17'h555d:	data_out=16'h8052;
17'h555e:	data_out=16'h1c5;
17'h555f:	data_out=16'h8009;
17'h5560:	data_out=16'h8405;
17'h5561:	data_out=16'h8217;
17'h5562:	data_out=16'hb0;
17'h5563:	data_out=16'h1ad;
17'h5564:	data_out=16'h8179;
17'h5565:	data_out=16'h80f3;
17'h5566:	data_out=16'hfe;
17'h5567:	data_out=16'h4a;
17'h5568:	data_out=16'h80bd;
17'h5569:	data_out=16'h80d0;
17'h556a:	data_out=16'h80da;
17'h556b:	data_out=16'h820e;
17'h556c:	data_out=16'h16f;
17'h556d:	data_out=16'h1b6;
17'h556e:	data_out=16'h80c9;
17'h556f:	data_out=16'h8109;
17'h5570:	data_out=16'h80c6;
17'h5571:	data_out=16'h81ee;
17'h5572:	data_out=16'h83c6;
17'h5573:	data_out=16'h82fe;
17'h5574:	data_out=16'h833b;
17'h5575:	data_out=16'h818d;
17'h5576:	data_out=16'h69;
17'h5577:	data_out=16'h844f;
17'h5578:	data_out=16'h821d;
17'h5579:	data_out=16'h8168;
17'h557a:	data_out=16'h194;
17'h557b:	data_out=16'h80ae;
17'h557c:	data_out=16'h8034;
17'h557d:	data_out=16'h8203;
17'h557e:	data_out=16'h821f;
17'h557f:	data_out=16'h82fc;
17'h5580:	data_out=16'h82f4;
17'h5581:	data_out=16'h4c9;
17'h5582:	data_out=16'h8506;
17'h5583:	data_out=16'h93;
17'h5584:	data_out=16'h88d0;
17'h5585:	data_out=16'h24b;
17'h5586:	data_out=16'h817e;
17'h5587:	data_out=16'h8810;
17'h5588:	data_out=16'h868c;
17'h5589:	data_out=16'h89ff;
17'h558a:	data_out=16'h84ec;
17'h558b:	data_out=16'h841;
17'h558c:	data_out=16'h89a5;
17'h558d:	data_out=16'h2d2;
17'h558e:	data_out=16'h831e;
17'h558f:	data_out=16'h8354;
17'h5590:	data_out=16'h842f;
17'h5591:	data_out=16'h8650;
17'h5592:	data_out=16'h80c4;
17'h5593:	data_out=16'h81c3;
17'h5594:	data_out=16'h788;
17'h5595:	data_out=16'h845a;
17'h5596:	data_out=16'h8551;
17'h5597:	data_out=16'h91a;
17'h5598:	data_out=16'h8353;
17'h5599:	data_out=16'h811a;
17'h559a:	data_out=16'h8662;
17'h559b:	data_out=16'h9ee;
17'h559c:	data_out=16'h249;
17'h559d:	data_out=16'h360;
17'h559e:	data_out=16'h69f;
17'h559f:	data_out=16'h87d5;
17'h55a0:	data_out=16'ha00;
17'h55a1:	data_out=16'h830f;
17'h55a2:	data_out=16'h8122;
17'h55a3:	data_out=16'h8a00;
17'h55a4:	data_out=16'h8a00;
17'h55a5:	data_out=16'h8891;
17'h55a6:	data_out=16'h8a00;
17'h55a7:	data_out=16'h797;
17'h55a8:	data_out=16'h82eb;
17'h55a9:	data_out=16'h42a;
17'h55aa:	data_out=16'h89c9;
17'h55ab:	data_out=16'h4e2;
17'h55ac:	data_out=16'h84e7;
17'h55ad:	data_out=16'h8750;
17'h55ae:	data_out=16'h845e;
17'h55af:	data_out=16'ha00;
17'h55b0:	data_out=16'h8a00;
17'h55b1:	data_out=16'h7f9;
17'h55b2:	data_out=16'h8a00;
17'h55b3:	data_out=16'h793;
17'h55b4:	data_out=16'hb8;
17'h55b5:	data_out=16'h87fd;
17'h55b6:	data_out=16'h8053;
17'h55b7:	data_out=16'h832b;
17'h55b8:	data_out=16'h35c;
17'h55b9:	data_out=16'h842;
17'h55ba:	data_out=16'h8640;
17'h55bb:	data_out=16'h863f;
17'h55bc:	data_out=16'h258;
17'h55bd:	data_out=16'h8303;
17'h55be:	data_out=16'h82e6;
17'h55bf:	data_out=16'h16d;
17'h55c0:	data_out=16'h8a00;
17'h55c1:	data_out=16'h24a;
17'h55c2:	data_out=16'h87ff;
17'h55c3:	data_out=16'h33;
17'h55c4:	data_out=16'h81a5;
17'h55c5:	data_out=16'h847f;
17'h55c6:	data_out=16'h232;
17'h55c7:	data_out=16'h89fa;
17'h55c8:	data_out=16'h801a;
17'h55c9:	data_out=16'h88de;
17'h55ca:	data_out=16'h87ae;
17'h55cb:	data_out=16'h8100;
17'h55cc:	data_out=16'h8a00;
17'h55cd:	data_out=16'h8038;
17'h55ce:	data_out=16'h84e6;
17'h55cf:	data_out=16'h8a00;
17'h55d0:	data_out=16'h8953;
17'h55d1:	data_out=16'h8698;
17'h55d2:	data_out=16'h8a00;
17'h55d3:	data_out=16'ha00;
17'h55d4:	data_out=16'h933;
17'h55d5:	data_out=16'h83ff;
17'h55d6:	data_out=16'h8a00;
17'h55d7:	data_out=16'h8a00;
17'h55d8:	data_out=16'h85ad;
17'h55d9:	data_out=16'h89ff;
17'h55da:	data_out=16'h9ff;
17'h55db:	data_out=16'h3f;
17'h55dc:	data_out=16'h9c6;
17'h55dd:	data_out=16'h8269;
17'h55de:	data_out=16'h9b1;
17'h55df:	data_out=16'h12d;
17'h55e0:	data_out=16'h8a00;
17'h55e1:	data_out=16'h82b3;
17'h55e2:	data_out=16'h9bc;
17'h55e3:	data_out=16'h823;
17'h55e4:	data_out=16'ha1;
17'h55e5:	data_out=16'hee;
17'h55e6:	data_out=16'h5f;
17'h55e7:	data_out=16'h82ce;
17'h55e8:	data_out=16'h830b;
17'h55e9:	data_out=16'h875e;
17'h55ea:	data_out=16'h832c;
17'h55eb:	data_out=16'h81fd;
17'h55ec:	data_out=16'h820a;
17'h55ed:	data_out=16'h7fe;
17'h55ee:	data_out=16'h832c;
17'h55ef:	data_out=16'h83c6;
17'h55f0:	data_out=16'h8325;
17'h55f1:	data_out=16'h85f4;
17'h55f2:	data_out=16'h88f9;
17'h55f3:	data_out=16'h857c;
17'h55f4:	data_out=16'h8a00;
17'h55f5:	data_out=16'h690;
17'h55f6:	data_out=16'h5b;
17'h55f7:	data_out=16'h8a00;
17'h55f8:	data_out=16'h80d7;
17'h55f9:	data_out=16'h8758;
17'h55fa:	data_out=16'h802;
17'h55fb:	data_out=16'h82d8;
17'h55fc:	data_out=16'h80dc;
17'h55fd:	data_out=16'h1ec;
17'h55fe:	data_out=16'h89ed;
17'h55ff:	data_out=16'h89c2;
17'h5600:	data_out=16'h8a00;
17'h5601:	data_out=16'h89a0;
17'h5602:	data_out=16'h2bd;
17'h5603:	data_out=16'h81a4;
17'h5604:	data_out=16'h3d;
17'h5605:	data_out=16'h9fb;
17'h5606:	data_out=16'ha00;
17'h5607:	data_out=16'h889;
17'h5608:	data_out=16'h88a3;
17'h5609:	data_out=16'h891f;
17'h560a:	data_out=16'h8a00;
17'h560b:	data_out=16'h9fd;
17'h560c:	data_out=16'h8a9;
17'h560d:	data_out=16'h954;
17'h560e:	data_out=16'h82a0;
17'h560f:	data_out=16'h6d1;
17'h5610:	data_out=16'h85b5;
17'h5611:	data_out=16'h39c;
17'h5612:	data_out=16'ha00;
17'h5613:	data_out=16'h340;
17'h5614:	data_out=16'h9ff;
17'h5615:	data_out=16'h8987;
17'h5616:	data_out=16'h8a00;
17'h5617:	data_out=16'h9f7;
17'h5618:	data_out=16'h8244;
17'h5619:	data_out=16'h484;
17'h561a:	data_out=16'h36f;
17'h561b:	data_out=16'h9e5;
17'h561c:	data_out=16'h8259;
17'h561d:	data_out=16'h82ad;
17'h561e:	data_out=16'h9f5;
17'h561f:	data_out=16'h887;
17'h5620:	data_out=16'h9f8;
17'h5621:	data_out=16'h81f1;
17'h5622:	data_out=16'h811d;
17'h5623:	data_out=16'h8a00;
17'h5624:	data_out=16'h8a00;
17'h5625:	data_out=16'h81d8;
17'h5626:	data_out=16'h8a00;
17'h5627:	data_out=16'h89e;
17'h5628:	data_out=16'h8078;
17'h5629:	data_out=16'h2f3;
17'h562a:	data_out=16'h81be;
17'h562b:	data_out=16'ha00;
17'h562c:	data_out=16'h89e2;
17'h562d:	data_out=16'h8a00;
17'h562e:	data_out=16'ha00;
17'h562f:	data_out=16'h9f0;
17'h5630:	data_out=16'h871d;
17'h5631:	data_out=16'h96c;
17'h5632:	data_out=16'h881d;
17'h5633:	data_out=16'ha00;
17'h5634:	data_out=16'h8a00;
17'h5635:	data_out=16'h617;
17'h5636:	data_out=16'h8281;
17'h5637:	data_out=16'h40b;
17'h5638:	data_out=16'h3d6;
17'h5639:	data_out=16'ha00;
17'h563a:	data_out=16'h8c;
17'h563b:	data_out=16'h860e;
17'h563c:	data_out=16'h823b;
17'h563d:	data_out=16'h89fe;
17'h563e:	data_out=16'h806a;
17'h563f:	data_out=16'h9fb;
17'h5640:	data_out=16'h8992;
17'h5641:	data_out=16'h836;
17'h5642:	data_out=16'h88fc;
17'h5643:	data_out=16'ha00;
17'h5644:	data_out=16'h80c0;
17'h5645:	data_out=16'h89b4;
17'h5646:	data_out=16'h850d;
17'h5647:	data_out=16'hde;
17'h5648:	data_out=16'ha00;
17'h5649:	data_out=16'h82ae;
17'h564a:	data_out=16'ha00;
17'h564b:	data_out=16'h868;
17'h564c:	data_out=16'h1ae;
17'h564d:	data_out=16'hb;
17'h564e:	data_out=16'ha00;
17'h564f:	data_out=16'h4b;
17'h5650:	data_out=16'h807e;
17'h5651:	data_out=16'hb5;
17'h5652:	data_out=16'h8a00;
17'h5653:	data_out=16'ha00;
17'h5654:	data_out=16'h52b;
17'h5655:	data_out=16'h84de;
17'h5656:	data_out=16'h8a00;
17'h5657:	data_out=16'h89fb;
17'h5658:	data_out=16'h89e9;
17'h5659:	data_out=16'h89ff;
17'h565a:	data_out=16'h9fe;
17'h565b:	data_out=16'h831e;
17'h565c:	data_out=16'h9d6;
17'h565d:	data_out=16'h83e6;
17'h565e:	data_out=16'h9f1;
17'h565f:	data_out=16'h2a3;
17'h5660:	data_out=16'h8a00;
17'h5661:	data_out=16'h837c;
17'h5662:	data_out=16'h9ee;
17'h5663:	data_out=16'ha00;
17'h5664:	data_out=16'h8335;
17'h5665:	data_out=16'h9f8;
17'h5666:	data_out=16'h90a;
17'h5667:	data_out=16'h536;
17'h5668:	data_out=16'h817f;
17'h5669:	data_out=16'h89fc;
17'h566a:	data_out=16'h8350;
17'h566b:	data_out=16'h42b;
17'h566c:	data_out=16'h8a00;
17'h566d:	data_out=16'ha00;
17'h566e:	data_out=16'h834f;
17'h566f:	data_out=16'h231;
17'h5670:	data_out=16'h82d2;
17'h5671:	data_out=16'ha00;
17'h5672:	data_out=16'h89ff;
17'h5673:	data_out=16'h8569;
17'h5674:	data_out=16'h873d;
17'h5675:	data_out=16'h892;
17'h5676:	data_out=16'h6f7;
17'h5677:	data_out=16'h89f7;
17'h5678:	data_out=16'h99c;
17'h5679:	data_out=16'h935;
17'h567a:	data_out=16'ha00;
17'h567b:	data_out=16'h803e;
17'h567c:	data_out=16'h1d5;
17'h567d:	data_out=16'ha00;
17'h567e:	data_out=16'h89c8;
17'h567f:	data_out=16'h8844;
17'h5680:	data_out=16'h8a00;
17'h5681:	data_out=16'h6c;
17'h5682:	data_out=16'h27f;
17'h5683:	data_out=16'h8a00;
17'h5684:	data_out=16'h8046;
17'h5685:	data_out=16'h7c8;
17'h5686:	data_out=16'h5a7;
17'h5687:	data_out=16'ha00;
17'h5688:	data_out=16'h81a0;
17'h5689:	data_out=16'h88ae;
17'h568a:	data_out=16'h8a00;
17'h568b:	data_out=16'h9fe;
17'h568c:	data_out=16'h9f0;
17'h568d:	data_out=16'h66e;
17'h568e:	data_out=16'h845f;
17'h568f:	data_out=16'h94f;
17'h5690:	data_out=16'h89f3;
17'h5691:	data_out=16'h77a;
17'h5692:	data_out=16'h9fa;
17'h5693:	data_out=16'h89fd;
17'h5694:	data_out=16'h9eb;
17'h5695:	data_out=16'h8a00;
17'h5696:	data_out=16'h8a00;
17'h5697:	data_out=16'h9de;
17'h5698:	data_out=16'h2d4;
17'h5699:	data_out=16'ha00;
17'h569a:	data_out=16'h77;
17'h569b:	data_out=16'h9b8;
17'h569c:	data_out=16'h8818;
17'h569d:	data_out=16'h5fa;
17'h569e:	data_out=16'h9e1;
17'h569f:	data_out=16'ha00;
17'h56a0:	data_out=16'h9eb;
17'h56a1:	data_out=16'h83c8;
17'h56a2:	data_out=16'h8359;
17'h56a3:	data_out=16'h8a00;
17'h56a4:	data_out=16'h8a00;
17'h56a5:	data_out=16'h89fc;
17'h56a6:	data_out=16'h8a00;
17'h56a7:	data_out=16'h9f7;
17'h56a8:	data_out=16'h825f;
17'h56a9:	data_out=16'h82e2;
17'h56aa:	data_out=16'h2fd;
17'h56ab:	data_out=16'ha00;
17'h56ac:	data_out=16'h8a00;
17'h56ad:	data_out=16'h8a00;
17'h56ae:	data_out=16'ha00;
17'h56af:	data_out=16'h9e5;
17'h56b0:	data_out=16'h894b;
17'h56b1:	data_out=16'h9aa;
17'h56b2:	data_out=16'h89f7;
17'h56b3:	data_out=16'h9ff;
17'h56b4:	data_out=16'h8a00;
17'h56b5:	data_out=16'h80c;
17'h56b6:	data_out=16'h88f;
17'h56b7:	data_out=16'h2d6;
17'h56b8:	data_out=16'h9f7;
17'h56b9:	data_out=16'h9fa;
17'h56ba:	data_out=16'h9db;
17'h56bb:	data_out=16'h8433;
17'h56bc:	data_out=16'h87c6;
17'h56bd:	data_out=16'h89fd;
17'h56be:	data_out=16'h822a;
17'h56bf:	data_out=16'h784;
17'h56c0:	data_out=16'h89fc;
17'h56c1:	data_out=16'h7c0;
17'h56c2:	data_out=16'h8a00;
17'h56c3:	data_out=16'h4de;
17'h56c4:	data_out=16'h583;
17'h56c5:	data_out=16'h8a00;
17'h56c6:	data_out=16'h8a00;
17'h56c7:	data_out=16'h11c;
17'h56c8:	data_out=16'ha00;
17'h56c9:	data_out=16'h89ff;
17'h56ca:	data_out=16'ha00;
17'h56cb:	data_out=16'h4e8;
17'h56cc:	data_out=16'h842d;
17'h56cd:	data_out=16'h80f4;
17'h56ce:	data_out=16'ha00;
17'h56cf:	data_out=16'h823e;
17'h56d0:	data_out=16'h8809;
17'h56d1:	data_out=16'h85c4;
17'h56d2:	data_out=16'h8a00;
17'h56d3:	data_out=16'ha00;
17'h56d4:	data_out=16'h9ee;
17'h56d5:	data_out=16'h89f4;
17'h56d6:	data_out=16'h89ff;
17'h56d7:	data_out=16'h89fd;
17'h56d8:	data_out=16'h89f2;
17'h56d9:	data_out=16'h89ff;
17'h56da:	data_out=16'h9f4;
17'h56db:	data_out=16'h173;
17'h56dc:	data_out=16'h9c0;
17'h56dd:	data_out=16'h81bc;
17'h56de:	data_out=16'h9de;
17'h56df:	data_out=16'h9fe;
17'h56e0:	data_out=16'h8a00;
17'h56e1:	data_out=16'h6c;
17'h56e2:	data_out=16'h9d3;
17'h56e3:	data_out=16'ha00;
17'h56e4:	data_out=16'h850f;
17'h56e5:	data_out=16'h808;
17'h56e6:	data_out=16'ha00;
17'h56e7:	data_out=16'h9fc;
17'h56e8:	data_out=16'h8352;
17'h56e9:	data_out=16'h8739;
17'h56ea:	data_out=16'h84e6;
17'h56eb:	data_out=16'h1e2;
17'h56ec:	data_out=16'h8a00;
17'h56ed:	data_out=16'ha00;
17'h56ee:	data_out=16'h84e4;
17'h56ef:	data_out=16'h8856;
17'h56f0:	data_out=16'h8498;
17'h56f1:	data_out=16'h9f6;
17'h56f2:	data_out=16'h8a00;
17'h56f3:	data_out=16'h8a00;
17'h56f4:	data_out=16'h897a;
17'h56f5:	data_out=16'h8222;
17'h56f6:	data_out=16'h9fc;
17'h56f7:	data_out=16'h89f2;
17'h56f8:	data_out=16'h17d;
17'h56f9:	data_out=16'h9c5;
17'h56fa:	data_out=16'h9f6;
17'h56fb:	data_out=16'h81c3;
17'h56fc:	data_out=16'ha00;
17'h56fd:	data_out=16'ha00;
17'h56fe:	data_out=16'h89ee;
17'h56ff:	data_out=16'h8839;
17'h5700:	data_out=16'h8a00;
17'h5701:	data_out=16'h9b0;
17'h5702:	data_out=16'h559;
17'h5703:	data_out=16'h89fd;
17'h5704:	data_out=16'h5af;
17'h5705:	data_out=16'h68f;
17'h5706:	data_out=16'h87eb;
17'h5707:	data_out=16'h9ff;
17'h5708:	data_out=16'h94;
17'h5709:	data_out=16'h89d0;
17'h570a:	data_out=16'h8a00;
17'h570b:	data_out=16'h9fd;
17'h570c:	data_out=16'h402;
17'h570d:	data_out=16'h8441;
17'h570e:	data_out=16'h819c;
17'h570f:	data_out=16'h9ed;
17'h5710:	data_out=16'h8a00;
17'h5711:	data_out=16'h527;
17'h5712:	data_out=16'h9fc;
17'h5713:	data_out=16'h89d4;
17'h5714:	data_out=16'h9f0;
17'h5715:	data_out=16'h8a00;
17'h5716:	data_out=16'h89fd;
17'h5717:	data_out=16'h9e5;
17'h5718:	data_out=16'h705;
17'h5719:	data_out=16'h9fd;
17'h571a:	data_out=16'h9fb;
17'h571b:	data_out=16'h9d7;
17'h571c:	data_out=16'h88cf;
17'h571d:	data_out=16'h58a;
17'h571e:	data_out=16'h9e2;
17'h571f:	data_out=16'ha00;
17'h5720:	data_out=16'h9f7;
17'h5721:	data_out=16'h80d7;
17'h5722:	data_out=16'h48d;
17'h5723:	data_out=16'h8a00;
17'h5724:	data_out=16'h8a00;
17'h5725:	data_out=16'h89fe;
17'h5726:	data_out=16'h8a00;
17'h5727:	data_out=16'h9fa;
17'h5728:	data_out=16'h205;
17'h5729:	data_out=16'h8268;
17'h572a:	data_out=16'h743;
17'h572b:	data_out=16'ha00;
17'h572c:	data_out=16'h89fe;
17'h572d:	data_out=16'h88c0;
17'h572e:	data_out=16'ha00;
17'h572f:	data_out=16'h9f5;
17'h5730:	data_out=16'h8378;
17'h5731:	data_out=16'h8fc;
17'h5732:	data_out=16'h8598;
17'h5733:	data_out=16'h9ff;
17'h5734:	data_out=16'h8860;
17'h5735:	data_out=16'h681;
17'h5736:	data_out=16'h9f4;
17'h5737:	data_out=16'h584;
17'h5738:	data_out=16'h9fd;
17'h5739:	data_out=16'h9fe;
17'h573a:	data_out=16'h437;
17'h573b:	data_out=16'h82ca;
17'h573c:	data_out=16'h868e;
17'h573d:	data_out=16'h89cc;
17'h573e:	data_out=16'h20b;
17'h573f:	data_out=16'h62c;
17'h5740:	data_out=16'h89f9;
17'h5741:	data_out=16'h85a;
17'h5742:	data_out=16'h8a00;
17'h5743:	data_out=16'h851a;
17'h5744:	data_out=16'h44b;
17'h5745:	data_out=16'h8a00;
17'h5746:	data_out=16'hdd;
17'h5747:	data_out=16'h87f5;
17'h5748:	data_out=16'h9ff;
17'h5749:	data_out=16'h89ff;
17'h574a:	data_out=16'ha00;
17'h574b:	data_out=16'h8245;
17'h574c:	data_out=16'h8a00;
17'h574d:	data_out=16'h8d8;
17'h574e:	data_out=16'ha00;
17'h574f:	data_out=16'h89ff;
17'h5750:	data_out=16'h14e;
17'h5751:	data_out=16'h89db;
17'h5752:	data_out=16'h8a00;
17'h5753:	data_out=16'ha00;
17'h5754:	data_out=16'h9fa;
17'h5755:	data_out=16'h89c9;
17'h5756:	data_out=16'h89ff;
17'h5757:	data_out=16'h89eb;
17'h5758:	data_out=16'h89e8;
17'h5759:	data_out=16'h8a00;
17'h575a:	data_out=16'h9fe;
17'h575b:	data_out=16'h892;
17'h575c:	data_out=16'h9d0;
17'h575d:	data_out=16'h78c;
17'h575e:	data_out=16'h9df;
17'h575f:	data_out=16'ha00;
17'h5760:	data_out=16'h89ff;
17'h5761:	data_out=16'h13;
17'h5762:	data_out=16'h8f0;
17'h5763:	data_out=16'ha00;
17'h5764:	data_out=16'h8a00;
17'h5765:	data_out=16'h8549;
17'h5766:	data_out=16'ha00;
17'h5767:	data_out=16'h9fa;
17'h5768:	data_out=16'h8015;
17'h5769:	data_out=16'h8875;
17'h576a:	data_out=16'h8241;
17'h576b:	data_out=16'h8a1;
17'h576c:	data_out=16'h8a00;
17'h576d:	data_out=16'ha00;
17'h576e:	data_out=16'h823e;
17'h576f:	data_out=16'h8229;
17'h5770:	data_out=16'h81e1;
17'h5771:	data_out=16'ha00;
17'h5772:	data_out=16'h8a00;
17'h5773:	data_out=16'h8a00;
17'h5774:	data_out=16'h839a;
17'h5775:	data_out=16'h86c0;
17'h5776:	data_out=16'h9fe;
17'h5777:	data_out=16'h89d6;
17'h5778:	data_out=16'h85f2;
17'h5779:	data_out=16'h9fd;
17'h577a:	data_out=16'ha00;
17'h577b:	data_out=16'h20c;
17'h577c:	data_out=16'ha00;
17'h577d:	data_out=16'ha00;
17'h577e:	data_out=16'h89f7;
17'h577f:	data_out=16'hd7;
17'h5780:	data_out=16'h89e8;
17'h5781:	data_out=16'h9f4;
17'h5782:	data_out=16'h9e2;
17'h5783:	data_out=16'h89f0;
17'h5784:	data_out=16'ha00;
17'h5785:	data_out=16'ha00;
17'h5786:	data_out=16'h8758;
17'h5787:	data_out=16'h9f5;
17'h5788:	data_out=16'h800f;
17'h5789:	data_out=16'h815f;
17'h578a:	data_out=16'h89e7;
17'h578b:	data_out=16'h80c7;
17'h578c:	data_out=16'h81ff;
17'h578d:	data_out=16'h89e9;
17'h578e:	data_out=16'h6f0;
17'h578f:	data_out=16'ha00;
17'h5790:	data_out=16'h2a;
17'h5791:	data_out=16'h9e4;
17'h5792:	data_out=16'h9eb;
17'h5793:	data_out=16'h89ea;
17'h5794:	data_out=16'h829;
17'h5795:	data_out=16'h86b5;
17'h5796:	data_out=16'h89e9;
17'h5797:	data_out=16'h359;
17'h5798:	data_out=16'h9fd;
17'h5799:	data_out=16'h9fa;
17'h579a:	data_out=16'ha00;
17'h579b:	data_out=16'h863;
17'h579c:	data_out=16'h89f1;
17'h579d:	data_out=16'h9f1;
17'h579e:	data_out=16'h9f5;
17'h579f:	data_out=16'ha00;
17'h57a0:	data_out=16'h9da;
17'h57a1:	data_out=16'h74c;
17'h57a2:	data_out=16'ha00;
17'h57a3:	data_out=16'h89ff;
17'h57a4:	data_out=16'h89ff;
17'h57a5:	data_out=16'h855d;
17'h57a6:	data_out=16'h89fe;
17'h57a7:	data_out=16'h9f0;
17'h57a8:	data_out=16'h7d7;
17'h57a9:	data_out=16'h358;
17'h57aa:	data_out=16'ha00;
17'h57ab:	data_out=16'ha00;
17'h57ac:	data_out=16'h89ec;
17'h57ad:	data_out=16'h7ec;
17'h57ae:	data_out=16'ha00;
17'h57af:	data_out=16'ha00;
17'h57b0:	data_out=16'h672;
17'h57b1:	data_out=16'h3a8;
17'h57b2:	data_out=16'h6c6;
17'h57b3:	data_out=16'h9fa;
17'h57b4:	data_out=16'h863d;
17'h57b5:	data_out=16'h7a8;
17'h57b6:	data_out=16'ha00;
17'h57b7:	data_out=16'h9ee;
17'h57b8:	data_out=16'h9fd;
17'h57b9:	data_out=16'h9ee;
17'h57ba:	data_out=16'h9dc;
17'h57bb:	data_out=16'h767;
17'h57bc:	data_out=16'h89ec;
17'h57bd:	data_out=16'h99e;
17'h57be:	data_out=16'h7db;
17'h57bf:	data_out=16'ha00;
17'h57c0:	data_out=16'ha00;
17'h57c1:	data_out=16'h88eb;
17'h57c2:	data_out=16'h89fc;
17'h57c3:	data_out=16'h8702;
17'h57c4:	data_out=16'h4a5;
17'h57c5:	data_out=16'h8738;
17'h57c6:	data_out=16'h441;
17'h57c7:	data_out=16'h9f3;
17'h57c8:	data_out=16'h9f7;
17'h57c9:	data_out=16'h86b6;
17'h57ca:	data_out=16'ha00;
17'h57cb:	data_out=16'h8400;
17'h57cc:	data_out=16'h8386;
17'h57cd:	data_out=16'ha00;
17'h57ce:	data_out=16'ha00;
17'h57cf:	data_out=16'h4ef;
17'h57d0:	data_out=16'h8f2;
17'h57d1:	data_out=16'h89e9;
17'h57d2:	data_out=16'h89fd;
17'h57d3:	data_out=16'ha00;
17'h57d4:	data_out=16'h9ff;
17'h57d5:	data_out=16'h89b1;
17'h57d6:	data_out=16'h89f3;
17'h57d7:	data_out=16'h889a;
17'h57d8:	data_out=16'h89e1;
17'h57d9:	data_out=16'h49;
17'h57da:	data_out=16'h9d8;
17'h57db:	data_out=16'h818d;
17'h57dc:	data_out=16'h967;
17'h57dd:	data_out=16'h9fd;
17'h57de:	data_out=16'h9e9;
17'h57df:	data_out=16'ha00;
17'h57e0:	data_out=16'h89f1;
17'h57e1:	data_out=16'h80a9;
17'h57e2:	data_out=16'h83f5;
17'h57e3:	data_out=16'h9ff;
17'h57e4:	data_out=16'h89f1;
17'h57e5:	data_out=16'h9e8;
17'h57e6:	data_out=16'ha00;
17'h57e7:	data_out=16'h9fc;
17'h57e8:	data_out=16'h784;
17'h57e9:	data_out=16'h89da;
17'h57ea:	data_out=16'h69d;
17'h57eb:	data_out=16'h9f9;
17'h57ec:	data_out=16'h89e0;
17'h57ed:	data_out=16'h9ff;
17'h57ee:	data_out=16'h69d;
17'h57ef:	data_out=16'h87e;
17'h57f0:	data_out=16'h6cb;
17'h57f1:	data_out=16'ha00;
17'h57f2:	data_out=16'h8762;
17'h57f3:	data_out=16'h80f3;
17'h57f4:	data_out=16'h5c4;
17'h57f5:	data_out=16'h89eb;
17'h57f6:	data_out=16'ha00;
17'h57f7:	data_out=16'h8783;
17'h57f8:	data_out=16'h8095;
17'h57f9:	data_out=16'h9fd;
17'h57fa:	data_out=16'h9ff;
17'h57fb:	data_out=16'h7da;
17'h57fc:	data_out=16'ha00;
17'h57fd:	data_out=16'ha00;
17'h57fe:	data_out=16'h89fe;
17'h57ff:	data_out=16'h95a;
17'h5800:	data_out=16'h89de;
17'h5801:	data_out=16'h9fd;
17'h5802:	data_out=16'h9dc;
17'h5803:	data_out=16'h89f4;
17'h5804:	data_out=16'ha00;
17'h5805:	data_out=16'h9ff;
17'h5806:	data_out=16'h89e9;
17'h5807:	data_out=16'h48e;
17'h5808:	data_out=16'h6a6;
17'h5809:	data_out=16'h89fc;
17'h580a:	data_out=16'h89c5;
17'h580b:	data_out=16'h88e4;
17'h580c:	data_out=16'h891a;
17'h580d:	data_out=16'h8a00;
17'h580e:	data_out=16'h9ff;
17'h580f:	data_out=16'ha00;
17'h5810:	data_out=16'h89f4;
17'h5811:	data_out=16'h9fa;
17'h5812:	data_out=16'h9d5;
17'h5813:	data_out=16'h89f6;
17'h5814:	data_out=16'h8465;
17'h5815:	data_out=16'h8831;
17'h5816:	data_out=16'h89f2;
17'h5817:	data_out=16'h895a;
17'h5818:	data_out=16'h9fb;
17'h5819:	data_out=16'ha00;
17'h581a:	data_out=16'ha00;
17'h581b:	data_out=16'ha3;
17'h581c:	data_out=16'h89ef;
17'h581d:	data_out=16'h9f1;
17'h581e:	data_out=16'h535;
17'h581f:	data_out=16'h75e;
17'h5820:	data_out=16'h9e8;
17'h5821:	data_out=16'ha00;
17'h5822:	data_out=16'ha00;
17'h5823:	data_out=16'h89ff;
17'h5824:	data_out=16'h89ff;
17'h5825:	data_out=16'h89f5;
17'h5826:	data_out=16'h89f8;
17'h5827:	data_out=16'h9fe;
17'h5828:	data_out=16'ha00;
17'h5829:	data_out=16'h7ea;
17'h582a:	data_out=16'ha00;
17'h582b:	data_out=16'ha00;
17'h582c:	data_out=16'h89f2;
17'h582d:	data_out=16'ha00;
17'h582e:	data_out=16'ha00;
17'h582f:	data_out=16'h9ff;
17'h5830:	data_out=16'h363;
17'h5831:	data_out=16'h85e0;
17'h5832:	data_out=16'h3b4;
17'h5833:	data_out=16'h9f6;
17'h5834:	data_out=16'h80a6;
17'h5835:	data_out=16'h8d6;
17'h5836:	data_out=16'ha00;
17'h5837:	data_out=16'h9f3;
17'h5838:	data_out=16'h9fe;
17'h5839:	data_out=16'h9cb;
17'h583a:	data_out=16'h332;
17'h583b:	data_out=16'h6e6;
17'h583c:	data_out=16'h898c;
17'h583d:	data_out=16'h97a;
17'h583e:	data_out=16'ha00;
17'h583f:	data_out=16'h9ff;
17'h5840:	data_out=16'ha00;
17'h5841:	data_out=16'h888c;
17'h5842:	data_out=16'h89fc;
17'h5843:	data_out=16'h8572;
17'h5844:	data_out=16'h832c;
17'h5845:	data_out=16'h897b;
17'h5846:	data_out=16'ha00;
17'h5847:	data_out=16'h84c3;
17'h5848:	data_out=16'h803;
17'h5849:	data_out=16'h89f8;
17'h584a:	data_out=16'ha00;
17'h584b:	data_out=16'h89ff;
17'h584c:	data_out=16'h89fd;
17'h584d:	data_out=16'ha00;
17'h584e:	data_out=16'ha00;
17'h584f:	data_out=16'h89fd;
17'h5850:	data_out=16'h1b;
17'h5851:	data_out=16'h89f0;
17'h5852:	data_out=16'h89f4;
17'h5853:	data_out=16'ha00;
17'h5854:	data_out=16'ha00;
17'h5855:	data_out=16'h89e0;
17'h5856:	data_out=16'h89ed;
17'h5857:	data_out=16'h82d0;
17'h5858:	data_out=16'h89f3;
17'h5859:	data_out=16'h3b1;
17'h585a:	data_out=16'h87e1;
17'h585b:	data_out=16'h9fe;
17'h585c:	data_out=16'h8ed;
17'h585d:	data_out=16'ha00;
17'h585e:	data_out=16'h9dd;
17'h585f:	data_out=16'ha00;
17'h5860:	data_out=16'h899a;
17'h5861:	data_out=16'h830c;
17'h5862:	data_out=16'h88f6;
17'h5863:	data_out=16'h9ff;
17'h5864:	data_out=16'h89d4;
17'h5865:	data_out=16'h8666;
17'h5866:	data_out=16'ha00;
17'h5867:	data_out=16'ha00;
17'h5868:	data_out=16'ha00;
17'h5869:	data_out=16'h881a;
17'h586a:	data_out=16'h9ff;
17'h586b:	data_out=16'h85a;
17'h586c:	data_out=16'h2bb;
17'h586d:	data_out=16'h9ff;
17'h586e:	data_out=16'h9ff;
17'h586f:	data_out=16'h8129;
17'h5870:	data_out=16'h9ff;
17'h5871:	data_out=16'ha00;
17'h5872:	data_out=16'h89ba;
17'h5873:	data_out=16'h8582;
17'h5874:	data_out=16'h1bf;
17'h5875:	data_out=16'h89f6;
17'h5876:	data_out=16'ha00;
17'h5877:	data_out=16'h89f2;
17'h5878:	data_out=16'h599;
17'h5879:	data_out=16'ha00;
17'h587a:	data_out=16'h6bf;
17'h587b:	data_out=16'ha00;
17'h587c:	data_out=16'ha00;
17'h587d:	data_out=16'ha00;
17'h587e:	data_out=16'h89fe;
17'h587f:	data_out=16'h841;
17'h5880:	data_out=16'h87a0;
17'h5881:	data_out=16'h5cb;
17'h5882:	data_out=16'h81bb;
17'h5883:	data_out=16'h89e9;
17'h5884:	data_out=16'h9ff;
17'h5885:	data_out=16'h87bc;
17'h5886:	data_out=16'h89d9;
17'h5887:	data_out=16'h8578;
17'h5888:	data_out=16'h9e5;
17'h5889:	data_out=16'h89e8;
17'h588a:	data_out=16'h89e0;
17'h588b:	data_out=16'h88af;
17'h588c:	data_out=16'h89c3;
17'h588d:	data_out=16'h8a00;
17'h588e:	data_out=16'h9fe;
17'h588f:	data_out=16'h80ed;
17'h5890:	data_out=16'h89c1;
17'h5891:	data_out=16'h8996;
17'h5892:	data_out=16'h29d;
17'h5893:	data_out=16'h89f0;
17'h5894:	data_out=16'h88a8;
17'h5895:	data_out=16'h8922;
17'h5896:	data_out=16'h89cb;
17'h5897:	data_out=16'h892f;
17'h5898:	data_out=16'h71e;
17'h5899:	data_out=16'ha00;
17'h589a:	data_out=16'h9ff;
17'h589b:	data_out=16'h89c4;
17'h589c:	data_out=16'h89e5;
17'h589d:	data_out=16'h8777;
17'h589e:	data_out=16'h8870;
17'h589f:	data_out=16'hd6;
17'h58a0:	data_out=16'ha00;
17'h58a1:	data_out=16'h9fe;
17'h58a2:	data_out=16'h8091;
17'h58a3:	data_out=16'h8a00;
17'h58a4:	data_out=16'h8a00;
17'h58a5:	data_out=16'h89c4;
17'h58a6:	data_out=16'h89e1;
17'h58a7:	data_out=16'h9db;
17'h58a8:	data_out=16'h9ff;
17'h58a9:	data_out=16'h9f3;
17'h58aa:	data_out=16'h8293;
17'h58ab:	data_out=16'ha00;
17'h58ac:	data_out=16'h89c6;
17'h58ad:	data_out=16'h8187;
17'h58ae:	data_out=16'ha00;
17'h58af:	data_out=16'h4ce;
17'h58b0:	data_out=16'h842d;
17'h58b1:	data_out=16'h89a3;
17'h58b2:	data_out=16'h84df;
17'h58b3:	data_out=16'h7c;
17'h58b4:	data_out=16'h869a;
17'h58b5:	data_out=16'h89a;
17'h58b6:	data_out=16'ha00;
17'h58b7:	data_out=16'h8425;
17'h58b8:	data_out=16'h8997;
17'h58b9:	data_out=16'h26b;
17'h58ba:	data_out=16'h89c8;
17'h58bb:	data_out=16'h83c5;
17'h58bc:	data_out=16'h8950;
17'h58bd:	data_out=16'h5ac;
17'h58be:	data_out=16'h9ff;
17'h58bf:	data_out=16'h87b7;
17'h58c0:	data_out=16'h806a;
17'h58c1:	data_out=16'h889f;
17'h58c2:	data_out=16'h89ff;
17'h58c3:	data_out=16'h319;
17'h58c4:	data_out=16'h8658;
17'h58c5:	data_out=16'h896c;
17'h58c6:	data_out=16'ha00;
17'h58c7:	data_out=16'h8607;
17'h58c8:	data_out=16'h874a;
17'h58c9:	data_out=16'h89d3;
17'h58ca:	data_out=16'h9fe;
17'h58cb:	data_out=16'h8a00;
17'h58cc:	data_out=16'h89f8;
17'h58cd:	data_out=16'h99a;
17'h58ce:	data_out=16'ha00;
17'h58cf:	data_out=16'h89fb;
17'h58d0:	data_out=16'h898b;
17'h58d1:	data_out=16'h89ee;
17'h58d2:	data_out=16'h89fe;
17'h58d3:	data_out=16'ha00;
17'h58d4:	data_out=16'ha00;
17'h58d5:	data_out=16'h89a1;
17'h58d6:	data_out=16'h89e8;
17'h58d7:	data_out=16'h2d;
17'h58d8:	data_out=16'h89ed;
17'h58d9:	data_out=16'h8913;
17'h58da:	data_out=16'h8999;
17'h58db:	data_out=16'h9ef;
17'h58dc:	data_out=16'h80b0;
17'h58dd:	data_out=16'h4ad;
17'h58de:	data_out=16'h8783;
17'h58df:	data_out=16'ha00;
17'h58e0:	data_out=16'h89de;
17'h58e1:	data_out=16'h86d2;
17'h58e2:	data_out=16'h894a;
17'h58e3:	data_out=16'h1e6;
17'h58e4:	data_out=16'h89db;
17'h58e5:	data_out=16'h875a;
17'h58e6:	data_out=16'ha00;
17'h58e7:	data_out=16'ha00;
17'h58e8:	data_out=16'h9fe;
17'h58e9:	data_out=16'h84b7;
17'h58ea:	data_out=16'h9fd;
17'h58eb:	data_out=16'h8853;
17'h58ec:	data_out=16'h832e;
17'h58ed:	data_out=16'h1b8;
17'h58ee:	data_out=16'h9fd;
17'h58ef:	data_out=16'h852e;
17'h58f0:	data_out=16'h9fe;
17'h58f1:	data_out=16'ha00;
17'h58f2:	data_out=16'h8982;
17'h58f3:	data_out=16'h8881;
17'h58f4:	data_out=16'h8559;
17'h58f5:	data_out=16'h89fc;
17'h58f6:	data_out=16'ha00;
17'h58f7:	data_out=16'h89c2;
17'h58f8:	data_out=16'ha00;
17'h58f9:	data_out=16'ha00;
17'h58fa:	data_out=16'h87f5;
17'h58fb:	data_out=16'h9ff;
17'h58fc:	data_out=16'ha00;
17'h58fd:	data_out=16'ha00;
17'h58fe:	data_out=16'h89ea;
17'h58ff:	data_out=16'h7e5;
17'h5900:	data_out=16'h9fe;
17'h5901:	data_out=16'h77d;
17'h5902:	data_out=16'h8963;
17'h5903:	data_out=16'h8908;
17'h5904:	data_out=16'h159;
17'h5905:	data_out=16'h87ed;
17'h5906:	data_out=16'h8a00;
17'h5907:	data_out=16'h89f2;
17'h5908:	data_out=16'h9e3;
17'h5909:	data_out=16'h8a00;
17'h590a:	data_out=16'h89ba;
17'h590b:	data_out=16'h8840;
17'h590c:	data_out=16'h89ea;
17'h590d:	data_out=16'h89db;
17'h590e:	data_out=16'h8ab;
17'h590f:	data_out=16'h88de;
17'h5910:	data_out=16'h89e1;
17'h5911:	data_out=16'h89e8;
17'h5912:	data_out=16'h889d;
17'h5913:	data_out=16'h898f;
17'h5914:	data_out=16'h8719;
17'h5915:	data_out=16'h8617;
17'h5916:	data_out=16'h8867;
17'h5917:	data_out=16'h8743;
17'h5918:	data_out=16'h10e;
17'h5919:	data_out=16'h9f6;
17'h591a:	data_out=16'h8146;
17'h591b:	data_out=16'h897a;
17'h591c:	data_out=16'h87eb;
17'h591d:	data_out=16'h8763;
17'h591e:	data_out=16'h8777;
17'h591f:	data_out=16'h851c;
17'h5920:	data_out=16'h9ef;
17'h5921:	data_out=16'h821;
17'h5922:	data_out=16'h897d;
17'h5923:	data_out=16'h8a00;
17'h5924:	data_out=16'h8a00;
17'h5925:	data_out=16'h89fe;
17'h5926:	data_out=16'h89d3;
17'h5927:	data_out=16'h3d0;
17'h5928:	data_out=16'h75f;
17'h5929:	data_out=16'ha00;
17'h592a:	data_out=16'h86bf;
17'h592b:	data_out=16'ha00;
17'h592c:	data_out=16'h8830;
17'h592d:	data_out=16'h88f4;
17'h592e:	data_out=16'h8173;
17'h592f:	data_out=16'h864c;
17'h5930:	data_out=16'h881a;
17'h5931:	data_out=16'h358;
17'h5932:	data_out=16'h8966;
17'h5933:	data_out=16'h8704;
17'h5934:	data_out=16'h970;
17'h5935:	data_out=16'h8251;
17'h5936:	data_out=16'ha00;
17'h5937:	data_out=16'h890d;
17'h5938:	data_out=16'h89ed;
17'h5939:	data_out=16'h8628;
17'h593a:	data_out=16'h89f5;
17'h593b:	data_out=16'h88d2;
17'h593c:	data_out=16'h87bf;
17'h593d:	data_out=16'h5bb;
17'h593e:	data_out=16'h759;
17'h593f:	data_out=16'h87ef;
17'h5940:	data_out=16'h86ae;
17'h5941:	data_out=16'h86b8;
17'h5942:	data_out=16'h8a00;
17'h5943:	data_out=16'ha00;
17'h5944:	data_out=16'h81da;
17'h5945:	data_out=16'h87ca;
17'h5946:	data_out=16'ha00;
17'h5947:	data_out=16'h89e4;
17'h5948:	data_out=16'h89fc;
17'h5949:	data_out=16'h89fe;
17'h594a:	data_out=16'h9eb;
17'h594b:	data_out=16'h8a00;
17'h594c:	data_out=16'h8a00;
17'h594d:	data_out=16'h899c;
17'h594e:	data_out=16'ha00;
17'h594f:	data_out=16'h8a00;
17'h5950:	data_out=16'h88db;
17'h5951:	data_out=16'h89ac;
17'h5952:	data_out=16'h8a00;
17'h5953:	data_out=16'h9c0;
17'h5954:	data_out=16'h969;
17'h5955:	data_out=16'h892e;
17'h5956:	data_out=16'h89e4;
17'h5957:	data_out=16'h85db;
17'h5958:	data_out=16'h89cc;
17'h5959:	data_out=16'h8976;
17'h595a:	data_out=16'h8961;
17'h595b:	data_out=16'h9e0;
17'h595c:	data_out=16'h89c8;
17'h595d:	data_out=16'h835e;
17'h595e:	data_out=16'h8793;
17'h595f:	data_out=16'h698;
17'h5960:	data_out=16'h89d8;
17'h5961:	data_out=16'h88af;
17'h5962:	data_out=16'h87d8;
17'h5963:	data_out=16'h86db;
17'h5964:	data_out=16'h882b;
17'h5965:	data_out=16'h8865;
17'h5966:	data_out=16'ha00;
17'h5967:	data_out=16'ha00;
17'h5968:	data_out=16'h7c0;
17'h5969:	data_out=16'hd9;
17'h596a:	data_out=16'h903;
17'h596b:	data_out=16'h87d3;
17'h596c:	data_out=16'ha00;
17'h596d:	data_out=16'h86e0;
17'h596e:	data_out=16'h900;
17'h596f:	data_out=16'h84e5;
17'h5970:	data_out=16'h8d0;
17'h5971:	data_out=16'h8096;
17'h5972:	data_out=16'h8964;
17'h5973:	data_out=16'h87c0;
17'h5974:	data_out=16'h8948;
17'h5975:	data_out=16'h89ed;
17'h5976:	data_out=16'ha00;
17'h5977:	data_out=16'h89f9;
17'h5978:	data_out=16'ha00;
17'h5979:	data_out=16'ha00;
17'h597a:	data_out=16'h86ec;
17'h597b:	data_out=16'h755;
17'h597c:	data_out=16'h9f9;
17'h597d:	data_out=16'h8df;
17'h597e:	data_out=16'h89e5;
17'h597f:	data_out=16'h141;
17'h5980:	data_out=16'h9fc;
17'h5981:	data_out=16'h9f7;
17'h5982:	data_out=16'h89aa;
17'h5983:	data_out=16'h87f0;
17'h5984:	data_out=16'h84ed;
17'h5985:	data_out=16'h885e;
17'h5986:	data_out=16'h8a00;
17'h5987:	data_out=16'h8a00;
17'h5988:	data_out=16'h9bf;
17'h5989:	data_out=16'h8a00;
17'h598a:	data_out=16'h898f;
17'h598b:	data_out=16'h878c;
17'h598c:	data_out=16'h8a00;
17'h598d:	data_out=16'h89e0;
17'h598e:	data_out=16'h5c8;
17'h598f:	data_out=16'h89a0;
17'h5990:	data_out=16'h89c8;
17'h5991:	data_out=16'h89f9;
17'h5992:	data_out=16'h89de;
17'h5993:	data_out=16'h89a4;
17'h5994:	data_out=16'h872e;
17'h5995:	data_out=16'hcc;
17'h5996:	data_out=16'h88c2;
17'h5997:	data_out=16'h8780;
17'h5998:	data_out=16'h8964;
17'h5999:	data_out=16'h9fa;
17'h599a:	data_out=16'h84b5;
17'h599b:	data_out=16'h8998;
17'h599c:	data_out=16'h8627;
17'h599d:	data_out=16'h8763;
17'h599e:	data_out=16'h87ea;
17'h599f:	data_out=16'h8767;
17'h59a0:	data_out=16'h9e3;
17'h59a1:	data_out=16'h4db;
17'h59a2:	data_out=16'h895c;
17'h59a3:	data_out=16'h8a00;
17'h59a4:	data_out=16'h8a00;
17'h59a5:	data_out=16'h89f7;
17'h59a6:	data_out=16'h89c8;
17'h59a7:	data_out=16'h181;
17'h59a8:	data_out=16'h3a9;
17'h59a9:	data_out=16'ha00;
17'h59aa:	data_out=16'h880a;
17'h59ab:	data_out=16'ha00;
17'h59ac:	data_out=16'h886d;
17'h59ad:	data_out=16'h88a2;
17'h59ae:	data_out=16'h896e;
17'h59af:	data_out=16'h871e;
17'h59b0:	data_out=16'h8340;
17'h59b1:	data_out=16'h7ea;
17'h59b2:	data_out=16'h8908;
17'h59b3:	data_out=16'h8800;
17'h59b4:	data_out=16'ha00;
17'h59b5:	data_out=16'h89cb;
17'h59b6:	data_out=16'h9f4;
17'h59b7:	data_out=16'h8967;
17'h59b8:	data_out=16'h89f8;
17'h59b9:	data_out=16'h880e;
17'h59ba:	data_out=16'h89f4;
17'h59bb:	data_out=16'h89ec;
17'h59bc:	data_out=16'h8565;
17'h59bd:	data_out=16'h9f9;
17'h59be:	data_out=16'h3a1;
17'h59bf:	data_out=16'h885c;
17'h59c0:	data_out=16'h8829;
17'h59c1:	data_out=16'h2a2;
17'h59c2:	data_out=16'h8a00;
17'h59c3:	data_out=16'ha00;
17'h59c4:	data_out=16'h30a;
17'h59c5:	data_out=16'h80fb;
17'h59c6:	data_out=16'ha00;
17'h59c7:	data_out=16'h89e8;
17'h59c8:	data_out=16'h8a00;
17'h59c9:	data_out=16'h89e1;
17'h59ca:	data_out=16'h8527;
17'h59cb:	data_out=16'h8a00;
17'h59cc:	data_out=16'h8a00;
17'h59cd:	data_out=16'h896e;
17'h59ce:	data_out=16'h4af;
17'h59cf:	data_out=16'h8a00;
17'h59d0:	data_out=16'h885c;
17'h59d1:	data_out=16'h89bf;
17'h59d2:	data_out=16'h8a00;
17'h59d3:	data_out=16'h8900;
17'h59d4:	data_out=16'h576;
17'h59d5:	data_out=16'h8941;
17'h59d6:	data_out=16'h8226;
17'h59d7:	data_out=16'h8693;
17'h59d8:	data_out=16'h89de;
17'h59d9:	data_out=16'h895f;
17'h59da:	data_out=16'h89d0;
17'h59db:	data_out=16'h9d4;
17'h59dc:	data_out=16'h89e3;
17'h59dd:	data_out=16'h84c4;
17'h59de:	data_out=16'h8762;
17'h59df:	data_out=16'h8960;
17'h59e0:	data_out=16'h89da;
17'h59e1:	data_out=16'h88fd;
17'h59e2:	data_out=16'h8748;
17'h59e3:	data_out=16'h883e;
17'h59e4:	data_out=16'h807e;
17'h59e5:	data_out=16'h8837;
17'h59e6:	data_out=16'ha00;
17'h59e7:	data_out=16'ha00;
17'h59e8:	data_out=16'h442;
17'h59e9:	data_out=16'h53;
17'h59ea:	data_out=16'h64d;
17'h59eb:	data_out=16'h886c;
17'h59ec:	data_out=16'ha00;
17'h59ed:	data_out=16'h8831;
17'h59ee:	data_out=16'h64a;
17'h59ef:	data_out=16'h851a;
17'h59f0:	data_out=16'h607;
17'h59f1:	data_out=16'h896f;
17'h59f2:	data_out=16'h8949;
17'h59f3:	data_out=16'h875d;
17'h59f4:	data_out=16'h848d;
17'h59f5:	data_out=16'h89f8;
17'h59f6:	data_out=16'ha00;
17'h59f7:	data_out=16'h89ef;
17'h59f8:	data_out=16'h9ff;
17'h59f9:	data_out=16'ha00;
17'h59fa:	data_out=16'h87a0;
17'h59fb:	data_out=16'h39b;
17'h59fc:	data_out=16'h838e;
17'h59fd:	data_out=16'h840e;
17'h59fe:	data_out=16'h89e3;
17'h59ff:	data_out=16'h87d6;
17'h5a00:	data_out=16'h99b;
17'h5a01:	data_out=16'h9d2;
17'h5a02:	data_out=16'h89ca;
17'h5a03:	data_out=16'h8865;
17'h5a04:	data_out=16'h8152;
17'h5a05:	data_out=16'h88bf;
17'h5a06:	data_out=16'h8a00;
17'h5a07:	data_out=16'h8a00;
17'h5a08:	data_out=16'h825;
17'h5a09:	data_out=16'h8a00;
17'h5a0a:	data_out=16'hfc;
17'h5a0b:	data_out=16'h9c1;
17'h5a0c:	data_out=16'h8a00;
17'h5a0d:	data_out=16'h8a00;
17'h5a0e:	data_out=16'h503;
17'h5a0f:	data_out=16'h89d4;
17'h5a10:	data_out=16'h8793;
17'h5a11:	data_out=16'h89fd;
17'h5a12:	data_out=16'h89fa;
17'h5a13:	data_out=16'h898c;
17'h5a14:	data_out=16'h85d5;
17'h5a15:	data_out=16'h84ab;
17'h5a16:	data_out=16'h89bc;
17'h5a17:	data_out=16'h8758;
17'h5a18:	data_out=16'h89fc;
17'h5a19:	data_out=16'ha00;
17'h5a1a:	data_out=16'h8680;
17'h5a1b:	data_out=16'h88e6;
17'h5a1c:	data_out=16'h84b4;
17'h5a1d:	data_out=16'h8467;
17'h5a1e:	data_out=16'h8793;
17'h5a1f:	data_out=16'h867a;
17'h5a20:	data_out=16'h9bd;
17'h5a21:	data_out=16'h3f7;
17'h5a22:	data_out=16'h87fd;
17'h5a23:	data_out=16'h8a00;
17'h5a24:	data_out=16'h8a00;
17'h5a25:	data_out=16'h89d3;
17'h5a26:	data_out=16'h89fb;
17'h5a27:	data_out=16'h67b;
17'h5a28:	data_out=16'h360;
17'h5a29:	data_out=16'ha00;
17'h5a2a:	data_out=16'h8806;
17'h5a2b:	data_out=16'h9f8;
17'h5a2c:	data_out=16'h897d;
17'h5a2d:	data_out=16'h894b;
17'h5a2e:	data_out=16'h8907;
17'h5a2f:	data_out=16'h876a;
17'h5a30:	data_out=16'h21f;
17'h5a31:	data_out=16'h1cc;
17'h5a32:	data_out=16'h8991;
17'h5a33:	data_out=16'h86c7;
17'h5a34:	data_out=16'h94f;
17'h5a35:	data_out=16'h870a;
17'h5a36:	data_out=16'h8030;
17'h5a37:	data_out=16'h8936;
17'h5a38:	data_out=16'h8a00;
17'h5a39:	data_out=16'h8742;
17'h5a3a:	data_out=16'h89f6;
17'h5a3b:	data_out=16'h89fb;
17'h5a3c:	data_out=16'h9f4;
17'h5a3d:	data_out=16'h9cc;
17'h5a3e:	data_out=16'h360;
17'h5a3f:	data_out=16'h88bb;
17'h5a40:	data_out=16'h8923;
17'h5a41:	data_out=16'h9d5;
17'h5a42:	data_out=16'h8a00;
17'h5a43:	data_out=16'ha00;
17'h5a44:	data_out=16'h11d;
17'h5a45:	data_out=16'h858c;
17'h5a46:	data_out=16'ha00;
17'h5a47:	data_out=16'h89f7;
17'h5a48:	data_out=16'h8a00;
17'h5a49:	data_out=16'h89b1;
17'h5a4a:	data_out=16'h87ba;
17'h5a4b:	data_out=16'h8a00;
17'h5a4c:	data_out=16'h89ec;
17'h5a4d:	data_out=16'h883c;
17'h5a4e:	data_out=16'h8137;
17'h5a4f:	data_out=16'h8a00;
17'h5a50:	data_out=16'h885f;
17'h5a51:	data_out=16'h89f8;
17'h5a52:	data_out=16'h8a00;
17'h5a53:	data_out=16'h88fb;
17'h5a54:	data_out=16'h8355;
17'h5a55:	data_out=16'h8844;
17'h5a56:	data_out=16'h27f;
17'h5a57:	data_out=16'h86ea;
17'h5a58:	data_out=16'h89f7;
17'h5a59:	data_out=16'h8949;
17'h5a5a:	data_out=16'h89e6;
17'h5a5b:	data_out=16'h91a;
17'h5a5c:	data_out=16'h89fc;
17'h5a5d:	data_out=16'h8540;
17'h5a5e:	data_out=16'h86b3;
17'h5a5f:	data_out=16'h89bf;
17'h5a60:	data_out=16'h8a00;
17'h5a61:	data_out=16'h89a6;
17'h5a62:	data_out=16'h85cb;
17'h5a63:	data_out=16'h878e;
17'h5a64:	data_out=16'h2fa;
17'h5a65:	data_out=16'h82b1;
17'h5a66:	data_out=16'h9fb;
17'h5a67:	data_out=16'ha00;
17'h5a68:	data_out=16'h37c;
17'h5a69:	data_out=16'h84e3;
17'h5a6a:	data_out=16'h5a9;
17'h5a6b:	data_out=16'h882b;
17'h5a6c:	data_out=16'h9e8;
17'h5a6d:	data_out=16'h8768;
17'h5a6e:	data_out=16'h5a6;
17'h5a6f:	data_out=16'h86e8;
17'h5a70:	data_out=16'h558;
17'h5a71:	data_out=16'h8995;
17'h5a72:	data_out=16'h8908;
17'h5a73:	data_out=16'h878e;
17'h5a74:	data_out=16'h81e1;
17'h5a75:	data_out=16'h89ff;
17'h5a76:	data_out=16'h9ff;
17'h5a77:	data_out=16'h89f9;
17'h5a78:	data_out=16'h9ff;
17'h5a79:	data_out=16'h9fd;
17'h5a7a:	data_out=16'h86e3;
17'h5a7b:	data_out=16'h35b;
17'h5a7c:	data_out=16'h89fa;
17'h5a7d:	data_out=16'h850a;
17'h5a7e:	data_out=16'h89b7;
17'h5a7f:	data_out=16'h8995;
17'h5a80:	data_out=16'h996;
17'h5a81:	data_out=16'h9ed;
17'h5a82:	data_out=16'h89bd;
17'h5a83:	data_out=16'h88e4;
17'h5a84:	data_out=16'h870d;
17'h5a85:	data_out=16'h8776;
17'h5a86:	data_out=16'h8a00;
17'h5a87:	data_out=16'h8a00;
17'h5a88:	data_out=16'h701;
17'h5a89:	data_out=16'h89fc;
17'h5a8a:	data_out=16'h9cc;
17'h5a8b:	data_out=16'h9b0;
17'h5a8c:	data_out=16'h8a00;
17'h5a8d:	data_out=16'h8a00;
17'h5a8e:	data_out=16'h570;
17'h5a8f:	data_out=16'h89e5;
17'h5a90:	data_out=16'h8203;
17'h5a91:	data_out=16'h80e0;
17'h5a92:	data_out=16'h8a00;
17'h5a93:	data_out=16'h88f1;
17'h5a94:	data_out=16'h82bc;
17'h5a95:	data_out=16'h888c;
17'h5a96:	data_out=16'h89cc;
17'h5a97:	data_out=16'h84e0;
17'h5a98:	data_out=16'h89ff;
17'h5a99:	data_out=16'ha00;
17'h5a9a:	data_out=16'h85d0;
17'h5a9b:	data_out=16'h8596;
17'h5a9c:	data_out=16'h803a;
17'h5a9d:	data_out=16'h537;
17'h5a9e:	data_out=16'h870c;
17'h5a9f:	data_out=16'h85cd;
17'h5aa0:	data_out=16'h841b;
17'h5aa1:	data_out=16'h44e;
17'h5aa2:	data_out=16'h885a;
17'h5aa3:	data_out=16'h89ff;
17'h5aa4:	data_out=16'h89ff;
17'h5aa5:	data_out=16'h8964;
17'h5aa6:	data_out=16'h230;
17'h5aa7:	data_out=16'h835;
17'h5aa8:	data_out=16'h47a;
17'h5aa9:	data_out=16'ha00;
17'h5aaa:	data_out=16'h882c;
17'h5aab:	data_out=16'h9ec;
17'h5aac:	data_out=16'h89a5;
17'h5aad:	data_out=16'h89e0;
17'h5aae:	data_out=16'h88de;
17'h5aaf:	data_out=16'h8775;
17'h5ab0:	data_out=16'h812f;
17'h5ab1:	data_out=16'h9d7;
17'h5ab2:	data_out=16'h8987;
17'h5ab3:	data_out=16'h855e;
17'h5ab4:	data_out=16'h9c2;
17'h5ab5:	data_out=16'h340;
17'h5ab6:	data_out=16'h84da;
17'h5ab7:	data_out=16'h886a;
17'h5ab8:	data_out=16'h8a00;
17'h5ab9:	data_out=16'h86ad;
17'h5aba:	data_out=16'h89f7;
17'h5abb:	data_out=16'h89db;
17'h5abc:	data_out=16'ha00;
17'h5abd:	data_out=16'h829f;
17'h5abe:	data_out=16'h485;
17'h5abf:	data_out=16'h8772;
17'h5ac0:	data_out=16'h8954;
17'h5ac1:	data_out=16'h9dd;
17'h5ac2:	data_out=16'h8a00;
17'h5ac3:	data_out=16'ha00;
17'h5ac4:	data_out=16'h9d7;
17'h5ac5:	data_out=16'h88bb;
17'h5ac6:	data_out=16'h9f4;
17'h5ac7:	data_out=16'h89ff;
17'h5ac8:	data_out=16'h8a00;
17'h5ac9:	data_out=16'h8918;
17'h5aca:	data_out=16'h885d;
17'h5acb:	data_out=16'h8a00;
17'h5acc:	data_out=16'h8a00;
17'h5acd:	data_out=16'h8927;
17'h5ace:	data_out=16'h87d0;
17'h5acf:	data_out=16'h8a00;
17'h5ad0:	data_out=16'h8929;
17'h5ad1:	data_out=16'h89f1;
17'h5ad2:	data_out=16'h8a00;
17'h5ad3:	data_out=16'h86f0;
17'h5ad4:	data_out=16'h875c;
17'h5ad5:	data_out=16'h8635;
17'h5ad6:	data_out=16'h6c5;
17'h5ad7:	data_out=16'h866b;
17'h5ad8:	data_out=16'h8964;
17'h5ad9:	data_out=16'h891e;
17'h5ada:	data_out=16'h896b;
17'h5adb:	data_out=16'h9e1;
17'h5adc:	data_out=16'h8799;
17'h5add:	data_out=16'h869d;
17'h5ade:	data_out=16'h8631;
17'h5adf:	data_out=16'h89f3;
17'h5ae0:	data_out=16'h89f5;
17'h5ae1:	data_out=16'h8901;
17'h5ae2:	data_out=16'h80ce;
17'h5ae3:	data_out=16'h85da;
17'h5ae4:	data_out=16'h9a8;
17'h5ae5:	data_out=16'h9ff;
17'h5ae6:	data_out=16'h9fd;
17'h5ae7:	data_out=16'ha00;
17'h5ae8:	data_out=16'h407;
17'h5ae9:	data_out=16'h8302;
17'h5aea:	data_out=16'h629;
17'h5aeb:	data_out=16'h8680;
17'h5aec:	data_out=16'h82c4;
17'h5aed:	data_out=16'h85cd;
17'h5aee:	data_out=16'h626;
17'h5aef:	data_out=16'h8692;
17'h5af0:	data_out=16'h5d1;
17'h5af1:	data_out=16'h89cd;
17'h5af2:	data_out=16'h8843;
17'h5af3:	data_out=16'h867a;
17'h5af4:	data_out=16'h85c3;
17'h5af5:	data_out=16'h89bd;
17'h5af6:	data_out=16'h9f6;
17'h5af7:	data_out=16'h89f6;
17'h5af8:	data_out=16'ha00;
17'h5af9:	data_out=16'h9f1;
17'h5afa:	data_out=16'h847c;
17'h5afb:	data_out=16'h483;
17'h5afc:	data_out=16'h89fb;
17'h5afd:	data_out=16'h85c3;
17'h5afe:	data_out=16'h8941;
17'h5aff:	data_out=16'h89c0;
17'h5b00:	data_out=16'h152;
17'h5b01:	data_out=16'h9f2;
17'h5b02:	data_out=16'h8905;
17'h5b03:	data_out=16'h8947;
17'h5b04:	data_out=16'h8a9;
17'h5b05:	data_out=16'h86d0;
17'h5b06:	data_out=16'h8a00;
17'h5b07:	data_out=16'h8a00;
17'h5b08:	data_out=16'h5f9;
17'h5b09:	data_out=16'h89ce;
17'h5b0a:	data_out=16'h9ea;
17'h5b0b:	data_out=16'h9e2;
17'h5b0c:	data_out=16'h8a00;
17'h5b0d:	data_out=16'h8a00;
17'h5b0e:	data_out=16'h9ff;
17'h5b0f:	data_out=16'h89a9;
17'h5b10:	data_out=16'h9f7;
17'h5b11:	data_out=16'h9fb;
17'h5b12:	data_out=16'h8a00;
17'h5b13:	data_out=16'h88c7;
17'h5b14:	data_out=16'h81bd;
17'h5b15:	data_out=16'h88b8;
17'h5b16:	data_out=16'h89d8;
17'h5b17:	data_out=16'h8528;
17'h5b18:	data_out=16'h8a00;
17'h5b19:	data_out=16'ha00;
17'h5b1a:	data_out=16'h8598;
17'h5b1b:	data_out=16'h545;
17'h5b1c:	data_out=16'h9db;
17'h5b1d:	data_out=16'h357;
17'h5b1e:	data_out=16'h86da;
17'h5b1f:	data_out=16'h86dd;
17'h5b20:	data_out=16'h84fd;
17'h5b21:	data_out=16'h9ff;
17'h5b22:	data_out=16'h84a3;
17'h5b23:	data_out=16'h89fa;
17'h5b24:	data_out=16'h89f9;
17'h5b25:	data_out=16'h88c0;
17'h5b26:	data_out=16'h989;
17'h5b27:	data_out=16'h9f8;
17'h5b28:	data_out=16'ha00;
17'h5b29:	data_out=16'ha00;
17'h5b2a:	data_out=16'h86a2;
17'h5b2b:	data_out=16'h9f1;
17'h5b2c:	data_out=16'h89b7;
17'h5b2d:	data_out=16'h8997;
17'h5b2e:	data_out=16'h86d1;
17'h5b2f:	data_out=16'h8704;
17'h5b30:	data_out=16'h3ea;
17'h5b31:	data_out=16'h9eb;
17'h5b32:	data_out=16'h81a7;
17'h5b33:	data_out=16'h8690;
17'h5b34:	data_out=16'h4d2;
17'h5b35:	data_out=16'h7c2;
17'h5b36:	data_out=16'h8234;
17'h5b37:	data_out=16'h8601;
17'h5b38:	data_out=16'h89f1;
17'h5b39:	data_out=16'h8864;
17'h5b3a:	data_out=16'h8983;
17'h5b3b:	data_out=16'h89b8;
17'h5b3c:	data_out=16'ha00;
17'h5b3d:	data_out=16'h162;
17'h5b3e:	data_out=16'ha00;
17'h5b3f:	data_out=16'h86cf;
17'h5b40:	data_out=16'h87fc;
17'h5b41:	data_out=16'h9ee;
17'h5b42:	data_out=16'h89fa;
17'h5b43:	data_out=16'ha00;
17'h5b44:	data_out=16'h9f7;
17'h5b45:	data_out=16'h88cd;
17'h5b46:	data_out=16'h9fd;
17'h5b47:	data_out=16'h89f7;
17'h5b48:	data_out=16'h89f1;
17'h5b49:	data_out=16'h8812;
17'h5b4a:	data_out=16'h88a9;
17'h5b4b:	data_out=16'h8a00;
17'h5b4c:	data_out=16'h8a00;
17'h5b4d:	data_out=16'h8729;
17'h5b4e:	data_out=16'h809f;
17'h5b4f:	data_out=16'h89ff;
17'h5b50:	data_out=16'h8982;
17'h5b51:	data_out=16'h89fe;
17'h5b52:	data_out=16'h8a00;
17'h5b53:	data_out=16'h80cf;
17'h5b54:	data_out=16'h8724;
17'h5b55:	data_out=16'h8479;
17'h5b56:	data_out=16'h9c3;
17'h5b57:	data_out=16'h66;
17'h5b58:	data_out=16'h9b7;
17'h5b59:	data_out=16'h8777;
17'h5b5a:	data_out=16'h88b8;
17'h5b5b:	data_out=16'h9f8;
17'h5b5c:	data_out=16'h849d;
17'h5b5d:	data_out=16'h8642;
17'h5b5e:	data_out=16'h84e8;
17'h5b5f:	data_out=16'h89ed;
17'h5b60:	data_out=16'h14;
17'h5b61:	data_out=16'h837e;
17'h5b62:	data_out=16'h831;
17'h5b63:	data_out=16'h86d1;
17'h5b64:	data_out=16'h9a5;
17'h5b65:	data_out=16'ha00;
17'h5b66:	data_out=16'h9f9;
17'h5b67:	data_out=16'ha00;
17'h5b68:	data_out=16'h9ff;
17'h5b69:	data_out=16'h342;
17'h5b6a:	data_out=16'h9ff;
17'h5b6b:	data_out=16'h8637;
17'h5b6c:	data_out=16'h84ff;
17'h5b6d:	data_out=16'h86c4;
17'h5b6e:	data_out=16'h9ff;
17'h5b6f:	data_out=16'h8688;
17'h5b70:	data_out=16'h9ff;
17'h5b71:	data_out=16'h89d3;
17'h5b72:	data_out=16'h85e5;
17'h5b73:	data_out=16'h84e6;
17'h5b74:	data_out=16'h807f;
17'h5b75:	data_out=16'h8786;
17'h5b76:	data_out=16'h9e8;
17'h5b77:	data_out=16'h89a6;
17'h5b78:	data_out=16'h9fe;
17'h5b79:	data_out=16'h9e0;
17'h5b7a:	data_out=16'h845b;
17'h5b7b:	data_out=16'ha00;
17'h5b7c:	data_out=16'h8a00;
17'h5b7d:	data_out=16'h8889;
17'h5b7e:	data_out=16'h628;
17'h5b7f:	data_out=16'h89de;
17'h5b80:	data_out=16'h8319;
17'h5b81:	data_out=16'h9f7;
17'h5b82:	data_out=16'h88b2;
17'h5b83:	data_out=16'h8954;
17'h5b84:	data_out=16'h600;
17'h5b85:	data_out=16'h879e;
17'h5b86:	data_out=16'h89fe;
17'h5b87:	data_out=16'h8a00;
17'h5b88:	data_out=16'h8483;
17'h5b89:	data_out=16'h89a2;
17'h5b8a:	data_out=16'h9fe;
17'h5b8b:	data_out=16'h9fe;
17'h5b8c:	data_out=16'h89ed;
17'h5b8d:	data_out=16'h8a00;
17'h5b8e:	data_out=16'ha00;
17'h5b8f:	data_out=16'h8961;
17'h5b90:	data_out=16'h6ce;
17'h5b91:	data_out=16'h9ff;
17'h5b92:	data_out=16'h8a00;
17'h5b93:	data_out=16'h8724;
17'h5b94:	data_out=16'h8441;
17'h5b95:	data_out=16'h8985;
17'h5b96:	data_out=16'h89e9;
17'h5b97:	data_out=16'h86bb;
17'h5b98:	data_out=16'h8a00;
17'h5b99:	data_out=16'ha00;
17'h5b9a:	data_out=16'h85cc;
17'h5b9b:	data_out=16'h9fe;
17'h5b9c:	data_out=16'h9ce;
17'h5b9d:	data_out=16'h9f5;
17'h5b9e:	data_out=16'h87d8;
17'h5b9f:	data_out=16'h886b;
17'h5ba0:	data_out=16'h852d;
17'h5ba1:	data_out=16'ha00;
17'h5ba2:	data_out=16'h8270;
17'h5ba3:	data_out=16'h89e6;
17'h5ba4:	data_out=16'h89e5;
17'h5ba5:	data_out=16'h8838;
17'h5ba6:	data_out=16'h9be;
17'h5ba7:	data_out=16'h9f9;
17'h5ba8:	data_out=16'ha00;
17'h5ba9:	data_out=16'ha00;
17'h5baa:	data_out=16'h849a;
17'h5bab:	data_out=16'h9e2;
17'h5bac:	data_out=16'h89db;
17'h5bad:	data_out=16'h818e;
17'h5bae:	data_out=16'h841c;
17'h5baf:	data_out=16'h866e;
17'h5bb0:	data_out=16'ha0;
17'h5bb1:	data_out=16'h9fb;
17'h5bb2:	data_out=16'hb5;
17'h5bb3:	data_out=16'h88e2;
17'h5bb4:	data_out=16'h868;
17'h5bb5:	data_out=16'h41e;
17'h5bb6:	data_out=16'h80fe;
17'h5bb7:	data_out=16'h665;
17'h5bb8:	data_out=16'h89b7;
17'h5bb9:	data_out=16'h8973;
17'h5bba:	data_out=16'h89a8;
17'h5bbb:	data_out=16'h895b;
17'h5bbc:	data_out=16'h9fe;
17'h5bbd:	data_out=16'h82dd;
17'h5bbe:	data_out=16'ha00;
17'h5bbf:	data_out=16'h87a2;
17'h5bc0:	data_out=16'h86ff;
17'h5bc1:	data_out=16'h9f0;
17'h5bc2:	data_out=16'h89c1;
17'h5bc3:	data_out=16'ha00;
17'h5bc4:	data_out=16'h826a;
17'h5bc5:	data_out=16'h89a1;
17'h5bc6:	data_out=16'h9fb;
17'h5bc7:	data_out=16'h89fb;
17'h5bc8:	data_out=16'h89d6;
17'h5bc9:	data_out=16'h8784;
17'h5bca:	data_out=16'h8884;
17'h5bcb:	data_out=16'h89ee;
17'h5bcc:	data_out=16'h89fb;
17'h5bcd:	data_out=16'h8519;
17'h5bce:	data_out=16'h81bf;
17'h5bcf:	data_out=16'h89ea;
17'h5bd0:	data_out=16'h89a7;
17'h5bd1:	data_out=16'h8a00;
17'h5bd2:	data_out=16'h89f1;
17'h5bd3:	data_out=16'h39d;
17'h5bd4:	data_out=16'h867c;
17'h5bd5:	data_out=16'h84ed;
17'h5bd6:	data_out=16'h9e9;
17'h5bd7:	data_out=16'h80a3;
17'h5bd8:	data_out=16'h9c4;
17'h5bd9:	data_out=16'h8668;
17'h5bda:	data_out=16'h88fa;
17'h5bdb:	data_out=16'h9fc;
17'h5bdc:	data_out=16'h815a;
17'h5bdd:	data_out=16'h8576;
17'h5bde:	data_out=16'h8427;
17'h5bdf:	data_out=16'h89e7;
17'h5be0:	data_out=16'h2f2;
17'h5be1:	data_out=16'h2d2;
17'h5be2:	data_out=16'ha00;
17'h5be3:	data_out=16'h88b5;
17'h5be4:	data_out=16'h9dd;
17'h5be5:	data_out=16'ha00;
17'h5be6:	data_out=16'h9f5;
17'h5be7:	data_out=16'h9f9;
17'h5be8:	data_out=16'ha00;
17'h5be9:	data_out=16'h882b;
17'h5bea:	data_out=16'ha00;
17'h5beb:	data_out=16'h867c;
17'h5bec:	data_out=16'h87e0;
17'h5bed:	data_out=16'h88b7;
17'h5bee:	data_out=16'ha00;
17'h5bef:	data_out=16'h877f;
17'h5bf0:	data_out=16'ha00;
17'h5bf1:	data_out=16'h89b1;
17'h5bf2:	data_out=16'h82bf;
17'h5bf3:	data_out=16'h2cc;
17'h5bf4:	data_out=16'h8304;
17'h5bf5:	data_out=16'h9bf;
17'h5bf6:	data_out=16'h9e6;
17'h5bf7:	data_out=16'h8953;
17'h5bf8:	data_out=16'ha00;
17'h5bf9:	data_out=16'h311;
17'h5bfa:	data_out=16'h8648;
17'h5bfb:	data_out=16'ha00;
17'h5bfc:	data_out=16'h8a00;
17'h5bfd:	data_out=16'h8949;
17'h5bfe:	data_out=16'h2b2;
17'h5bff:	data_out=16'h89ee;
17'h5c00:	data_out=16'h862c;
17'h5c01:	data_out=16'h9e0;
17'h5c02:	data_out=16'h45b;
17'h5c03:	data_out=16'h8969;
17'h5c04:	data_out=16'h8374;
17'h5c05:	data_out=16'h89fb;
17'h5c06:	data_out=16'h89ef;
17'h5c07:	data_out=16'h8a00;
17'h5c08:	data_out=16'h8060;
17'h5c09:	data_out=16'h895c;
17'h5c0a:	data_out=16'h9cd;
17'h5c0b:	data_out=16'ha00;
17'h5c0c:	data_out=16'h89e7;
17'h5c0d:	data_out=16'h8a00;
17'h5c0e:	data_out=16'ha00;
17'h5c0f:	data_out=16'h87bb;
17'h5c10:	data_out=16'h99c;
17'h5c11:	data_out=16'ha00;
17'h5c12:	data_out=16'h8a00;
17'h5c13:	data_out=16'h8791;
17'h5c14:	data_out=16'h8757;
17'h5c15:	data_out=16'h89f7;
17'h5c16:	data_out=16'h8a00;
17'h5c17:	data_out=16'h8949;
17'h5c18:	data_out=16'h8a00;
17'h5c19:	data_out=16'ha00;
17'h5c1a:	data_out=16'h88cd;
17'h5c1b:	data_out=16'h9ff;
17'h5c1c:	data_out=16'h256;
17'h5c1d:	data_out=16'h9dc;
17'h5c1e:	data_out=16'h88a9;
17'h5c1f:	data_out=16'h8930;
17'h5c20:	data_out=16'h8380;
17'h5c21:	data_out=16'ha00;
17'h5c22:	data_out=16'h5c1;
17'h5c23:	data_out=16'h8437;
17'h5c24:	data_out=16'h8437;
17'h5c25:	data_out=16'h864b;
17'h5c26:	data_out=16'h9c2;
17'h5c27:	data_out=16'h9fa;
17'h5c28:	data_out=16'ha00;
17'h5c29:	data_out=16'h9f0;
17'h5c2a:	data_out=16'hbd;
17'h5c2b:	data_out=16'h9f5;
17'h5c2c:	data_out=16'h8a00;
17'h5c2d:	data_out=16'h81f6;
17'h5c2e:	data_out=16'h8008;
17'h5c2f:	data_out=16'h84f5;
17'h5c30:	data_out=16'h89fc;
17'h5c31:	data_out=16'h53c;
17'h5c32:	data_out=16'h86bc;
17'h5c33:	data_out=16'h8972;
17'h5c34:	data_out=16'h383;
17'h5c35:	data_out=16'h8004;
17'h5c36:	data_out=16'h4c7;
17'h5c37:	data_out=16'h9f1;
17'h5c38:	data_out=16'h89a0;
17'h5c39:	data_out=16'h899c;
17'h5c3a:	data_out=16'h88ff;
17'h5c3b:	data_out=16'h8771;
17'h5c3c:	data_out=16'h9dd;
17'h5c3d:	data_out=16'h835e;
17'h5c3e:	data_out=16'ha00;
17'h5c3f:	data_out=16'h89fb;
17'h5c40:	data_out=16'h8665;
17'h5c41:	data_out=16'h9ed;
17'h5c42:	data_out=16'h8151;
17'h5c43:	data_out=16'ha00;
17'h5c44:	data_out=16'h838a;
17'h5c45:	data_out=16'h89fb;
17'h5c46:	data_out=16'h9dc;
17'h5c47:	data_out=16'h89e0;
17'h5c48:	data_out=16'h89cf;
17'h5c49:	data_out=16'h856a;
17'h5c4a:	data_out=16'h8446;
17'h5c4b:	data_out=16'h89f9;
17'h5c4c:	data_out=16'h89f1;
17'h5c4d:	data_out=16'h201;
17'h5c4e:	data_out=16'h81f7;
17'h5c4f:	data_out=16'h896f;
17'h5c50:	data_out=16'h89e6;
17'h5c51:	data_out=16'h8a00;
17'h5c52:	data_out=16'h8872;
17'h5c53:	data_out=16'h9f9;
17'h5c54:	data_out=16'h81ae;
17'h5c55:	data_out=16'h858e;
17'h5c56:	data_out=16'h66a;
17'h5c57:	data_out=16'h331;
17'h5c58:	data_out=16'h88af;
17'h5c59:	data_out=16'h86a1;
17'h5c5a:	data_out=16'h898a;
17'h5c5b:	data_out=16'h3f8;
17'h5c5c:	data_out=16'h8892;
17'h5c5d:	data_out=16'h835b;
17'h5c5e:	data_out=16'h8340;
17'h5c5f:	data_out=16'h89f7;
17'h5c60:	data_out=16'h6fd;
17'h5c61:	data_out=16'h85dd;
17'h5c62:	data_out=16'ha00;
17'h5c63:	data_out=16'h8963;
17'h5c64:	data_out=16'h9b0;
17'h5c65:	data_out=16'h8387;
17'h5c66:	data_out=16'h9f9;
17'h5c67:	data_out=16'h9e8;
17'h5c68:	data_out=16'ha00;
17'h5c69:	data_out=16'h85e7;
17'h5c6a:	data_out=16'ha00;
17'h5c6b:	data_out=16'h8967;
17'h5c6c:	data_out=16'h89ff;
17'h5c6d:	data_out=16'h8966;
17'h5c6e:	data_out=16'ha00;
17'h5c6f:	data_out=16'h89eb;
17'h5c70:	data_out=16'ha00;
17'h5c71:	data_out=16'h89d9;
17'h5c72:	data_out=16'h863e;
17'h5c73:	data_out=16'h84c3;
17'h5c74:	data_out=16'h8a00;
17'h5c75:	data_out=16'h811b;
17'h5c76:	data_out=16'h9f8;
17'h5c77:	data_out=16'h873a;
17'h5c78:	data_out=16'ha00;
17'h5c79:	data_out=16'h8612;
17'h5c7a:	data_out=16'h87fa;
17'h5c7b:	data_out=16'ha00;
17'h5c7c:	data_out=16'h8a00;
17'h5c7d:	data_out=16'h89a8;
17'h5c7e:	data_out=16'h9fd;
17'h5c7f:	data_out=16'h8a00;
17'h5c80:	data_out=16'h87bd;
17'h5c81:	data_out=16'h7fe;
17'h5c82:	data_out=16'h9d1;
17'h5c83:	data_out=16'h899b;
17'h5c84:	data_out=16'h43;
17'h5c85:	data_out=16'h89d7;
17'h5c86:	data_out=16'h8a00;
17'h5c87:	data_out=16'h8a00;
17'h5c88:	data_out=16'h8119;
17'h5c89:	data_out=16'h874f;
17'h5c8a:	data_out=16'h9e7;
17'h5c8b:	data_out=16'ha00;
17'h5c8c:	data_out=16'h83be;
17'h5c8d:	data_out=16'h8a00;
17'h5c8e:	data_out=16'ha00;
17'h5c8f:	data_out=16'h8399;
17'h5c90:	data_out=16'h8282;
17'h5c91:	data_out=16'ha00;
17'h5c92:	data_out=16'h8a00;
17'h5c93:	data_out=16'h8915;
17'h5c94:	data_out=16'h8999;
17'h5c95:	data_out=16'h89ec;
17'h5c96:	data_out=16'h89e9;
17'h5c97:	data_out=16'h89aa;
17'h5c98:	data_out=16'h8a00;
17'h5c99:	data_out=16'h9fc;
17'h5c9a:	data_out=16'h88a8;
17'h5c9b:	data_out=16'h81a;
17'h5c9c:	data_out=16'h89bd;
17'h5c9d:	data_out=16'h9ea;
17'h5c9e:	data_out=16'h88ff;
17'h5c9f:	data_out=16'h89ad;
17'h5ca0:	data_out=16'h81d5;
17'h5ca1:	data_out=16'ha00;
17'h5ca2:	data_out=16'h8104;
17'h5ca3:	data_out=16'h9d5;
17'h5ca4:	data_out=16'h9d2;
17'h5ca5:	data_out=16'h82ce;
17'h5ca6:	data_out=16'h9ca;
17'h5ca7:	data_out=16'h9cd;
17'h5ca8:	data_out=16'ha00;
17'h5ca9:	data_out=16'h9e9;
17'h5caa:	data_out=16'h9a1;
17'h5cab:	data_out=16'h9e2;
17'h5cac:	data_out=16'h89e9;
17'h5cad:	data_out=16'h87e4;
17'h5cae:	data_out=16'h45e;
17'h5caf:	data_out=16'h8356;
17'h5cb0:	data_out=16'h8a00;
17'h5cb1:	data_out=16'h39e;
17'h5cb2:	data_out=16'h82f6;
17'h5cb3:	data_out=16'h89ca;
17'h5cb4:	data_out=16'h847c;
17'h5cb5:	data_out=16'h5b8;
17'h5cb6:	data_out=16'h64d;
17'h5cb7:	data_out=16'h9ef;
17'h5cb8:	data_out=16'h898d;
17'h5cb9:	data_out=16'h89ce;
17'h5cba:	data_out=16'h8543;
17'h5cbb:	data_out=16'h86;
17'h5cbc:	data_out=16'h9f1;
17'h5cbd:	data_out=16'h812b;
17'h5cbe:	data_out=16'ha00;
17'h5cbf:	data_out=16'h89d9;
17'h5cc0:	data_out=16'h81d2;
17'h5cc1:	data_out=16'h99b;
17'h5cc2:	data_out=16'h8476;
17'h5cc3:	data_out=16'ha00;
17'h5cc4:	data_out=16'h819b;
17'h5cc5:	data_out=16'h89ef;
17'h5cc6:	data_out=16'h9cb;
17'h5cc7:	data_out=16'h89fc;
17'h5cc8:	data_out=16'h89f4;
17'h5cc9:	data_out=16'h8157;
17'h5cca:	data_out=16'h2b;
17'h5ccb:	data_out=16'h8583;
17'h5ccc:	data_out=16'h886b;
17'h5ccd:	data_out=16'h8397;
17'h5cce:	data_out=16'h8232;
17'h5ccf:	data_out=16'h8305;
17'h5cd0:	data_out=16'h89eb;
17'h5cd1:	data_out=16'h8a00;
17'h5cd2:	data_out=16'h974;
17'h5cd3:	data_out=16'h9e7;
17'h5cd4:	data_out=16'h181;
17'h5cd5:	data_out=16'h85a9;
17'h5cd6:	data_out=16'h645;
17'h5cd7:	data_out=16'h9ed;
17'h5cd8:	data_out=16'h89b0;
17'h5cd9:	data_out=16'h8226;
17'h5cda:	data_out=16'h89d4;
17'h5cdb:	data_out=16'h80fc;
17'h5cdc:	data_out=16'h89ab;
17'h5cdd:	data_out=16'hc7;
17'h5cde:	data_out=16'h8182;
17'h5cdf:	data_out=16'h8988;
17'h5ce0:	data_out=16'h9af;
17'h5ce1:	data_out=16'h8384;
17'h5ce2:	data_out=16'ha00;
17'h5ce3:	data_out=16'h89c1;
17'h5ce4:	data_out=16'h935;
17'h5ce5:	data_out=16'h83c6;
17'h5ce6:	data_out=16'h9e4;
17'h5ce7:	data_out=16'h3d2;
17'h5ce8:	data_out=16'ha00;
17'h5ce9:	data_out=16'h8702;
17'h5cea:	data_out=16'ha00;
17'h5ceb:	data_out=16'h891c;
17'h5cec:	data_out=16'h8976;
17'h5ced:	data_out=16'h89c3;
17'h5cee:	data_out=16'ha00;
17'h5cef:	data_out=16'h89fc;
17'h5cf0:	data_out=16'ha00;
17'h5cf1:	data_out=16'h89b1;
17'h5cf2:	data_out=16'h85d8;
17'h5cf3:	data_out=16'h83fc;
17'h5cf4:	data_out=16'h8a00;
17'h5cf5:	data_out=16'h8629;
17'h5cf6:	data_out=16'h9d3;
17'h5cf7:	data_out=16'h834a;
17'h5cf8:	data_out=16'ha00;
17'h5cf9:	data_out=16'h8a00;
17'h5cfa:	data_out=16'h89b2;
17'h5cfb:	data_out=16'ha00;
17'h5cfc:	data_out=16'h8a00;
17'h5cfd:	data_out=16'h89cd;
17'h5cfe:	data_out=16'h3f2;
17'h5cff:	data_out=16'h8a00;
17'h5d00:	data_out=16'h8740;
17'h5d01:	data_out=16'h516;
17'h5d02:	data_out=16'h52e;
17'h5d03:	data_out=16'h89ad;
17'h5d04:	data_out=16'h50b;
17'h5d05:	data_out=16'h88ed;
17'h5d06:	data_out=16'h8a00;
17'h5d07:	data_out=16'h865d;
17'h5d08:	data_out=16'h8312;
17'h5d09:	data_out=16'h89cf;
17'h5d0a:	data_out=16'h9ff;
17'h5d0b:	data_out=16'ha00;
17'h5d0c:	data_out=16'h84f4;
17'h5d0d:	data_out=16'h8a00;
17'h5d0e:	data_out=16'ha00;
17'h5d0f:	data_out=16'h849f;
17'h5d10:	data_out=16'h891b;
17'h5d11:	data_out=16'ha00;
17'h5d12:	data_out=16'h8a00;
17'h5d13:	data_out=16'h857a;
17'h5d14:	data_out=16'h89b7;
17'h5d15:	data_out=16'h886b;
17'h5d16:	data_out=16'h8998;
17'h5d17:	data_out=16'h89ca;
17'h5d18:	data_out=16'h8a00;
17'h5d19:	data_out=16'h9f7;
17'h5d1a:	data_out=16'h86a3;
17'h5d1b:	data_out=16'ha00;
17'h5d1c:	data_out=16'h89cc;
17'h5d1d:	data_out=16'h8a2;
17'h5d1e:	data_out=16'h88cc;
17'h5d1f:	data_out=16'h89f7;
17'h5d20:	data_out=16'h154;
17'h5d21:	data_out=16'h9ff;
17'h5d22:	data_out=16'h884e;
17'h5d23:	data_out=16'ha00;
17'h5d24:	data_out=16'ha00;
17'h5d25:	data_out=16'h844e;
17'h5d26:	data_out=16'h9eb;
17'h5d27:	data_out=16'h5fc;
17'h5d28:	data_out=16'h9fe;
17'h5d29:	data_out=16'h7f7;
17'h5d2a:	data_out=16'h700;
17'h5d2b:	data_out=16'h82eb;
17'h5d2c:	data_out=16'h89df;
17'h5d2d:	data_out=16'h88fd;
17'h5d2e:	data_out=16'h80d3;
17'h5d2f:	data_out=16'h82b9;
17'h5d30:	data_out=16'h8a00;
17'h5d31:	data_out=16'h9ff;
17'h5d32:	data_out=16'h8345;
17'h5d33:	data_out=16'h89db;
17'h5d34:	data_out=16'h89eb;
17'h5d35:	data_out=16'h9bb;
17'h5d36:	data_out=16'h4ce;
17'h5d37:	data_out=16'h9ee;
17'h5d38:	data_out=16'h89dd;
17'h5d39:	data_out=16'h89db;
17'h5d3a:	data_out=16'h85bc;
17'h5d3b:	data_out=16'h9d8;
17'h5d3c:	data_out=16'ha00;
17'h5d3d:	data_out=16'h17e;
17'h5d3e:	data_out=16'h9fe;
17'h5d3f:	data_out=16'h88f6;
17'h5d40:	data_out=16'h7be;
17'h5d41:	data_out=16'h16d;
17'h5d42:	data_out=16'h89f7;
17'h5d43:	data_out=16'ha00;
17'h5d44:	data_out=16'h9ef;
17'h5d45:	data_out=16'h887e;
17'h5d46:	data_out=16'h87a0;
17'h5d47:	data_out=16'h89fc;
17'h5d48:	data_out=16'h89fb;
17'h5d49:	data_out=16'h814c;
17'h5d4a:	data_out=16'h58b;
17'h5d4b:	data_out=16'h881d;
17'h5d4c:	data_out=16'h89f4;
17'h5d4d:	data_out=16'h8958;
17'h5d4e:	data_out=16'h83f7;
17'h5d4f:	data_out=16'h83a6;
17'h5d50:	data_out=16'h89f1;
17'h5d51:	data_out=16'h89f0;
17'h5d52:	data_out=16'h984;
17'h5d53:	data_out=16'h791;
17'h5d54:	data_out=16'h138;
17'h5d55:	data_out=16'h5d5;
17'h5d56:	data_out=16'h8290;
17'h5d57:	data_out=16'hf;
17'h5d58:	data_out=16'h89b9;
17'h5d59:	data_out=16'h80c4;
17'h5d5a:	data_out=16'h89f2;
17'h5d5b:	data_out=16'h4a3;
17'h5d5c:	data_out=16'h890b;
17'h5d5d:	data_out=16'h807f;
17'h5d5e:	data_out=16'h8141;
17'h5d5f:	data_out=16'h89fe;
17'h5d60:	data_out=16'h2b2;
17'h5d61:	data_out=16'h9d2;
17'h5d62:	data_out=16'ha00;
17'h5d63:	data_out=16'h89e1;
17'h5d64:	data_out=16'h8473;
17'h5d65:	data_out=16'h84b3;
17'h5d66:	data_out=16'h9e0;
17'h5d67:	data_out=16'h8214;
17'h5d68:	data_out=16'h9fe;
17'h5d69:	data_out=16'h88b2;
17'h5d6a:	data_out=16'ha00;
17'h5d6b:	data_out=16'h84cf;
17'h5d6c:	data_out=16'h89c5;
17'h5d6d:	data_out=16'h89e0;
17'h5d6e:	data_out=16'ha00;
17'h5d6f:	data_out=16'h89ce;
17'h5d70:	data_out=16'ha00;
17'h5d71:	data_out=16'h8a00;
17'h5d72:	data_out=16'h86aa;
17'h5d73:	data_out=16'h84c2;
17'h5d74:	data_out=16'h8a00;
17'h5d75:	data_out=16'h9e4;
17'h5d76:	data_out=16'h9bf;
17'h5d77:	data_out=16'h85cc;
17'h5d78:	data_out=16'h9ff;
17'h5d79:	data_out=16'h8a00;
17'h5d7a:	data_out=16'h89d4;
17'h5d7b:	data_out=16'h9fe;
17'h5d7c:	data_out=16'h8a00;
17'h5d7d:	data_out=16'h89e8;
17'h5d7e:	data_out=16'h5da;
17'h5d7f:	data_out=16'h89ff;
17'h5d80:	data_out=16'h89d2;
17'h5d81:	data_out=16'h8567;
17'h5d82:	data_out=16'h876c;
17'h5d83:	data_out=16'h89d4;
17'h5d84:	data_out=16'h6e8;
17'h5d85:	data_out=16'h366;
17'h5d86:	data_out=16'h8a00;
17'h5d87:	data_out=16'h8442;
17'h5d88:	data_out=16'h89c4;
17'h5d89:	data_out=16'h8935;
17'h5d8a:	data_out=16'h9fd;
17'h5d8b:	data_out=16'h81a1;
17'h5d8c:	data_out=16'h89e0;
17'h5d8d:	data_out=16'h8a00;
17'h5d8e:	data_out=16'ha00;
17'h5d8f:	data_out=16'h80bb;
17'h5d90:	data_out=16'h89c3;
17'h5d91:	data_out=16'ha00;
17'h5d92:	data_out=16'h8a00;
17'h5d93:	data_out=16'h13e;
17'h5d94:	data_out=16'h89d6;
17'h5d95:	data_out=16'h87ce;
17'h5d96:	data_out=16'h8852;
17'h5d97:	data_out=16'h89f7;
17'h5d98:	data_out=16'h89f6;
17'h5d99:	data_out=16'h9f4;
17'h5d9a:	data_out=16'h87b2;
17'h5d9b:	data_out=16'h31b;
17'h5d9c:	data_out=16'h89ee;
17'h5d9d:	data_out=16'h13c;
17'h5d9e:	data_out=16'h884c;
17'h5d9f:	data_out=16'h89fc;
17'h5da0:	data_out=16'hf;
17'h5da1:	data_out=16'ha00;
17'h5da2:	data_out=16'h89af;
17'h5da3:	data_out=16'ha00;
17'h5da4:	data_out=16'ha00;
17'h5da5:	data_out=16'h84f9;
17'h5da6:	data_out=16'h8591;
17'h5da7:	data_out=16'h82c1;
17'h5da8:	data_out=16'h9ff;
17'h5da9:	data_out=16'h75d;
17'h5daa:	data_out=16'h728;
17'h5dab:	data_out=16'h89b0;
17'h5dac:	data_out=16'h88a1;
17'h5dad:	data_out=16'h898b;
17'h5dae:	data_out=16'h8397;
17'h5daf:	data_out=16'h8923;
17'h5db0:	data_out=16'h8a00;
17'h5db1:	data_out=16'h9f4;
17'h5db2:	data_out=16'h8794;
17'h5db3:	data_out=16'h89fb;
17'h5db4:	data_out=16'h89f1;
17'h5db5:	data_out=16'h5dc;
17'h5db6:	data_out=16'h8290;
17'h5db7:	data_out=16'h8023;
17'h5db8:	data_out=16'h89f5;
17'h5db9:	data_out=16'h89f7;
17'h5dba:	data_out=16'h844b;
17'h5dbb:	data_out=16'h9da;
17'h5dbc:	data_out=16'h223;
17'h5dbd:	data_out=16'h25;
17'h5dbe:	data_out=16'h9ff;
17'h5dbf:	data_out=16'h346;
17'h5dc0:	data_out=16'h9f4;
17'h5dc1:	data_out=16'h8a00;
17'h5dc2:	data_out=16'h89e1;
17'h5dc3:	data_out=16'ha00;
17'h5dc4:	data_out=16'h9ec;
17'h5dc5:	data_out=16'h87c3;
17'h5dc6:	data_out=16'h88e7;
17'h5dc7:	data_out=16'h88b5;
17'h5dc8:	data_out=16'h89fb;
17'h5dc9:	data_out=16'h8329;
17'h5dca:	data_out=16'h478;
17'h5dcb:	data_out=16'h89e5;
17'h5dcc:	data_out=16'h8894;
17'h5dcd:	data_out=16'h89ad;
17'h5dce:	data_out=16'h8a00;
17'h5dcf:	data_out=16'h812f;
17'h5dd0:	data_out=16'h89f3;
17'h5dd1:	data_out=16'h80f2;
17'h5dd2:	data_out=16'h9ae;
17'h5dd3:	data_out=16'h8367;
17'h5dd4:	data_out=16'h8390;
17'h5dd5:	data_out=16'h923;
17'h5dd6:	data_out=16'h89a7;
17'h5dd7:	data_out=16'h37;
17'h5dd8:	data_out=16'h89e4;
17'h5dd9:	data_out=16'h80b1;
17'h5dda:	data_out=16'h8a00;
17'h5ddb:	data_out=16'h9aa;
17'h5ddc:	data_out=16'h89e6;
17'h5ddd:	data_out=16'h8576;
17'h5dde:	data_out=16'h86ed;
17'h5ddf:	data_out=16'h89ac;
17'h5de0:	data_out=16'h818f;
17'h5de1:	data_out=16'h972;
17'h5de2:	data_out=16'h5b;
17'h5de3:	data_out=16'h89fe;
17'h5de4:	data_out=16'h89d6;
17'h5de5:	data_out=16'h8398;
17'h5de6:	data_out=16'h9dd;
17'h5de7:	data_out=16'h80d0;
17'h5de8:	data_out=16'ha00;
17'h5de9:	data_out=16'h89be;
17'h5dea:	data_out=16'ha00;
17'h5deb:	data_out=16'h80a1;
17'h5dec:	data_out=16'h89e0;
17'h5ded:	data_out=16'h89fc;
17'h5dee:	data_out=16'ha00;
17'h5def:	data_out=16'h85a7;
17'h5df0:	data_out=16'ha00;
17'h5df1:	data_out=16'h81c6;
17'h5df2:	data_out=16'h88c7;
17'h5df3:	data_out=16'h87ac;
17'h5df4:	data_out=16'h8a00;
17'h5df5:	data_out=16'h31d;
17'h5df6:	data_out=16'h878c;
17'h5df7:	data_out=16'h8956;
17'h5df8:	data_out=16'h9e7;
17'h5df9:	data_out=16'h8a00;
17'h5dfa:	data_out=16'h89ee;
17'h5dfb:	data_out=16'h9ff;
17'h5dfc:	data_out=16'h89fb;
17'h5dfd:	data_out=16'h89d8;
17'h5dfe:	data_out=16'h68b;
17'h5dff:	data_out=16'h89ff;
17'h5e00:	data_out=16'h8965;
17'h5e01:	data_out=16'h8240;
17'h5e02:	data_out=16'h895f;
17'h5e03:	data_out=16'h8963;
17'h5e04:	data_out=16'h80c8;
17'h5e05:	data_out=16'h926;
17'h5e06:	data_out=16'h8a00;
17'h5e07:	data_out=16'h8665;
17'h5e08:	data_out=16'h8987;
17'h5e09:	data_out=16'h89f0;
17'h5e0a:	data_out=16'h7b6;
17'h5e0b:	data_out=16'h887f;
17'h5e0c:	data_out=16'h89b3;
17'h5e0d:	data_out=16'h89ea;
17'h5e0e:	data_out=16'h9fc;
17'h5e0f:	data_out=16'h84a7;
17'h5e10:	data_out=16'h89f2;
17'h5e11:	data_out=16'ha00;
17'h5e12:	data_out=16'h88d0;
17'h5e13:	data_out=16'h4eb;
17'h5e14:	data_out=16'h89eb;
17'h5e15:	data_out=16'h880;
17'h5e16:	data_out=16'h65c;
17'h5e17:	data_out=16'h89fa;
17'h5e18:	data_out=16'h86e6;
17'h5e19:	data_out=16'h8ed;
17'h5e1a:	data_out=16'h86af;
17'h5e1b:	data_out=16'h8742;
17'h5e1c:	data_out=16'h89ca;
17'h5e1d:	data_out=16'h83ba;
17'h5e1e:	data_out=16'h8928;
17'h5e1f:	data_out=16'h89ff;
17'h5e20:	data_out=16'h8695;
17'h5e21:	data_out=16'h9fa;
17'h5e22:	data_out=16'h89f8;
17'h5e23:	data_out=16'ha00;
17'h5e24:	data_out=16'ha00;
17'h5e25:	data_out=16'h8866;
17'h5e26:	data_out=16'h8812;
17'h5e27:	data_out=16'h87b4;
17'h5e28:	data_out=16'h9f8;
17'h5e29:	data_out=16'h871;
17'h5e2a:	data_out=16'h7c8;
17'h5e2b:	data_out=16'h89fa;
17'h5e2c:	data_out=16'h6af;
17'h5e2d:	data_out=16'h89d9;
17'h5e2e:	data_out=16'h8897;
17'h5e2f:	data_out=16'h893a;
17'h5e30:	data_out=16'h8a00;
17'h5e31:	data_out=16'h9fe;
17'h5e32:	data_out=16'h89fd;
17'h5e33:	data_out=16'h89ff;
17'h5e34:	data_out=16'h89c7;
17'h5e35:	data_out=16'h8960;
17'h5e36:	data_out=16'h88cf;
17'h5e37:	data_out=16'h88be;
17'h5e38:	data_out=16'h8a00;
17'h5e39:	data_out=16'h89fe;
17'h5e3a:	data_out=16'h8738;
17'h5e3b:	data_out=16'h80;
17'h5e3c:	data_out=16'h8526;
17'h5e3d:	data_out=16'h85a2;
17'h5e3e:	data_out=16'h9f8;
17'h5e3f:	data_out=16'h922;
17'h5e40:	data_out=16'h8ca;
17'h5e41:	data_out=16'h8a00;
17'h5e42:	data_out=16'h89b8;
17'h5e43:	data_out=16'h9fe;
17'h5e44:	data_out=16'h9d2;
17'h5e45:	data_out=16'h8c3;
17'h5e46:	data_out=16'h897d;
17'h5e47:	data_out=16'h890b;
17'h5e48:	data_out=16'h89fd;
17'h5e49:	data_out=16'h872a;
17'h5e4a:	data_out=16'h82d1;
17'h5e4b:	data_out=16'h89c1;
17'h5e4c:	data_out=16'h87eb;
17'h5e4d:	data_out=16'h89f8;
17'h5e4e:	data_out=16'h8a00;
17'h5e4f:	data_out=16'h81bc;
17'h5e50:	data_out=16'h89f2;
17'h5e51:	data_out=16'h1b6;
17'h5e52:	data_out=16'h96e;
17'h5e53:	data_out=16'h89b1;
17'h5e54:	data_out=16'h89bf;
17'h5e55:	data_out=16'h3ce;
17'h5e56:	data_out=16'h89aa;
17'h5e57:	data_out=16'h8651;
17'h5e58:	data_out=16'h89ac;
17'h5e59:	data_out=16'h8723;
17'h5e5a:	data_out=16'h89e2;
17'h5e5b:	data_out=16'h895;
17'h5e5c:	data_out=16'h93;
17'h5e5d:	data_out=16'h886c;
17'h5e5e:	data_out=16'h87aa;
17'h5e5f:	data_out=16'h89f4;
17'h5e60:	data_out=16'h87be;
17'h5e61:	data_out=16'h665;
17'h5e62:	data_out=16'h87df;
17'h5e63:	data_out=16'h8a00;
17'h5e64:	data_out=16'h89c2;
17'h5e65:	data_out=16'h89b2;
17'h5e66:	data_out=16'h826b;
17'h5e67:	data_out=16'h369;
17'h5e68:	data_out=16'h9fa;
17'h5e69:	data_out=16'h896f;
17'h5e6a:	data_out=16'h9fd;
17'h5e6b:	data_out=16'h8276;
17'h5e6c:	data_out=16'h4b4;
17'h5e6d:	data_out=16'h8a00;
17'h5e6e:	data_out=16'h9fd;
17'h5e6f:	data_out=16'h971;
17'h5e70:	data_out=16'h9fc;
17'h5e71:	data_out=16'h977;
17'h5e72:	data_out=16'h80dd;
17'h5e73:	data_out=16'h888c;
17'h5e74:	data_out=16'h8a00;
17'h5e75:	data_out=16'h9ad;
17'h5e76:	data_out=16'h89e2;
17'h5e77:	data_out=16'h89ce;
17'h5e78:	data_out=16'h999;
17'h5e79:	data_out=16'h89ff;
17'h5e7a:	data_out=16'h89fd;
17'h5e7b:	data_out=16'h9f8;
17'h5e7c:	data_out=16'h8089;
17'h5e7d:	data_out=16'h89ff;
17'h5e7e:	data_out=16'h32a;
17'h5e7f:	data_out=16'h89ff;
17'h5e80:	data_out=16'h8e3;
17'h5e81:	data_out=16'h9e7;
17'h5e82:	data_out=16'h894d;
17'h5e83:	data_out=16'h89f2;
17'h5e84:	data_out=16'h8ce;
17'h5e85:	data_out=16'h8b5;
17'h5e86:	data_out=16'h8a00;
17'h5e87:	data_out=16'h8195;
17'h5e88:	data_out=16'h891f;
17'h5e89:	data_out=16'h898a;
17'h5e8a:	data_out=16'h9d7;
17'h5e8b:	data_out=16'h88ea;
17'h5e8c:	data_out=16'h8954;
17'h5e8d:	data_out=16'h89bd;
17'h5e8e:	data_out=16'h9fe;
17'h5e8f:	data_out=16'h5a;
17'h5e90:	data_out=16'h89f5;
17'h5e91:	data_out=16'ha00;
17'h5e92:	data_out=16'h1ed;
17'h5e93:	data_out=16'h3fc;
17'h5e94:	data_out=16'h89c8;
17'h5e95:	data_out=16'h9ff;
17'h5e96:	data_out=16'h59f;
17'h5e97:	data_out=16'h89ee;
17'h5e98:	data_out=16'h9fc;
17'h5e99:	data_out=16'h85e;
17'h5e9a:	data_out=16'h7b8;
17'h5e9b:	data_out=16'h8942;
17'h5e9c:	data_out=16'h89d8;
17'h5e9d:	data_out=16'h50a;
17'h5e9e:	data_out=16'h88a2;
17'h5e9f:	data_out=16'h8922;
17'h5ea0:	data_out=16'h8527;
17'h5ea1:	data_out=16'h9fe;
17'h5ea2:	data_out=16'h89fd;
17'h5ea3:	data_out=16'ha00;
17'h5ea4:	data_out=16'ha00;
17'h5ea5:	data_out=16'h88be;
17'h5ea6:	data_out=16'h898c;
17'h5ea7:	data_out=16'h86d5;
17'h5ea8:	data_out=16'h9fc;
17'h5ea9:	data_out=16'h3de;
17'h5eaa:	data_out=16'h9f0;
17'h5eab:	data_out=16'h89ef;
17'h5eac:	data_out=16'h644;
17'h5ead:	data_out=16'h89d0;
17'h5eae:	data_out=16'h85c5;
17'h5eaf:	data_out=16'h88c3;
17'h5eb0:	data_out=16'h8a00;
17'h5eb1:	data_out=16'h9ff;
17'h5eb2:	data_out=16'h89eb;
17'h5eb3:	data_out=16'h89ea;
17'h5eb4:	data_out=16'h36d;
17'h5eb5:	data_out=16'h8991;
17'h5eb6:	data_out=16'h87ee;
17'h5eb7:	data_out=16'h893f;
17'h5eb8:	data_out=16'h8a00;
17'h5eb9:	data_out=16'h89e3;
17'h5eba:	data_out=16'h864a;
17'h5ebb:	data_out=16'h4b;
17'h5ebc:	data_out=16'h89bd;
17'h5ebd:	data_out=16'h9f2;
17'h5ebe:	data_out=16'h9fc;
17'h5ebf:	data_out=16'h89d;
17'h5ec0:	data_out=16'h9cb;
17'h5ec1:	data_out=16'h89f2;
17'h5ec2:	data_out=16'h89cf;
17'h5ec3:	data_out=16'h9e3;
17'h5ec4:	data_out=16'h9ce;
17'h5ec5:	data_out=16'h9ec;
17'h5ec6:	data_out=16'h89c9;
17'h5ec7:	data_out=16'h819e;
17'h5ec8:	data_out=16'h88b9;
17'h5ec9:	data_out=16'h888d;
17'h5eca:	data_out=16'h9e6;
17'h5ecb:	data_out=16'h8994;
17'h5ecc:	data_out=16'h802b;
17'h5ecd:	data_out=16'h89fb;
17'h5ece:	data_out=16'h81ea;
17'h5ecf:	data_out=16'h996;
17'h5ed0:	data_out=16'h89f4;
17'h5ed1:	data_out=16'h85e1;
17'h5ed2:	data_out=16'h9dc;
17'h5ed3:	data_out=16'h8968;
17'h5ed4:	data_out=16'h88d7;
17'h5ed5:	data_out=16'h8808;
17'h5ed6:	data_out=16'h898d;
17'h5ed7:	data_out=16'h82e3;
17'h5ed8:	data_out=16'h899b;
17'h5ed9:	data_out=16'h9d3;
17'h5eda:	data_out=16'h89c6;
17'h5edb:	data_out=16'h9cd;
17'h5edc:	data_out=16'h1fc;
17'h5edd:	data_out=16'h713;
17'h5ede:	data_out=16'h87e0;
17'h5edf:	data_out=16'h9fa;
17'h5ee0:	data_out=16'h27d;
17'h5ee1:	data_out=16'h668;
17'h5ee2:	data_out=16'h894e;
17'h5ee3:	data_out=16'h89eb;
17'h5ee4:	data_out=16'h86c5;
17'h5ee5:	data_out=16'h88ff;
17'h5ee6:	data_out=16'h8635;
17'h5ee7:	data_out=16'h9dd;
17'h5ee8:	data_out=16'h9fe;
17'h5ee9:	data_out=16'h8964;
17'h5eea:	data_out=16'h9fe;
17'h5eeb:	data_out=16'h825;
17'h5eec:	data_out=16'h917;
17'h5eed:	data_out=16'h89ea;
17'h5eee:	data_out=16'h9fe;
17'h5eef:	data_out=16'h97c;
17'h5ef0:	data_out=16'h9fe;
17'h5ef1:	data_out=16'h9f1;
17'h5ef2:	data_out=16'h623;
17'h5ef3:	data_out=16'h646;
17'h5ef4:	data_out=16'h8a00;
17'h5ef5:	data_out=16'h845d;
17'h5ef6:	data_out=16'h8933;
17'h5ef7:	data_out=16'h89c9;
17'h5ef8:	data_out=16'h49c;
17'h5ef9:	data_out=16'h89a2;
17'h5efa:	data_out=16'h89c9;
17'h5efb:	data_out=16'h9fc;
17'h5efc:	data_out=16'h9fc;
17'h5efd:	data_out=16'h87c6;
17'h5efe:	data_out=16'h81d8;
17'h5eff:	data_out=16'h89ff;
17'h5f00:	data_out=16'ha00;
17'h5f01:	data_out=16'h9ff;
17'h5f02:	data_out=16'h298;
17'h5f03:	data_out=16'h89fa;
17'h5f04:	data_out=16'h9ff;
17'h5f05:	data_out=16'h9dc;
17'h5f06:	data_out=16'h8a00;
17'h5f07:	data_out=16'ha00;
17'h5f08:	data_out=16'h855b;
17'h5f09:	data_out=16'h89fb;
17'h5f0a:	data_out=16'h9ff;
17'h5f0b:	data_out=16'h89ec;
17'h5f0c:	data_out=16'h77;
17'h5f0d:	data_out=16'h8951;
17'h5f0e:	data_out=16'ha00;
17'h5f0f:	data_out=16'ha00;
17'h5f10:	data_out=16'h8a00;
17'h5f11:	data_out=16'ha00;
17'h5f12:	data_out=16'h78d;
17'h5f13:	data_out=16'h1ca;
17'h5f14:	data_out=16'h89fb;
17'h5f15:	data_out=16'ha00;
17'h5f16:	data_out=16'h9f5;
17'h5f17:	data_out=16'h89fc;
17'h5f18:	data_out=16'ha00;
17'h5f19:	data_out=16'h89f5;
17'h5f1a:	data_out=16'h9d7;
17'h5f1b:	data_out=16'h89d7;
17'h5f1c:	data_out=16'h89f7;
17'h5f1d:	data_out=16'h859;
17'h5f1e:	data_out=16'h883b;
17'h5f1f:	data_out=16'h6fa;
17'h5f20:	data_out=16'h8803;
17'h5f21:	data_out=16'ha00;
17'h5f22:	data_out=16'h8a00;
17'h5f23:	data_out=16'ha00;
17'h5f24:	data_out=16'ha00;
17'h5f25:	data_out=16'h83c9;
17'h5f26:	data_out=16'h775;
17'h5f27:	data_out=16'h881a;
17'h5f28:	data_out=16'ha00;
17'h5f29:	data_out=16'h867f;
17'h5f2a:	data_out=16'h9ff;
17'h5f2b:	data_out=16'h8a00;
17'h5f2c:	data_out=16'h9f5;
17'h5f2d:	data_out=16'h89e5;
17'h5f2e:	data_out=16'h83d3;
17'h5f2f:	data_out=16'h89a6;
17'h5f30:	data_out=16'h66e;
17'h5f31:	data_out=16'ha00;
17'h5f32:	data_out=16'h98b;
17'h5f33:	data_out=16'h89fe;
17'h5f34:	data_out=16'h8445;
17'h5f35:	data_out=16'h9a9;
17'h5f36:	data_out=16'h886b;
17'h5f37:	data_out=16'h822c;
17'h5f38:	data_out=16'h888a;
17'h5f39:	data_out=16'h89fc;
17'h5f3a:	data_out=16'h9c6;
17'h5f3b:	data_out=16'h8e7;
17'h5f3c:	data_out=16'h8a00;
17'h5f3d:	data_out=16'ha00;
17'h5f3e:	data_out=16'ha00;
17'h5f3f:	data_out=16'h9dd;
17'h5f40:	data_out=16'h9f2;
17'h5f41:	data_out=16'h89fe;
17'h5f42:	data_out=16'h89e2;
17'h5f43:	data_out=16'h696;
17'h5f44:	data_out=16'h95b;
17'h5f45:	data_out=16'ha00;
17'h5f46:	data_out=16'h89ef;
17'h5f47:	data_out=16'h9fd;
17'h5f48:	data_out=16'h886c;
17'h5f49:	data_out=16'h808a;
17'h5f4a:	data_out=16'h5e0;
17'h5f4b:	data_out=16'h89ec;
17'h5f4c:	data_out=16'h9fe;
17'h5f4d:	data_out=16'h89ff;
17'h5f4e:	data_out=16'hb4;
17'h5f4f:	data_out=16'h9e4;
17'h5f50:	data_out=16'h89fa;
17'h5f51:	data_out=16'h328;
17'h5f52:	data_out=16'h9fe;
17'h5f53:	data_out=16'h89e0;
17'h5f54:	data_out=16'h8934;
17'h5f55:	data_out=16'h867d;
17'h5f56:	data_out=16'h992;
17'h5f57:	data_out=16'ha00;
17'h5f58:	data_out=16'h89cf;
17'h5f59:	data_out=16'ha00;
17'h5f5a:	data_out=16'h89ff;
17'h5f5b:	data_out=16'h9f5;
17'h5f5c:	data_out=16'h89f0;
17'h5f5d:	data_out=16'h922;
17'h5f5e:	data_out=16'h891a;
17'h5f5f:	data_out=16'ha00;
17'h5f60:	data_out=16'h9fc;
17'h5f61:	data_out=16'h9f2;
17'h5f62:	data_out=16'h89e5;
17'h5f63:	data_out=16'h89fe;
17'h5f64:	data_out=16'h89fb;
17'h5f65:	data_out=16'h8906;
17'h5f66:	data_out=16'h8981;
17'h5f67:	data_out=16'h803b;
17'h5f68:	data_out=16'ha00;
17'h5f69:	data_out=16'h899d;
17'h5f6a:	data_out=16'ha00;
17'h5f6b:	data_out=16'h9e2;
17'h5f6c:	data_out=16'ha00;
17'h5f6d:	data_out=16'h89fe;
17'h5f6e:	data_out=16'ha00;
17'h5f6f:	data_out=16'h9b5;
17'h5f70:	data_out=16'ha00;
17'h5f71:	data_out=16'ha00;
17'h5f72:	data_out=16'h9f1;
17'h5f73:	data_out=16'h9e1;
17'h5f74:	data_out=16'h7a4;
17'h5f75:	data_out=16'h89b1;
17'h5f76:	data_out=16'h89e4;
17'h5f77:	data_out=16'h89f3;
17'h5f78:	data_out=16'h89ff;
17'h5f79:	data_out=16'h8997;
17'h5f7a:	data_out=16'h89fd;
17'h5f7b:	data_out=16'ha00;
17'h5f7c:	data_out=16'ha00;
17'h5f7d:	data_out=16'h8536;
17'h5f7e:	data_out=16'h84b5;
17'h5f7f:	data_out=16'h5da;
17'h5f80:	data_out=16'h8a8;
17'h5f81:	data_out=16'h8278;
17'h5f82:	data_out=16'h9ff;
17'h5f83:	data_out=16'h89ee;
17'h5f84:	data_out=16'ha00;
17'h5f85:	data_out=16'h9f9;
17'h5f86:	data_out=16'h9ce;
17'h5f87:	data_out=16'ha00;
17'h5f88:	data_out=16'h494;
17'h5f89:	data_out=16'h28b;
17'h5f8a:	data_out=16'ha00;
17'h5f8b:	data_out=16'h89ea;
17'h5f8c:	data_out=16'h662;
17'h5f8d:	data_out=16'h9e8;
17'h5f8e:	data_out=16'ha00;
17'h5f8f:	data_out=16'h9ff;
17'h5f90:	data_out=16'h8a00;
17'h5f91:	data_out=16'h9f6;
17'h5f92:	data_out=16'h9fc;
17'h5f93:	data_out=16'h594;
17'h5f94:	data_out=16'h89f8;
17'h5f95:	data_out=16'ha00;
17'h5f96:	data_out=16'h9ff;
17'h5f97:	data_out=16'h89f8;
17'h5f98:	data_out=16'ha00;
17'h5f99:	data_out=16'h8a00;
17'h5f9a:	data_out=16'h9f7;
17'h5f9b:	data_out=16'h89df;
17'h5f9c:	data_out=16'h85db;
17'h5f9d:	data_out=16'h84d8;
17'h5f9e:	data_out=16'h9e2;
17'h5f9f:	data_out=16'h9fd;
17'h5fa0:	data_out=16'h89f3;
17'h5fa1:	data_out=16'ha00;
17'h5fa2:	data_out=16'h89f6;
17'h5fa3:	data_out=16'ha00;
17'h5fa4:	data_out=16'ha00;
17'h5fa5:	data_out=16'ha00;
17'h5fa6:	data_out=16'h9ff;
17'h5fa7:	data_out=16'h89e6;
17'h5fa8:	data_out=16'ha00;
17'h5fa9:	data_out=16'h123;
17'h5faa:	data_out=16'h9fd;
17'h5fab:	data_out=16'h8a00;
17'h5fac:	data_out=16'h9fd;
17'h5fad:	data_out=16'h89e1;
17'h5fae:	data_out=16'h9fd;
17'h5faf:	data_out=16'h89f9;
17'h5fb0:	data_out=16'h9f6;
17'h5fb1:	data_out=16'h646;
17'h5fb2:	data_out=16'h9ff;
17'h5fb3:	data_out=16'h89ff;
17'h5fb4:	data_out=16'h89d9;
17'h5fb5:	data_out=16'h8f3;
17'h5fb6:	data_out=16'h75c;
17'h5fb7:	data_out=16'h9fe;
17'h5fb8:	data_out=16'h8845;
17'h5fb9:	data_out=16'h89ff;
17'h5fba:	data_out=16'h9de;
17'h5fbb:	data_out=16'h839;
17'h5fbc:	data_out=16'h89f5;
17'h5fbd:	data_out=16'ha00;
17'h5fbe:	data_out=16'ha00;
17'h5fbf:	data_out=16'h9f9;
17'h5fc0:	data_out=16'ha00;
17'h5fc1:	data_out=16'h89f4;
17'h5fc2:	data_out=16'h9c5;
17'h5fc3:	data_out=16'h82c4;
17'h5fc4:	data_out=16'h284;
17'h5fc5:	data_out=16'ha00;
17'h5fc6:	data_out=16'h86e4;
17'h5fc7:	data_out=16'h9e0;
17'h5fc8:	data_out=16'h357;
17'h5fc9:	data_out=16'ha00;
17'h5fca:	data_out=16'h1;
17'h5fcb:	data_out=16'h366;
17'h5fcc:	data_out=16'ha00;
17'h5fcd:	data_out=16'h89fb;
17'h5fce:	data_out=16'h8c2;
17'h5fcf:	data_out=16'ha00;
17'h5fd0:	data_out=16'h89fd;
17'h5fd1:	data_out=16'ha00;
17'h5fd2:	data_out=16'ha00;
17'h5fd3:	data_out=16'h89ed;
17'h5fd4:	data_out=16'h89f1;
17'h5fd5:	data_out=16'ha00;
17'h5fd6:	data_out=16'h9ff;
17'h5fd7:	data_out=16'ha00;
17'h5fd8:	data_out=16'h96b;
17'h5fd9:	data_out=16'ha00;
17'h5fda:	data_out=16'h89f7;
17'h5fdb:	data_out=16'h990;
17'h5fdc:	data_out=16'h89f5;
17'h5fdd:	data_out=16'h9db;
17'h5fde:	data_out=16'h89f0;
17'h5fdf:	data_out=16'h9ff;
17'h5fe0:	data_out=16'h9fe;
17'h5fe1:	data_out=16'ha00;
17'h5fe2:	data_out=16'h89cf;
17'h5fe3:	data_out=16'h8a00;
17'h5fe4:	data_out=16'h8a00;
17'h5fe5:	data_out=16'h89f6;
17'h5fe6:	data_out=16'h89ed;
17'h5fe7:	data_out=16'h89db;
17'h5fe8:	data_out=16'ha00;
17'h5fe9:	data_out=16'h4c6;
17'h5fea:	data_out=16'ha00;
17'h5feb:	data_out=16'h8d8;
17'h5fec:	data_out=16'ha00;
17'h5fed:	data_out=16'h8a00;
17'h5fee:	data_out=16'ha00;
17'h5fef:	data_out=16'h9e6;
17'h5ff0:	data_out=16'ha00;
17'h5ff1:	data_out=16'ha00;
17'h5ff2:	data_out=16'ha00;
17'h5ff3:	data_out=16'ha00;
17'h5ff4:	data_out=16'ha00;
17'h5ff5:	data_out=16'h9ee;
17'h5ff6:	data_out=16'h89eb;
17'h5ff7:	data_out=16'h6ea;
17'h5ff8:	data_out=16'h8a00;
17'h5ff9:	data_out=16'h661;
17'h5ffa:	data_out=16'h89fd;
17'h5ffb:	data_out=16'ha00;
17'h5ffc:	data_out=16'h9ff;
17'h5ffd:	data_out=16'h986;
17'h5ffe:	data_out=16'h837f;
17'h5fff:	data_out=16'h8b1;
17'h6000:	data_out=16'h8cf;
17'h6001:	data_out=16'h7fb;
17'h6002:	data_out=16'ha00;
17'h6003:	data_out=16'h6b2;
17'h6004:	data_out=16'ha00;
17'h6005:	data_out=16'ha00;
17'h6006:	data_out=16'h7b0;
17'h6007:	data_out=16'ha00;
17'h6008:	data_out=16'h9d8;
17'h6009:	data_out=16'h97b;
17'h600a:	data_out=16'ha00;
17'h600b:	data_out=16'h8a00;
17'h600c:	data_out=16'h948;
17'h600d:	data_out=16'ha00;
17'h600e:	data_out=16'ha00;
17'h600f:	data_out=16'ha00;
17'h6010:	data_out=16'h89ff;
17'h6011:	data_out=16'h962;
17'h6012:	data_out=16'ha00;
17'h6013:	data_out=16'ha00;
17'h6014:	data_out=16'h8371;
17'h6015:	data_out=16'ha00;
17'h6016:	data_out=16'ha00;
17'h6017:	data_out=16'h89d9;
17'h6018:	data_out=16'ha00;
17'h6019:	data_out=16'h8a00;
17'h601a:	data_out=16'ha00;
17'h601b:	data_out=16'h873b;
17'h601c:	data_out=16'h97c;
17'h601d:	data_out=16'h677;
17'h601e:	data_out=16'ha00;
17'h601f:	data_out=16'ha00;
17'h6020:	data_out=16'h7b9;
17'h6021:	data_out=16'ha00;
17'h6022:	data_out=16'h8397;
17'h6023:	data_out=16'ha00;
17'h6024:	data_out=16'ha00;
17'h6025:	data_out=16'ha00;
17'h6026:	data_out=16'h9ff;
17'h6027:	data_out=16'h3a9;
17'h6028:	data_out=16'ha00;
17'h6029:	data_out=16'h834a;
17'h602a:	data_out=16'ha00;
17'h602b:	data_out=16'h8a00;
17'h602c:	data_out=16'ha00;
17'h602d:	data_out=16'h89fe;
17'h602e:	data_out=16'ha00;
17'h602f:	data_out=16'h87c9;
17'h6030:	data_out=16'ha00;
17'h6031:	data_out=16'h8828;
17'h6032:	data_out=16'ha00;
17'h6033:	data_out=16'h8214;
17'h6034:	data_out=16'h89f3;
17'h6035:	data_out=16'h9f2;
17'h6036:	data_out=16'h9fd;
17'h6037:	data_out=16'ha00;
17'h6038:	data_out=16'h82a9;
17'h6039:	data_out=16'h1c6;
17'h603a:	data_out=16'h9ee;
17'h603b:	data_out=16'h891;
17'h603c:	data_out=16'h4c9;
17'h603d:	data_out=16'ha00;
17'h603e:	data_out=16'ha00;
17'h603f:	data_out=16'ha00;
17'h6040:	data_out=16'ha00;
17'h6041:	data_out=16'h654;
17'h6042:	data_out=16'ha00;
17'h6043:	data_out=16'h463;
17'h6044:	data_out=16'h52c;
17'h6045:	data_out=16'ha00;
17'h6046:	data_out=16'h86d2;
17'h6047:	data_out=16'h9ed;
17'h6048:	data_out=16'ha00;
17'h6049:	data_out=16'ha00;
17'h604a:	data_out=16'h532;
17'h604b:	data_out=16'ha00;
17'h604c:	data_out=16'ha00;
17'h604d:	data_out=16'h86df;
17'h604e:	data_out=16'h9fa;
17'h604f:	data_out=16'ha00;
17'h6050:	data_out=16'h799;
17'h6051:	data_out=16'ha00;
17'h6052:	data_out=16'ha00;
17'h6053:	data_out=16'h89f4;
17'h6054:	data_out=16'h74b;
17'h6055:	data_out=16'ha00;
17'h6056:	data_out=16'ha00;
17'h6057:	data_out=16'ha00;
17'h6058:	data_out=16'h9ff;
17'h6059:	data_out=16'ha00;
17'h605a:	data_out=16'h89fb;
17'h605b:	data_out=16'h9e2;
17'h605c:	data_out=16'h89ef;
17'h605d:	data_out=16'ha00;
17'h605e:	data_out=16'h87f1;
17'h605f:	data_out=16'ha00;
17'h6060:	data_out=16'h9ff;
17'h6061:	data_out=16'ha00;
17'h6062:	data_out=16'h8962;
17'h6063:	data_out=16'h845d;
17'h6064:	data_out=16'h8a00;
17'h6065:	data_out=16'h8a00;
17'h6066:	data_out=16'h89f3;
17'h6067:	data_out=16'h88cb;
17'h6068:	data_out=16'ha00;
17'h6069:	data_out=16'h9f5;
17'h606a:	data_out=16'ha00;
17'h606b:	data_out=16'ha00;
17'h606c:	data_out=16'ha00;
17'h606d:	data_out=16'h8366;
17'h606e:	data_out=16'ha00;
17'h606f:	data_out=16'ha00;
17'h6070:	data_out=16'ha00;
17'h6071:	data_out=16'ha00;
17'h6072:	data_out=16'ha00;
17'h6073:	data_out=16'ha00;
17'h6074:	data_out=16'ha00;
17'h6075:	data_out=16'ha00;
17'h6076:	data_out=16'h89fd;
17'h6077:	data_out=16'ha00;
17'h6078:	data_out=16'h1e1;
17'h6079:	data_out=16'h9ff;
17'h607a:	data_out=16'h81b2;
17'h607b:	data_out=16'ha00;
17'h607c:	data_out=16'ha00;
17'h607d:	data_out=16'h9ff;
17'h607e:	data_out=16'h847d;
17'h607f:	data_out=16'h9f9;
17'h6080:	data_out=16'h751;
17'h6081:	data_out=16'h935;
17'h6082:	data_out=16'ha00;
17'h6083:	data_out=16'h92d;
17'h6084:	data_out=16'ha00;
17'h6085:	data_out=16'ha00;
17'h6086:	data_out=16'h7c4;
17'h6087:	data_out=16'h9fa;
17'h6088:	data_out=16'h9ff;
17'h6089:	data_out=16'h83a;
17'h608a:	data_out=16'ha00;
17'h608b:	data_out=16'h89ff;
17'h608c:	data_out=16'h9b2;
17'h608d:	data_out=16'h9fc;
17'h608e:	data_out=16'ha00;
17'h608f:	data_out=16'ha00;
17'h6090:	data_out=16'h8a5;
17'h6091:	data_out=16'ha00;
17'h6092:	data_out=16'h344;
17'h6093:	data_out=16'h877;
17'h6094:	data_out=16'h3ae;
17'h6095:	data_out=16'ha00;
17'h6096:	data_out=16'ha00;
17'h6097:	data_out=16'h89ea;
17'h6098:	data_out=16'ha00;
17'h6099:	data_out=16'h8a00;
17'h609a:	data_out=16'ha00;
17'h609b:	data_out=16'h85f0;
17'h609c:	data_out=16'h9e8;
17'h609d:	data_out=16'h7ff;
17'h609e:	data_out=16'ha00;
17'h609f:	data_out=16'h9ff;
17'h60a0:	data_out=16'h9cc;
17'h60a1:	data_out=16'ha00;
17'h60a2:	data_out=16'h82e7;
17'h60a3:	data_out=16'ha00;
17'h60a4:	data_out=16'ha00;
17'h60a5:	data_out=16'ha00;
17'h60a6:	data_out=16'ha00;
17'h60a7:	data_out=16'h8c6;
17'h60a8:	data_out=16'ha00;
17'h60a9:	data_out=16'h883e;
17'h60aa:	data_out=16'ha00;
17'h60ab:	data_out=16'h8a00;
17'h60ac:	data_out=16'ha00;
17'h60ad:	data_out=16'h89ff;
17'h60ae:	data_out=16'ha00;
17'h60af:	data_out=16'h4ef;
17'h60b0:	data_out=16'ha00;
17'h60b1:	data_out=16'h89fe;
17'h60b2:	data_out=16'ha00;
17'h60b3:	data_out=16'h5a4;
17'h60b4:	data_out=16'h820d;
17'h60b5:	data_out=16'h9fb;
17'h60b6:	data_out=16'h9ff;
17'h60b7:	data_out=16'ha00;
17'h60b8:	data_out=16'h59a;
17'h60b9:	data_out=16'h7d5;
17'h60ba:	data_out=16'h359;
17'h60bb:	data_out=16'h97f;
17'h60bc:	data_out=16'h9f7;
17'h60bd:	data_out=16'ha00;
17'h60be:	data_out=16'ha00;
17'h60bf:	data_out=16'ha00;
17'h60c0:	data_out=16'ha00;
17'h60c1:	data_out=16'h9e3;
17'h60c2:	data_out=16'ha00;
17'h60c3:	data_out=16'h20a;
17'h60c4:	data_out=16'h70d;
17'h60c5:	data_out=16'ha00;
17'h60c6:	data_out=16'h8466;
17'h60c7:	data_out=16'h9f9;
17'h60c8:	data_out=16'h9bd;
17'h60c9:	data_out=16'ha00;
17'h60ca:	data_out=16'h919;
17'h60cb:	data_out=16'h75d;
17'h60cc:	data_out=16'ha00;
17'h60cd:	data_out=16'h8434;
17'h60ce:	data_out=16'ha00;
17'h60cf:	data_out=16'ha00;
17'h60d0:	data_out=16'h98c;
17'h60d1:	data_out=16'ha00;
17'h60d2:	data_out=16'ha00;
17'h60d3:	data_out=16'h87e8;
17'h60d4:	data_out=16'h9f6;
17'h60d5:	data_out=16'ha00;
17'h60d6:	data_out=16'ha00;
17'h60d7:	data_out=16'ha00;
17'h60d8:	data_out=16'ha00;
17'h60d9:	data_out=16'ha00;
17'h60da:	data_out=16'h89fd;
17'h60db:	data_out=16'ha00;
17'h60dc:	data_out=16'h1fa;
17'h60dd:	data_out=16'ha00;
17'h60de:	data_out=16'h4a8;
17'h60df:	data_out=16'ha00;
17'h60e0:	data_out=16'ha00;
17'h60e1:	data_out=16'ha00;
17'h60e2:	data_out=16'h8974;
17'h60e3:	data_out=16'h50e;
17'h60e4:	data_out=16'h8a00;
17'h60e5:	data_out=16'h88be;
17'h60e6:	data_out=16'h8a00;
17'h60e7:	data_out=16'h85df;
17'h60e8:	data_out=16'ha00;
17'h60e9:	data_out=16'h9f9;
17'h60ea:	data_out=16'ha00;
17'h60eb:	data_out=16'ha00;
17'h60ec:	data_out=16'h9a5;
17'h60ed:	data_out=16'h566;
17'h60ee:	data_out=16'ha00;
17'h60ef:	data_out=16'ha00;
17'h60f0:	data_out=16'ha00;
17'h60f1:	data_out=16'ha00;
17'h60f2:	data_out=16'ha00;
17'h60f3:	data_out=16'ha00;
17'h60f4:	data_out=16'ha00;
17'h60f5:	data_out=16'ha00;
17'h60f6:	data_out=16'h8a00;
17'h60f7:	data_out=16'ha00;
17'h60f8:	data_out=16'h44f;
17'h60f9:	data_out=16'ha00;
17'h60fa:	data_out=16'h5fb;
17'h60fb:	data_out=16'ha00;
17'h60fc:	data_out=16'ha00;
17'h60fd:	data_out=16'h9fd;
17'h60fe:	data_out=16'he;
17'h60ff:	data_out=16'ha00;
17'h6100:	data_out=16'h3e7;
17'h6101:	data_out=16'h5c3;
17'h6102:	data_out=16'ha00;
17'h6103:	data_out=16'h5b9;
17'h6104:	data_out=16'ha00;
17'h6105:	data_out=16'ha00;
17'h6106:	data_out=16'h385;
17'h6107:	data_out=16'h652;
17'h6108:	data_out=16'ha00;
17'h6109:	data_out=16'h811b;
17'h610a:	data_out=16'h6bf;
17'h610b:	data_out=16'h8a00;
17'h610c:	data_out=16'h99b;
17'h610d:	data_out=16'h798;
17'h610e:	data_out=16'h5ae;
17'h610f:	data_out=16'ha00;
17'h6110:	data_out=16'h1e2;
17'h6111:	data_out=16'h9db;
17'h6112:	data_out=16'h9;
17'h6113:	data_out=16'h4df;
17'h6114:	data_out=16'h31a;
17'h6115:	data_out=16'ha00;
17'h6116:	data_out=16'ha00;
17'h6117:	data_out=16'h8207;
17'h6118:	data_out=16'h964;
17'h6119:	data_out=16'h8a00;
17'h611a:	data_out=16'ha00;
17'h611b:	data_out=16'h8473;
17'h611c:	data_out=16'ha00;
17'h611d:	data_out=16'h557;
17'h611e:	data_out=16'h5e1;
17'h611f:	data_out=16'h9f7;
17'h6120:	data_out=16'h99e;
17'h6121:	data_out=16'h59b;
17'h6122:	data_out=16'h849c;
17'h6123:	data_out=16'h7e1;
17'h6124:	data_out=16'h7e9;
17'h6125:	data_out=16'h227;
17'h6126:	data_out=16'h810e;
17'h6127:	data_out=16'h559;
17'h6128:	data_out=16'h583;
17'h6129:	data_out=16'h8292;
17'h612a:	data_out=16'h66b;
17'h612b:	data_out=16'h8a00;
17'h612c:	data_out=16'ha00;
17'h612d:	data_out=16'h8a00;
17'h612e:	data_out=16'h9f9;
17'h612f:	data_out=16'h3b6;
17'h6130:	data_out=16'ha00;
17'h6131:	data_out=16'h85a1;
17'h6132:	data_out=16'ha00;
17'h6133:	data_out=16'h440;
17'h6134:	data_out=16'h81e1;
17'h6135:	data_out=16'ha00;
17'h6136:	data_out=16'ha00;
17'h6137:	data_out=16'ha00;
17'h6138:	data_out=16'h8ad;
17'h6139:	data_out=16'h54c;
17'h613a:	data_out=16'h8078;
17'h613b:	data_out=16'h993;
17'h613c:	data_out=16'h7e4;
17'h613d:	data_out=16'ha00;
17'h613e:	data_out=16'h584;
17'h613f:	data_out=16'ha00;
17'h6140:	data_out=16'ha00;
17'h6141:	data_out=16'ha00;
17'h6142:	data_out=16'h140;
17'h6143:	data_out=16'h1e0;
17'h6144:	data_out=16'h9aa;
17'h6145:	data_out=16'ha00;
17'h6146:	data_out=16'h8715;
17'h6147:	data_out=16'h21b;
17'h6148:	data_out=16'h35;
17'h6149:	data_out=16'h2d8;
17'h614a:	data_out=16'h9ef;
17'h614b:	data_out=16'h8264;
17'h614c:	data_out=16'h716;
17'h614d:	data_out=16'h84bc;
17'h614e:	data_out=16'ha00;
17'h614f:	data_out=16'h6f2;
17'h6150:	data_out=16'h9fd;
17'h6151:	data_out=16'ha00;
17'h6152:	data_out=16'h87c;
17'h6153:	data_out=16'h80ea;
17'h6154:	data_out=16'h9b8;
17'h6155:	data_out=16'h9ff;
17'h6156:	data_out=16'ha00;
17'h6157:	data_out=16'ha00;
17'h6158:	data_out=16'ha00;
17'h6159:	data_out=16'ha00;
17'h615a:	data_out=16'h850a;
17'h615b:	data_out=16'ha00;
17'h615c:	data_out=16'h4f0;
17'h615d:	data_out=16'ha00;
17'h615e:	data_out=16'h2d8;
17'h615f:	data_out=16'h53e;
17'h6160:	data_out=16'h824b;
17'h6161:	data_out=16'ha00;
17'h6162:	data_out=16'h831b;
17'h6163:	data_out=16'h3f5;
17'h6164:	data_out=16'h85fb;
17'h6165:	data_out=16'h863f;
17'h6166:	data_out=16'h8a00;
17'h6167:	data_out=16'h83df;
17'h6168:	data_out=16'h58e;
17'h6169:	data_out=16'ha00;
17'h616a:	data_out=16'h5be;
17'h616b:	data_out=16'ha00;
17'h616c:	data_out=16'h7f4;
17'h616d:	data_out=16'h40f;
17'h616e:	data_out=16'h5be;
17'h616f:	data_out=16'h77f;
17'h6170:	data_out=16'h5b6;
17'h6171:	data_out=16'ha00;
17'h6172:	data_out=16'ha00;
17'h6173:	data_out=16'ha00;
17'h6174:	data_out=16'ha00;
17'h6175:	data_out=16'h997;
17'h6176:	data_out=16'h8a00;
17'h6177:	data_out=16'ha00;
17'h6178:	data_out=16'haa;
17'h6179:	data_out=16'ha00;
17'h617a:	data_out=16'h3f4;
17'h617b:	data_out=16'h584;
17'h617c:	data_out=16'h762;
17'h617d:	data_out=16'h4df;
17'h617e:	data_out=16'h83ca;
17'h617f:	data_out=16'ha00;
17'h6180:	data_out=16'h8348;
17'h6181:	data_out=16'h8161;
17'h6182:	data_out=16'h8125;
17'h6183:	data_out=16'h80bb;
17'h6184:	data_out=16'h34a;
17'h6185:	data_out=16'h109;
17'h6186:	data_out=16'h12e;
17'h6187:	data_out=16'h8a;
17'h6188:	data_out=16'h839a;
17'h6189:	data_out=16'h81e6;
17'h618a:	data_out=16'h80ec;
17'h618b:	data_out=16'h834b;
17'h618c:	data_out=16'h32c;
17'h618d:	data_out=16'h8062;
17'h618e:	data_out=16'h6d;
17'h618f:	data_out=16'h80fc;
17'h6190:	data_out=16'h8117;
17'h6191:	data_out=16'h10c;
17'h6192:	data_out=16'h8232;
17'h6193:	data_out=16'h9c;
17'h6194:	data_out=16'h81b9;
17'h6195:	data_out=16'h8017;
17'h6196:	data_out=16'h80c5;
17'h6197:	data_out=16'h81d9;
17'h6198:	data_out=16'h8012;
17'h6199:	data_out=16'h22c;
17'h619a:	data_out=16'h2e9;
17'h619b:	data_out=16'h825d;
17'h619c:	data_out=16'h80da;
17'h619d:	data_out=16'h832e;
17'h619e:	data_out=16'h826c;
17'h619f:	data_out=16'h2a;
17'h61a0:	data_out=16'h82bb;
17'h61a1:	data_out=16'h5d;
17'h61a2:	data_out=16'h800f;
17'h61a3:	data_out=16'hf1;
17'h61a4:	data_out=16'hf1;
17'h61a5:	data_out=16'h165;
17'h61a6:	data_out=16'h84b1;
17'h61a7:	data_out=16'h8415;
17'h61a8:	data_out=16'h68;
17'h61a9:	data_out=16'h8096;
17'h61aa:	data_out=16'h830e;
17'h61ab:	data_out=16'h84ee;
17'h61ac:	data_out=16'h80eb;
17'h61ad:	data_out=16'h800b;
17'h61ae:	data_out=16'h8263;
17'h61af:	data_out=16'h8185;
17'h61b0:	data_out=16'h292;
17'h61b1:	data_out=16'h81fa;
17'h61b2:	data_out=16'h28e;
17'h61b3:	data_out=16'h826d;
17'h61b4:	data_out=16'h80f5;
17'h61b5:	data_out=16'h1b8;
17'h61b6:	data_out=16'h828b;
17'h61b7:	data_out=16'h811f;
17'h61b8:	data_out=16'h252;
17'h61b9:	data_out=16'h8249;
17'h61ba:	data_out=16'h8185;
17'h61bb:	data_out=16'h80eb;
17'h61bc:	data_out=16'h821f;
17'h61bd:	data_out=16'h8212;
17'h61be:	data_out=16'h63;
17'h61bf:	data_out=16'h223;
17'h61c0:	data_out=16'h301;
17'h61c1:	data_out=16'h820f;
17'h61c2:	data_out=16'h338;
17'h61c3:	data_out=16'h1f0;
17'h61c4:	data_out=16'h812d;
17'h61c5:	data_out=16'h8080;
17'h61c6:	data_out=16'h8228;
17'h61c7:	data_out=16'h8106;
17'h61c8:	data_out=16'h8148;
17'h61c9:	data_out=16'h169;
17'h61ca:	data_out=16'h237;
17'h61cb:	data_out=16'h2e1;
17'h61cc:	data_out=16'h2a9;
17'h61cd:	data_out=16'ha;
17'h61ce:	data_out=16'h810c;
17'h61cf:	data_out=16'h201;
17'h61d0:	data_out=16'h29c;
17'h61d1:	data_out=16'h80fc;
17'h61d2:	data_out=16'h103;
17'h61d3:	data_out=16'h83c9;
17'h61d4:	data_out=16'h81d2;
17'h61d5:	data_out=16'h81d6;
17'h61d6:	data_out=16'h80f4;
17'h61d7:	data_out=16'h6;
17'h61d8:	data_out=16'h81ed;
17'h61d9:	data_out=16'h217;
17'h61da:	data_out=16'h82a8;
17'h61db:	data_out=16'h8033;
17'h61dc:	data_out=16'h8173;
17'h61dd:	data_out=16'h80e2;
17'h61de:	data_out=16'h8108;
17'h61df:	data_out=16'h8054;
17'h61e0:	data_out=16'h827f;
17'h61e1:	data_out=16'h1f;
17'h61e2:	data_out=16'h8285;
17'h61e3:	data_out=16'h822a;
17'h61e4:	data_out=16'h821c;
17'h61e5:	data_out=16'h1e0;
17'h61e6:	data_out=16'h1af;
17'h61e7:	data_out=16'h81b7;
17'h61e8:	data_out=16'h5c;
17'h61e9:	data_out=16'h8304;
17'h61ea:	data_out=16'h71;
17'h61eb:	data_out=16'h1f6;
17'h61ec:	data_out=16'h81b4;
17'h61ed:	data_out=16'h8260;
17'h61ee:	data_out=16'h6a;
17'h61ef:	data_out=16'h131;
17'h61f0:	data_out=16'h6c;
17'h61f1:	data_out=16'h8298;
17'h61f2:	data_out=16'h1ee;
17'h61f3:	data_out=16'h1a2;
17'h61f4:	data_out=16'h277;
17'h61f5:	data_out=16'hea;
17'h61f6:	data_out=16'h84fd;
17'h61f7:	data_out=16'h2e7;
17'h61f8:	data_out=16'h1e6;
17'h61f9:	data_out=16'h82cb;
17'h61fa:	data_out=16'h81f6;
17'h61fb:	data_out=16'h5a;
17'h61fc:	data_out=16'h8097;
17'h61fd:	data_out=16'h122;
17'h61fe:	data_out=16'h81fa;
17'h61ff:	data_out=16'h291;
17'h6200:	data_out=16'h10;
17'h6201:	data_out=16'he;
17'h6202:	data_out=16'ha;
17'h6203:	data_out=16'h5;
17'h6204:	data_out=16'hd;
17'h6205:	data_out=16'h0;
17'h6206:	data_out=16'h8003;
17'h6207:	data_out=16'he;
17'h6208:	data_out=16'h8001;
17'h6209:	data_out=16'h8003;
17'h620a:	data_out=16'hb;
17'h620b:	data_out=16'h8003;
17'h620c:	data_out=16'hf;
17'h620d:	data_out=16'h3;
17'h620e:	data_out=16'h8002;
17'h620f:	data_out=16'hb;
17'h6210:	data_out=16'h1;
17'h6211:	data_out=16'hc;
17'h6212:	data_out=16'h1;
17'h6213:	data_out=16'h3;
17'h6214:	data_out=16'h1;
17'h6215:	data_out=16'hf;
17'h6216:	data_out=16'hf;
17'h6217:	data_out=16'h8004;
17'h6218:	data_out=16'hd;
17'h6219:	data_out=16'h8001;
17'h621a:	data_out=16'h4;
17'h621b:	data_out=16'hb;
17'h621c:	data_out=16'h8;
17'h621d:	data_out=16'h3;
17'h621e:	data_out=16'h8001;
17'h621f:	data_out=16'h8;
17'h6220:	data_out=16'h2;
17'h6221:	data_out=16'h8006;
17'h6222:	data_out=16'h8005;
17'h6223:	data_out=16'h8002;
17'h6224:	data_out=16'h1;
17'h6225:	data_out=16'h1;
17'h6226:	data_out=16'hc;
17'h6227:	data_out=16'h0;
17'h6228:	data_out=16'h8002;
17'h6229:	data_out=16'h8;
17'h622a:	data_out=16'h5;
17'h622b:	data_out=16'h8004;
17'h622c:	data_out=16'hd;
17'h622d:	data_out=16'h9;
17'h622e:	data_out=16'hb;
17'h622f:	data_out=16'h8004;
17'h6230:	data_out=16'h7;
17'h6231:	data_out=16'h8001;
17'h6232:	data_out=16'h6;
17'h6233:	data_out=16'h6;
17'h6234:	data_out=16'h8001;
17'h6235:	data_out=16'h2;
17'h6236:	data_out=16'h9;
17'h6237:	data_out=16'hf;
17'h6238:	data_out=16'h8000;
17'h6239:	data_out=16'hb;
17'h623a:	data_out=16'hc;
17'h623b:	data_out=16'hf;
17'h623c:	data_out=16'h1;
17'h623d:	data_out=16'h8003;
17'h623e:	data_out=16'h4;
17'h623f:	data_out=16'h8;
17'h6240:	data_out=16'h0;
17'h6241:	data_out=16'h5;
17'h6242:	data_out=16'hc;
17'h6243:	data_out=16'h8001;
17'h6244:	data_out=16'hc;
17'h6245:	data_out=16'h4;
17'h6246:	data_out=16'h3;
17'h6247:	data_out=16'hf;
17'h6248:	data_out=16'hb;
17'h6249:	data_out=16'hc;
17'h624a:	data_out=16'h1;
17'h624b:	data_out=16'h10;
17'h624c:	data_out=16'h8;
17'h624d:	data_out=16'hb;
17'h624e:	data_out=16'he;
17'h624f:	data_out=16'hd;
17'h6250:	data_out=16'hf;
17'h6251:	data_out=16'h10;
17'h6252:	data_out=16'h1;
17'h6253:	data_out=16'hc;
17'h6254:	data_out=16'h8001;
17'h6255:	data_out=16'hd;
17'h6256:	data_out=16'hf;
17'h6257:	data_out=16'h2;
17'h6258:	data_out=16'hc;
17'h6259:	data_out=16'hb;
17'h625a:	data_out=16'h8003;
17'h625b:	data_out=16'he;
17'h625c:	data_out=16'h9;
17'h625d:	data_out=16'hc;
17'h625e:	data_out=16'h6;
17'h625f:	data_out=16'hb;
17'h6260:	data_out=16'h7;
17'h6261:	data_out=16'h8000;
17'h6262:	data_out=16'h8005;
17'h6263:	data_out=16'h8003;
17'h6264:	data_out=16'h7;
17'h6265:	data_out=16'h8;
17'h6266:	data_out=16'h8003;
17'h6267:	data_out=16'h3;
17'h6268:	data_out=16'h8000;
17'h6269:	data_out=16'h0;
17'h626a:	data_out=16'h8004;
17'h626b:	data_out=16'hb;
17'h626c:	data_out=16'hf;
17'h626d:	data_out=16'hc;
17'h626e:	data_out=16'h8001;
17'h626f:	data_out=16'he;
17'h6270:	data_out=16'ha;
17'h6271:	data_out=16'h5;
17'h6272:	data_out=16'hc;
17'h6273:	data_out=16'h12;
17'h6274:	data_out=16'ha;
17'h6275:	data_out=16'ha;
17'h6276:	data_out=16'h2;
17'h6277:	data_out=16'h6;
17'h6278:	data_out=16'h5;
17'h6279:	data_out=16'h7;
17'h627a:	data_out=16'h8001;
17'h627b:	data_out=16'h8003;
17'h627c:	data_out=16'h8000;
17'h627d:	data_out=16'h8;
17'h627e:	data_out=16'hf;
17'h627f:	data_out=16'hc;
17'h6280:	data_out=16'ha0;
17'h6281:	data_out=16'h64;
17'h6282:	data_out=16'h8004;
17'h6283:	data_out=16'h8013;
17'h6284:	data_out=16'h8083;
17'h6285:	data_out=16'hc4;
17'h6286:	data_out=16'hc5;
17'h6287:	data_out=16'h800a;
17'h6288:	data_out=16'h14b;
17'h6289:	data_out=16'h67;
17'h628a:	data_out=16'h8027;
17'h628b:	data_out=16'hde;
17'h628c:	data_out=16'h59;
17'h628d:	data_out=16'h8073;
17'h628e:	data_out=16'h8015;
17'h628f:	data_out=16'h4e;
17'h6290:	data_out=16'h80a4;
17'h6291:	data_out=16'h8020;
17'h6292:	data_out=16'h7c;
17'h6293:	data_out=16'h808e;
17'h6294:	data_out=16'h11;
17'h6295:	data_out=16'h8087;
17'h6296:	data_out=16'h8092;
17'h6297:	data_out=16'h1c;
17'h6298:	data_out=16'h8064;
17'h6299:	data_out=16'h3e;
17'h629a:	data_out=16'h809d;
17'h629b:	data_out=16'h7c;
17'h629c:	data_out=16'h10b;
17'h629d:	data_out=16'h8b;
17'h629e:	data_out=16'hec;
17'h629f:	data_out=16'h52;
17'h62a0:	data_out=16'h16f;
17'h62a1:	data_out=16'h8019;
17'h62a2:	data_out=16'h49;
17'h62a3:	data_out=16'h810f;
17'h62a4:	data_out=16'h8105;
17'h62a5:	data_out=16'h7;
17'h62a6:	data_out=16'h8a;
17'h62a7:	data_out=16'heb;
17'h62a8:	data_out=16'h8010;
17'h62a9:	data_out=16'h8097;
17'h62aa:	data_out=16'h37;
17'h62ab:	data_out=16'hdd;
17'h62ac:	data_out=16'h8021;
17'h62ad:	data_out=16'h80bc;
17'h62ae:	data_out=16'h803d;
17'h62af:	data_out=16'h105;
17'h62b0:	data_out=16'h806c;
17'h62b1:	data_out=16'h6e;
17'h62b2:	data_out=16'h8068;
17'h62b3:	data_out=16'h51;
17'h62b4:	data_out=16'h800c;
17'h62b5:	data_out=16'h89;
17'h62b6:	data_out=16'h16f;
17'h62b7:	data_out=16'h14;
17'h62b8:	data_out=16'hff;
17'h62b9:	data_out=16'h6f;
17'h62ba:	data_out=16'h8075;
17'h62bb:	data_out=16'h4b;
17'h62bc:	data_out=16'h73;
17'h62bd:	data_out=16'h2a;
17'h62be:	data_out=16'h8009;
17'h62bf:	data_out=16'h21;
17'h62c0:	data_out=16'h80d8;
17'h62c1:	data_out=16'h137;
17'h62c2:	data_out=16'hc;
17'h62c3:	data_out=16'h84;
17'h62c4:	data_out=16'h80a8;
17'h62c5:	data_out=16'h8103;
17'h62c6:	data_out=16'h103;
17'h62c7:	data_out=16'h806c;
17'h62c8:	data_out=16'h806b;
17'h62c9:	data_out=16'h8024;
17'h62ca:	data_out=16'h8089;
17'h62cb:	data_out=16'h58;
17'h62cc:	data_out=16'h8084;
17'h62cd:	data_out=16'h83;
17'h62ce:	data_out=16'h15;
17'h62cf:	data_out=16'h808b;
17'h62d0:	data_out=16'h80e9;
17'h62d1:	data_out=16'hc;
17'h62d2:	data_out=16'h80f5;
17'h62d3:	data_out=16'h1b0;
17'h62d4:	data_out=16'h166;
17'h62d5:	data_out=16'he3;
17'h62d6:	data_out=16'h8082;
17'h62d7:	data_out=16'h809e;
17'h62d8:	data_out=16'h8001;
17'h62d9:	data_out=16'h8094;
17'h62da:	data_out=16'h8004;
17'h62db:	data_out=16'h13f;
17'h62dc:	data_out=16'h8f;
17'h62dd:	data_out=16'h805c;
17'h62de:	data_out=16'h10c;
17'h62df:	data_out=16'h8022;
17'h62e0:	data_out=16'h8074;
17'h62e1:	data_out=16'h8003;
17'h62e2:	data_out=16'h146;
17'h62e3:	data_out=16'h48;
17'h62e4:	data_out=16'h8;
17'h62e5:	data_out=16'h804d;
17'h62e6:	data_out=16'hf;
17'h62e7:	data_out=16'h8050;
17'h62e8:	data_out=16'h800e;
17'h62e9:	data_out=16'hac;
17'h62ea:	data_out=16'h801c;
17'h62eb:	data_out=16'h800a;
17'h62ec:	data_out=16'h80a1;
17'h62ed:	data_out=16'h62;
17'h62ee:	data_out=16'h8014;
17'h62ef:	data_out=16'h5a;
17'h62f0:	data_out=16'h801f;
17'h62f1:	data_out=16'h805d;
17'h62f2:	data_out=16'h80fa;
17'h62f3:	data_out=16'h8012;
17'h62f4:	data_out=16'h8067;
17'h62f5:	data_out=16'h92;
17'h62f6:	data_out=16'hd3;
17'h62f7:	data_out=16'h80ff;
17'h62f8:	data_out=16'h8c;
17'h62f9:	data_out=16'h8006;
17'h62fa:	data_out=16'h1a;
17'h62fb:	data_out=16'h8013;
17'h62fc:	data_out=16'h64;
17'h62fd:	data_out=16'h10d;
17'h62fe:	data_out=16'h6f;
17'h62ff:	data_out=16'h8139;
17'h6300:	data_out=16'h5a3;
17'h6301:	data_out=16'h2e1;
17'h6302:	data_out=16'h80d0;
17'h6303:	data_out=16'h29d;
17'h6304:	data_out=16'h81c3;
17'h6305:	data_out=16'h8158;
17'h6306:	data_out=16'h83a2;
17'h6307:	data_out=16'h8051;
17'h6308:	data_out=16'h802a;
17'h6309:	data_out=16'h3a3;
17'h630a:	data_out=16'h1c7;
17'h630b:	data_out=16'h81bf;
17'h630c:	data_out=16'h8616;
17'h630d:	data_out=16'h80b4;
17'h630e:	data_out=16'h8136;
17'h630f:	data_out=16'h808b;
17'h6310:	data_out=16'h3c7;
17'h6311:	data_out=16'h8144;
17'h6312:	data_out=16'h224;
17'h6313:	data_out=16'hc;
17'h6314:	data_out=16'h193;
17'h6315:	data_out=16'h15;
17'h6316:	data_out=16'h803e;
17'h6317:	data_out=16'hd6;
17'h6318:	data_out=16'h80c4;
17'h6319:	data_out=16'h28d;
17'h631a:	data_out=16'h828c;
17'h631b:	data_out=16'h1e7;
17'h631c:	data_out=16'h80a4;
17'h631d:	data_out=16'h429;
17'h631e:	data_out=16'h2cf;
17'h631f:	data_out=16'h82b6;
17'h6320:	data_out=16'ha00;
17'h6321:	data_out=16'h8135;
17'h6322:	data_out=16'h796;
17'h6323:	data_out=16'h8508;
17'h6324:	data_out=16'h8507;
17'h6325:	data_out=16'h2f9;
17'h6326:	data_out=16'h8233;
17'h6327:	data_out=16'h546;
17'h6328:	data_out=16'h811d;
17'h6329:	data_out=16'h2bc;
17'h632a:	data_out=16'hf5;
17'h632b:	data_out=16'h62d;
17'h632c:	data_out=16'h802b;
17'h632d:	data_out=16'h18a;
17'h632e:	data_out=16'h96;
17'h632f:	data_out=16'h710;
17'h6330:	data_out=16'h8647;
17'h6331:	data_out=16'h35d;
17'h6332:	data_out=16'h85d5;
17'h6333:	data_out=16'h2f3;
17'h6334:	data_out=16'hbc;
17'h6335:	data_out=16'h854d;
17'h6336:	data_out=16'h1a7;
17'h6337:	data_out=16'h80e4;
17'h6338:	data_out=16'h8015;
17'h6339:	data_out=16'h366;
17'h633a:	data_out=16'h74d;
17'h633b:	data_out=16'h82f4;
17'h633c:	data_out=16'h8067;
17'h633d:	data_out=16'h4d7;
17'h633e:	data_out=16'h811f;
17'h633f:	data_out=16'h82b3;
17'h6340:	data_out=16'h30;
17'h6341:	data_out=16'h815b;
17'h6342:	data_out=16'h2c3;
17'h6343:	data_out=16'h8401;
17'h6344:	data_out=16'h81a7;
17'h6345:	data_out=16'h810f;
17'h6346:	data_out=16'h18e;
17'h6347:	data_out=16'h306;
17'h6348:	data_out=16'h287;
17'h6349:	data_out=16'h318;
17'h634a:	data_out=16'h8147;
17'h634b:	data_out=16'hd7;
17'h634c:	data_out=16'h133;
17'h634d:	data_out=16'h817;
17'h634e:	data_out=16'h80b1;
17'h634f:	data_out=16'h15f;
17'h6350:	data_out=16'h803b;
17'h6351:	data_out=16'h8731;
17'h6352:	data_out=16'h84e5;
17'h6353:	data_out=16'h761;
17'h6354:	data_out=16'h79b;
17'h6355:	data_out=16'h859c;
17'h6356:	data_out=16'h155;
17'h6357:	data_out=16'h20b;
17'h6358:	data_out=16'h83f4;
17'h6359:	data_out=16'h141;
17'h635a:	data_out=16'h104;
17'h635b:	data_out=16'h8530;
17'h635c:	data_out=16'h226;
17'h635d:	data_out=16'h379;
17'h635e:	data_out=16'h64c;
17'h635f:	data_out=16'h2d6;
17'h6360:	data_out=16'h8389;
17'h6361:	data_out=16'h83e2;
17'h6362:	data_out=16'h82a0;
17'h6363:	data_out=16'h2b2;
17'h6364:	data_out=16'h171;
17'h6365:	data_out=16'h1ee;
17'h6366:	data_out=16'h260;
17'h6367:	data_out=16'h275;
17'h6368:	data_out=16'h8122;
17'h6369:	data_out=16'h81b5;
17'h636a:	data_out=16'h814a;
17'h636b:	data_out=16'h8008;
17'h636c:	data_out=16'h833;
17'h636d:	data_out=16'h2dd;
17'h636e:	data_out=16'h8152;
17'h636f:	data_out=16'h2a;
17'h6370:	data_out=16'h813e;
17'h6371:	data_out=16'h830c;
17'h6372:	data_out=16'h831b;
17'h6373:	data_out=16'h8186;
17'h6374:	data_out=16'h866d;
17'h6375:	data_out=16'h8861;
17'h6376:	data_out=16'h36f;
17'h6377:	data_out=16'h8207;
17'h6378:	data_out=16'h8377;
17'h6379:	data_out=16'h80e8;
17'h637a:	data_out=16'h20a;
17'h637b:	data_out=16'h8113;
17'h637c:	data_out=16'h18;
17'h637d:	data_out=16'h847e;
17'h637e:	data_out=16'h241;
17'h637f:	data_out=16'h8105;
17'h6380:	data_out=16'h83b3;
17'h6381:	data_out=16'ha00;
17'h6382:	data_out=16'h3f8;
17'h6383:	data_out=16'h432;
17'h6384:	data_out=16'h8858;
17'h6385:	data_out=16'h8055;
17'h6386:	data_out=16'h8161;
17'h6387:	data_out=16'h274;
17'h6388:	data_out=16'h97;
17'h6389:	data_out=16'h822e;
17'h638a:	data_out=16'h82d1;
17'h638b:	data_out=16'ha00;
17'h638c:	data_out=16'h8978;
17'h638d:	data_out=16'h596;
17'h638e:	data_out=16'h8296;
17'h638f:	data_out=16'h719;
17'h6390:	data_out=16'h63d;
17'h6391:	data_out=16'h851c;
17'h6392:	data_out=16'ha00;
17'h6393:	data_out=16'h123;
17'h6394:	data_out=16'h9fe;
17'h6395:	data_out=16'h865b;
17'h6396:	data_out=16'h87c8;
17'h6397:	data_out=16'h9fc;
17'h6398:	data_out=16'h815a;
17'h6399:	data_out=16'h1d6;
17'h639a:	data_out=16'h87cb;
17'h639b:	data_out=16'h9fd;
17'h639c:	data_out=16'h8183;
17'h639d:	data_out=16'ha00;
17'h639e:	data_out=16'h9fc;
17'h639f:	data_out=16'h8663;
17'h63a0:	data_out=16'ha00;
17'h63a1:	data_out=16'h8262;
17'h63a2:	data_out=16'h88f;
17'h63a3:	data_out=16'h8a00;
17'h63a4:	data_out=16'h8a00;
17'h63a5:	data_out=16'h261;
17'h63a6:	data_out=16'h8a00;
17'h63a7:	data_out=16'ha00;
17'h63a8:	data_out=16'h81c3;
17'h63a9:	data_out=16'h9d6;
17'h63aa:	data_out=16'h5a4;
17'h63ab:	data_out=16'ha00;
17'h63ac:	data_out=16'h878a;
17'h63ad:	data_out=16'hbd;
17'h63ae:	data_out=16'h9f2;
17'h63af:	data_out=16'ha00;
17'h63b0:	data_out=16'h8a00;
17'h63b1:	data_out=16'h8ec;
17'h63b2:	data_out=16'h89ff;
17'h63b3:	data_out=16'ha00;
17'h63b4:	data_out=16'h256;
17'h63b5:	data_out=16'h899c;
17'h63b6:	data_out=16'h9e6;
17'h63b7:	data_out=16'h4ca;
17'h63b8:	data_out=16'h247;
17'h63b9:	data_out=16'ha00;
17'h63ba:	data_out=16'h9fd;
17'h63bb:	data_out=16'h8901;
17'h63bc:	data_out=16'h7cd;
17'h63bd:	data_out=16'h9;
17'h63be:	data_out=16'h81b3;
17'h63bf:	data_out=16'h818e;
17'h63c0:	data_out=16'h89dd;
17'h63c1:	data_out=16'h37f;
17'h63c2:	data_out=16'h540;
17'h63c3:	data_out=16'h8341;
17'h63c4:	data_out=16'h837d;
17'h63c5:	data_out=16'h8684;
17'h63c6:	data_out=16'h7a7;
17'h63c7:	data_out=16'h37b;
17'h63c8:	data_out=16'ha00;
17'h63c9:	data_out=16'h14b;
17'h63ca:	data_out=16'h176;
17'h63cb:	data_out=16'h9f8;
17'h63cc:	data_out=16'h5c4;
17'h63cd:	data_out=16'h985;
17'h63ce:	data_out=16'h940;
17'h63cf:	data_out=16'h407;
17'h63d0:	data_out=16'h88ac;
17'h63d1:	data_out=16'h8a00;
17'h63d2:	data_out=16'h8a00;
17'h63d3:	data_out=16'ha00;
17'h63d4:	data_out=16'ha00;
17'h63d5:	data_out=16'h88e8;
17'h63d6:	data_out=16'h8517;
17'h63d7:	data_out=16'h8331;
17'h63d8:	data_out=16'h85a0;
17'h63d9:	data_out=16'h875c;
17'h63da:	data_out=16'ha00;
17'h63db:	data_out=16'h882b;
17'h63dc:	data_out=16'h9ff;
17'h63dd:	data_out=16'h8e2;
17'h63de:	data_out=16'ha00;
17'h63df:	data_out=16'h77d;
17'h63e0:	data_out=16'h8a00;
17'h63e1:	data_out=16'h8866;
17'h63e2:	data_out=16'h9f7;
17'h63e3:	data_out=16'ha00;
17'h63e4:	data_out=16'h3ed;
17'h63e5:	data_out=16'ha00;
17'h63e6:	data_out=16'h34a;
17'h63e7:	data_out=16'h707;
17'h63e8:	data_out=16'h822d;
17'h63e9:	data_out=16'h80bd;
17'h63ea:	data_out=16'h831a;
17'h63eb:	data_out=16'h83e7;
17'h63ec:	data_out=16'h7f2;
17'h63ed:	data_out=16'ha00;
17'h63ee:	data_out=16'h8305;
17'h63ef:	data_out=16'h81c2;
17'h63f0:	data_out=16'h82b7;
17'h63f1:	data_out=16'h2b2;
17'h63f2:	data_out=16'h89ff;
17'h63f3:	data_out=16'h8582;
17'h63f4:	data_out=16'h8a00;
17'h63f5:	data_out=16'h8005;
17'h63f6:	data_out=16'h4f9;
17'h63f7:	data_out=16'h89ce;
17'h63f8:	data_out=16'h8538;
17'h63f9:	data_out=16'h7d7;
17'h63fa:	data_out=16'ha00;
17'h63fb:	data_out=16'h819d;
17'h63fc:	data_out=16'h256;
17'h63fd:	data_out=16'h12d;
17'h63fe:	data_out=16'h8395;
17'h63ff:	data_out=16'h89f3;
17'h6400:	data_out=16'h8a00;
17'h6401:	data_out=16'h8138;
17'h6402:	data_out=16'h404;
17'h6403:	data_out=16'h8939;
17'h6404:	data_out=16'h524;
17'h6405:	data_out=16'h9ff;
17'h6406:	data_out=16'ha00;
17'h6407:	data_out=16'h9fe;
17'h6408:	data_out=16'h89c5;
17'h6409:	data_out=16'h8942;
17'h640a:	data_out=16'h8a00;
17'h640b:	data_out=16'h9fb;
17'h640c:	data_out=16'h2fe;
17'h640d:	data_out=16'h142;
17'h640e:	data_out=16'h84f8;
17'h640f:	data_out=16'h696;
17'h6410:	data_out=16'h89ef;
17'h6411:	data_out=16'h9f6;
17'h6412:	data_out=16'h9f0;
17'h6413:	data_out=16'h84e4;
17'h6414:	data_out=16'h9fb;
17'h6415:	data_out=16'h8a00;
17'h6416:	data_out=16'h89ff;
17'h6417:	data_out=16'h9ee;
17'h6418:	data_out=16'h8631;
17'h6419:	data_out=16'ha00;
17'h641a:	data_out=16'h9fd;
17'h641b:	data_out=16'h9df;
17'h641c:	data_out=16'h6a4;
17'h641d:	data_out=16'h5d5;
17'h641e:	data_out=16'h9d1;
17'h641f:	data_out=16'h6d9;
17'h6420:	data_out=16'h9f3;
17'h6421:	data_out=16'h8454;
17'h6422:	data_out=16'h81f6;
17'h6423:	data_out=16'h8a00;
17'h6424:	data_out=16'h8a00;
17'h6425:	data_out=16'h89f3;
17'h6426:	data_out=16'h8a00;
17'h6427:	data_out=16'h9f8;
17'h6428:	data_out=16'h8247;
17'h6429:	data_out=16'h322;
17'h642a:	data_out=16'h88e8;
17'h642b:	data_out=16'ha00;
17'h642c:	data_out=16'h89ff;
17'h642d:	data_out=16'h8a00;
17'h642e:	data_out=16'h9e8;
17'h642f:	data_out=16'h9ef;
17'h6430:	data_out=16'h872a;
17'h6431:	data_out=16'h9fb;
17'h6432:	data_out=16'h874e;
17'h6433:	data_out=16'ha00;
17'h6434:	data_out=16'h89fc;
17'h6435:	data_out=16'h85b;
17'h6436:	data_out=16'h876c;
17'h6437:	data_out=16'h711;
17'h6438:	data_out=16'ha00;
17'h6439:	data_out=16'ha00;
17'h643a:	data_out=16'h8152;
17'h643b:	data_out=16'h89cc;
17'h643c:	data_out=16'h1a7;
17'h643d:	data_out=16'h89ff;
17'h643e:	data_out=16'h8220;
17'h643f:	data_out=16'h9fe;
17'h6440:	data_out=16'h894a;
17'h6441:	data_out=16'h80d0;
17'h6442:	data_out=16'h8a00;
17'h6443:	data_out=16'ha00;
17'h6444:	data_out=16'h122;
17'h6445:	data_out=16'h8a00;
17'h6446:	data_out=16'h80d9;
17'h6447:	data_out=16'h895a;
17'h6448:	data_out=16'ha00;
17'h6449:	data_out=16'h89fc;
17'h644a:	data_out=16'ha00;
17'h644b:	data_out=16'h5e6;
17'h644c:	data_out=16'h8819;
17'h644d:	data_out=16'hb5;
17'h644e:	data_out=16'h982;
17'h644f:	data_out=16'h89f7;
17'h6450:	data_out=16'h853b;
17'h6451:	data_out=16'h891b;
17'h6452:	data_out=16'h8a00;
17'h6453:	data_out=16'ha00;
17'h6454:	data_out=16'h9ee;
17'h6455:	data_out=16'h89f3;
17'h6456:	data_out=16'h8a00;
17'h6457:	data_out=16'h89ff;
17'h6458:	data_out=16'h89f6;
17'h6459:	data_out=16'h89e4;
17'h645a:	data_out=16'h9f6;
17'h645b:	data_out=16'h7db;
17'h645c:	data_out=16'h9f7;
17'h645d:	data_out=16'h88c6;
17'h645e:	data_out=16'h9f2;
17'h645f:	data_out=16'h5f9;
17'h6460:	data_out=16'h8a00;
17'h6461:	data_out=16'h3c7;
17'h6462:	data_out=16'h99a;
17'h6463:	data_out=16'ha00;
17'h6464:	data_out=16'h804d;
17'h6465:	data_out=16'h9fe;
17'h6466:	data_out=16'ha00;
17'h6467:	data_out=16'ha00;
17'h6468:	data_out=16'h83b5;
17'h6469:	data_out=16'h8a00;
17'h646a:	data_out=16'h856c;
17'h646b:	data_out=16'h9fc;
17'h646c:	data_out=16'h8a00;
17'h646d:	data_out=16'ha00;
17'h646e:	data_out=16'h856b;
17'h646f:	data_out=16'h58e;
17'h6470:	data_out=16'h8528;
17'h6471:	data_out=16'h9ed;
17'h6472:	data_out=16'h89ec;
17'h6473:	data_out=16'h105;
17'h6474:	data_out=16'h87b2;
17'h6475:	data_out=16'h940;
17'h6476:	data_out=16'ha00;
17'h6477:	data_out=16'h89fc;
17'h6478:	data_out=16'h9f6;
17'h6479:	data_out=16'h44a;
17'h647a:	data_out=16'ha00;
17'h647b:	data_out=16'h81f4;
17'h647c:	data_out=16'h4ba;
17'h647d:	data_out=16'ha00;
17'h647e:	data_out=16'h899e;
17'h647f:	data_out=16'h8776;
17'h6480:	data_out=16'h8a00;
17'h6481:	data_out=16'h9c8;
17'h6482:	data_out=16'h98e;
17'h6483:	data_out=16'h89fe;
17'h6484:	data_out=16'h9ea;
17'h6485:	data_out=16'h9f5;
17'h6486:	data_out=16'ha00;
17'h6487:	data_out=16'ha00;
17'h6488:	data_out=16'h8319;
17'h6489:	data_out=16'h877e;
17'h648a:	data_out=16'h8a00;
17'h648b:	data_out=16'h9fb;
17'h648c:	data_out=16'h9e7;
17'h648d:	data_out=16'h84c7;
17'h648e:	data_out=16'h8450;
17'h648f:	data_out=16'h9ed;
17'h6490:	data_out=16'h89f3;
17'h6491:	data_out=16'h9e5;
17'h6492:	data_out=16'h9fd;
17'h6493:	data_out=16'h89f4;
17'h6494:	data_out=16'h9f6;
17'h6495:	data_out=16'h8a00;
17'h6496:	data_out=16'h89fd;
17'h6497:	data_out=16'h9ee;
17'h6498:	data_out=16'h45d;
17'h6499:	data_out=16'h9fc;
17'h649a:	data_out=16'h9f4;
17'h649b:	data_out=16'h9cf;
17'h649c:	data_out=16'h81b0;
17'h649d:	data_out=16'h9e8;
17'h649e:	data_out=16'h9ed;
17'h649f:	data_out=16'ha00;
17'h64a0:	data_out=16'h9e0;
17'h64a1:	data_out=16'h8380;
17'h64a2:	data_out=16'h979;
17'h64a3:	data_out=16'h8a00;
17'h64a4:	data_out=16'h8a00;
17'h64a5:	data_out=16'h89e4;
17'h64a6:	data_out=16'h8a00;
17'h64a7:	data_out=16'h9f6;
17'h64a8:	data_out=16'h822d;
17'h64a9:	data_out=16'h8520;
17'h64aa:	data_out=16'h5fb;
17'h64ab:	data_out=16'ha00;
17'h64ac:	data_out=16'h89fe;
17'h64ad:	data_out=16'h8a00;
17'h64ae:	data_out=16'ha00;
17'h64af:	data_out=16'h9e9;
17'h64b0:	data_out=16'h844a;
17'h64b1:	data_out=16'h9eb;
17'h64b2:	data_out=16'h8428;
17'h64b3:	data_out=16'ha00;
17'h64b4:	data_out=16'h880d;
17'h64b5:	data_out=16'h909;
17'h64b6:	data_out=16'h4ea;
17'h64b7:	data_out=16'h9ec;
17'h64b8:	data_out=16'h9ec;
17'h64b9:	data_out=16'ha00;
17'h64ba:	data_out=16'h9e9;
17'h64bb:	data_out=16'h83b8;
17'h64bc:	data_out=16'h80e8;
17'h64bd:	data_out=16'h8934;
17'h64be:	data_out=16'h8224;
17'h64bf:	data_out=16'h9f5;
17'h64c0:	data_out=16'h857d;
17'h64c1:	data_out=16'h625;
17'h64c2:	data_out=16'h8a00;
17'h64c3:	data_out=16'h810;
17'h64c4:	data_out=16'h9f7;
17'h64c5:	data_out=16'h8a00;
17'h64c6:	data_out=16'h80f2;
17'h64c7:	data_out=16'h63f;
17'h64c8:	data_out=16'ha00;
17'h64c9:	data_out=16'h89f7;
17'h64ca:	data_out=16'ha00;
17'h64cb:	data_out=16'h2c0;
17'h64cc:	data_out=16'h87bb;
17'h64cd:	data_out=16'h9f3;
17'h64ce:	data_out=16'ha00;
17'h64cf:	data_out=16'h8569;
17'h64d0:	data_out=16'h133;
17'h64d1:	data_out=16'h89ed;
17'h64d2:	data_out=16'h89fd;
17'h64d3:	data_out=16'ha00;
17'h64d4:	data_out=16'h9e1;
17'h64d5:	data_out=16'h89e7;
17'h64d6:	data_out=16'h8a00;
17'h64d7:	data_out=16'h89f3;
17'h64d8:	data_out=16'h89f0;
17'h64d9:	data_out=16'h89da;
17'h64da:	data_out=16'h9fc;
17'h64db:	data_out=16'h853;
17'h64dc:	data_out=16'h9eb;
17'h64dd:	data_out=16'h63b;
17'h64de:	data_out=16'h9e3;
17'h64df:	data_out=16'h9fc;
17'h64e0:	data_out=16'h8a00;
17'h64e1:	data_out=16'h9ce;
17'h64e2:	data_out=16'h9df;
17'h64e3:	data_out=16'ha00;
17'h64e4:	data_out=16'h81f0;
17'h64e5:	data_out=16'h9f5;
17'h64e6:	data_out=16'ha00;
17'h64e7:	data_out=16'h9fd;
17'h64e8:	data_out=16'h82eb;
17'h64e9:	data_out=16'h89fb;
17'h64ea:	data_out=16'h8503;
17'h64eb:	data_out=16'h9f2;
17'h64ec:	data_out=16'h8a00;
17'h64ed:	data_out=16'ha00;
17'h64ee:	data_out=16'h8500;
17'h64ef:	data_out=16'h209;
17'h64f0:	data_out=16'h849c;
17'h64f1:	data_out=16'ha00;
17'h64f2:	data_out=16'h89e6;
17'h64f3:	data_out=16'h89f1;
17'h64f4:	data_out=16'h8502;
17'h64f5:	data_out=16'h430;
17'h64f6:	data_out=16'ha00;
17'h64f7:	data_out=16'h89ea;
17'h64f8:	data_out=16'h7c0;
17'h64f9:	data_out=16'h9d4;
17'h64fa:	data_out=16'ha00;
17'h64fb:	data_out=16'h8220;
17'h64fc:	data_out=16'ha00;
17'h64fd:	data_out=16'ha00;
17'h64fe:	data_out=16'h898b;
17'h64ff:	data_out=16'h8173;
17'h6500:	data_out=16'h8a00;
17'h6501:	data_out=16'h9cc;
17'h6502:	data_out=16'h9e2;
17'h6503:	data_out=16'h8a00;
17'h6504:	data_out=16'h9ef;
17'h6505:	data_out=16'h9fc;
17'h6506:	data_out=16'h8502;
17'h6507:	data_out=16'h9fd;
17'h6508:	data_out=16'h35f;
17'h6509:	data_out=16'h8913;
17'h650a:	data_out=16'h8a00;
17'h650b:	data_out=16'h9fa;
17'h650c:	data_out=16'h89b1;
17'h650d:	data_out=16'h89ed;
17'h650e:	data_out=16'h564;
17'h650f:	data_out=16'ha00;
17'h6510:	data_out=16'h89fd;
17'h6511:	data_out=16'h9e4;
17'h6512:	data_out=16'h9f6;
17'h6513:	data_out=16'h89f0;
17'h6514:	data_out=16'h9c9;
17'h6515:	data_out=16'h89fc;
17'h6516:	data_out=16'h89fc;
17'h6517:	data_out=16'h70a;
17'h6518:	data_out=16'ha00;
17'h6519:	data_out=16'h9f6;
17'h651a:	data_out=16'h9ff;
17'h651b:	data_out=16'h95f;
17'h651c:	data_out=16'h8034;
17'h651d:	data_out=16'h9dd;
17'h651e:	data_out=16'h9f8;
17'h651f:	data_out=16'ha00;
17'h6520:	data_out=16'h9e7;
17'h6521:	data_out=16'h618;
17'h6522:	data_out=16'ha00;
17'h6523:	data_out=16'h8a00;
17'h6524:	data_out=16'h8a00;
17'h6525:	data_out=16'h89d9;
17'h6526:	data_out=16'h8a00;
17'h6527:	data_out=16'h9ee;
17'h6528:	data_out=16'h786;
17'h6529:	data_out=16'h8168;
17'h652a:	data_out=16'h9fe;
17'h652b:	data_out=16'ha00;
17'h652c:	data_out=16'h89fd;
17'h652d:	data_out=16'h16f;
17'h652e:	data_out=16'ha00;
17'h652f:	data_out=16'h9df;
17'h6530:	data_out=16'hca;
17'h6531:	data_out=16'h8e2;
17'h6532:	data_out=16'h183;
17'h6533:	data_out=16'ha00;
17'h6534:	data_out=16'h853d;
17'h6535:	data_out=16'h959;
17'h6536:	data_out=16'h9f3;
17'h6537:	data_out=16'h9fc;
17'h6538:	data_out=16'h9f1;
17'h6539:	data_out=16'ha00;
17'h653a:	data_out=16'h9eb;
17'h653b:	data_out=16'h874d;
17'h653c:	data_out=16'h10d;
17'h653d:	data_out=16'h92e;
17'h653e:	data_out=16'h790;
17'h653f:	data_out=16'h9fc;
17'h6540:	data_out=16'h92;
17'h6541:	data_out=16'h8403;
17'h6542:	data_out=16'h8a00;
17'h6543:	data_out=16'h89b0;
17'h6544:	data_out=16'ha00;
17'h6545:	data_out=16'h89fc;
17'h6546:	data_out=16'h797;
17'h6547:	data_out=16'h19e;
17'h6548:	data_out=16'ha00;
17'h6549:	data_out=16'h89ed;
17'h654a:	data_out=16'ha00;
17'h654b:	data_out=16'h8575;
17'h654c:	data_out=16'h89f1;
17'h654d:	data_out=16'ha00;
17'h654e:	data_out=16'ha00;
17'h654f:	data_out=16'h86fb;
17'h6550:	data_out=16'h98a;
17'h6551:	data_out=16'h89e3;
17'h6552:	data_out=16'h89ff;
17'h6553:	data_out=16'ha00;
17'h6554:	data_out=16'h9e9;
17'h6555:	data_out=16'h89c2;
17'h6556:	data_out=16'h89ff;
17'h6557:	data_out=16'h8985;
17'h6558:	data_out=16'h89e2;
17'h6559:	data_out=16'h843b;
17'h655a:	data_out=16'h9ed;
17'h655b:	data_out=16'h9fb;
17'h655c:	data_out=16'h997;
17'h655d:	data_out=16'h9cc;
17'h655e:	data_out=16'h9b7;
17'h655f:	data_out=16'ha00;
17'h6560:	data_out=16'h89ff;
17'h6561:	data_out=16'h9d5;
17'h6562:	data_out=16'h49c;
17'h6563:	data_out=16'ha00;
17'h6564:	data_out=16'h21;
17'h6565:	data_out=16'h9ee;
17'h6566:	data_out=16'ha00;
17'h6567:	data_out=16'ha00;
17'h6568:	data_out=16'h6ac;
17'h6569:	data_out=16'h8714;
17'h656a:	data_out=16'h4e1;
17'h656b:	data_out=16'h9f7;
17'h656c:	data_out=16'h8a00;
17'h656d:	data_out=16'ha00;
17'h656e:	data_out=16'h4e3;
17'h656f:	data_out=16'hc4;
17'h6570:	data_out=16'h52a;
17'h6571:	data_out=16'ha00;
17'h6572:	data_out=16'h8682;
17'h6573:	data_out=16'h4e;
17'h6574:	data_out=16'h800c;
17'h6575:	data_out=16'h89d7;
17'h6576:	data_out=16'ha00;
17'h6577:	data_out=16'h8955;
17'h6578:	data_out=16'h8423;
17'h6579:	data_out=16'ha00;
17'h657a:	data_out=16'ha00;
17'h657b:	data_out=16'h792;
17'h657c:	data_out=16'ha00;
17'h657d:	data_out=16'ha00;
17'h657e:	data_out=16'h8995;
17'h657f:	data_out=16'h9e1;
17'h6580:	data_out=16'h89f8;
17'h6581:	data_out=16'h9f6;
17'h6582:	data_out=16'h9e2;
17'h6583:	data_out=16'h89ff;
17'h6584:	data_out=16'h9ff;
17'h6585:	data_out=16'ha00;
17'h6586:	data_out=16'h899d;
17'h6587:	data_out=16'h340;
17'h6588:	data_out=16'h9e5;
17'h6589:	data_out=16'h89fd;
17'h658a:	data_out=16'h89e4;
17'h658b:	data_out=16'h8900;
17'h658c:	data_out=16'h88bd;
17'h658d:	data_out=16'h89fe;
17'h658e:	data_out=16'h9ff;
17'h658f:	data_out=16'ha00;
17'h6590:	data_out=16'h89fc;
17'h6591:	data_out=16'h9e7;
17'h6592:	data_out=16'h9da;
17'h6593:	data_out=16'h89fa;
17'h6594:	data_out=16'h86da;
17'h6595:	data_out=16'h89f7;
17'h6596:	data_out=16'h89f5;
17'h6597:	data_out=16'h8987;
17'h6598:	data_out=16'h9fc;
17'h6599:	data_out=16'h9fa;
17'h659a:	data_out=16'ha00;
17'h659b:	data_out=16'h59;
17'h659c:	data_out=16'h89f9;
17'h659d:	data_out=16'h9dc;
17'h659e:	data_out=16'h3fe;
17'h659f:	data_out=16'h85fd;
17'h65a0:	data_out=16'h99a;
17'h65a1:	data_out=16'ha00;
17'h65a2:	data_out=16'ha00;
17'h65a3:	data_out=16'h89ff;
17'h65a4:	data_out=16'h89ff;
17'h65a5:	data_out=16'h89ef;
17'h65a6:	data_out=16'h89f8;
17'h65a7:	data_out=16'h9da;
17'h65a8:	data_out=16'ha00;
17'h65a9:	data_out=16'h690;
17'h65aa:	data_out=16'ha00;
17'h65ab:	data_out=16'ha00;
17'h65ac:	data_out=16'h89f6;
17'h65ad:	data_out=16'h9f4;
17'h65ae:	data_out=16'ha00;
17'h65af:	data_out=16'h9d6;
17'h65b0:	data_out=16'h9ff;
17'h65b1:	data_out=16'h82a7;
17'h65b2:	data_out=16'h9dc;
17'h65b3:	data_out=16'h4de;
17'h65b4:	data_out=16'h201;
17'h65b5:	data_out=16'h5bc;
17'h65b6:	data_out=16'ha00;
17'h65b7:	data_out=16'h9fa;
17'h65b8:	data_out=16'h9ee;
17'h65b9:	data_out=16'h5cd;
17'h65ba:	data_out=16'h800b;
17'h65bb:	data_out=16'h8516;
17'h65bc:	data_out=16'h8668;
17'h65bd:	data_out=16'h8188;
17'h65be:	data_out=16'ha00;
17'h65bf:	data_out=16'h9ac;
17'h65c0:	data_out=16'h336;
17'h65c1:	data_out=16'h89df;
17'h65c2:	data_out=16'h89fd;
17'h65c3:	data_out=16'h88d9;
17'h65c4:	data_out=16'h85ee;
17'h65c5:	data_out=16'h89f7;
17'h65c6:	data_out=16'ha00;
17'h65c7:	data_out=16'h85a6;
17'h65c8:	data_out=16'h93c;
17'h65c9:	data_out=16'h89f8;
17'h65ca:	data_out=16'ha00;
17'h65cb:	data_out=16'h89ff;
17'h65cc:	data_out=16'h89ee;
17'h65cd:	data_out=16'ha00;
17'h65ce:	data_out=16'ha00;
17'h65cf:	data_out=16'h8513;
17'h65d0:	data_out=16'h1cd;
17'h65d1:	data_out=16'h89ec;
17'h65d2:	data_out=16'h89f9;
17'h65d3:	data_out=16'ha00;
17'h65d4:	data_out=16'h9d1;
17'h65d5:	data_out=16'h89dd;
17'h65d6:	data_out=16'h89fd;
17'h65d7:	data_out=16'h89dd;
17'h65d8:	data_out=16'h89ec;
17'h65d9:	data_out=16'h146;
17'h65da:	data_out=16'h209;
17'h65db:	data_out=16'h9fa;
17'h65dc:	data_out=16'h922;
17'h65dd:	data_out=16'h9ec;
17'h65de:	data_out=16'h987;
17'h65df:	data_out=16'ha00;
17'h65e0:	data_out=16'h89c7;
17'h65e1:	data_out=16'h1c1;
17'h65e2:	data_out=16'h8953;
17'h65e3:	data_out=16'h7fe;
17'h65e4:	data_out=16'h8a00;
17'h65e5:	data_out=16'h8678;
17'h65e6:	data_out=16'h9fc;
17'h65e7:	data_out=16'h9fd;
17'h65e8:	data_out=16'ha00;
17'h65e9:	data_out=16'h88b5;
17'h65ea:	data_out=16'h9ff;
17'h65eb:	data_out=16'h6a9;
17'h65ec:	data_out=16'h944;
17'h65ed:	data_out=16'h7f5;
17'h65ee:	data_out=16'h9ff;
17'h65ef:	data_out=16'h110;
17'h65f0:	data_out=16'h9ff;
17'h65f1:	data_out=16'ha00;
17'h65f2:	data_out=16'h8538;
17'h65f3:	data_out=16'h21a;
17'h65f4:	data_out=16'h9fc;
17'h65f5:	data_out=16'h89e6;
17'h65f6:	data_out=16'ha00;
17'h65f7:	data_out=16'h89f2;
17'h65f8:	data_out=16'h44d;
17'h65f9:	data_out=16'h9ff;
17'h65fa:	data_out=16'h214;
17'h65fb:	data_out=16'ha00;
17'h65fc:	data_out=16'ha00;
17'h65fd:	data_out=16'h696;
17'h65fe:	data_out=16'h89f9;
17'h65ff:	data_out=16'h777;
17'h6600:	data_out=16'h64f;
17'h6601:	data_out=16'h9eb;
17'h6602:	data_out=16'h9df;
17'h6603:	data_out=16'h89ed;
17'h6604:	data_out=16'h9ff;
17'h6605:	data_out=16'h8734;
17'h6606:	data_out=16'h89eb;
17'h6607:	data_out=16'h89db;
17'h6608:	data_out=16'h9d1;
17'h6609:	data_out=16'h89fc;
17'h660a:	data_out=16'h89e3;
17'h660b:	data_out=16'h88d2;
17'h660c:	data_out=16'h897c;
17'h660d:	data_out=16'h8a00;
17'h660e:	data_out=16'ha00;
17'h660f:	data_out=16'h9fc;
17'h6610:	data_out=16'h89e8;
17'h6611:	data_out=16'h8771;
17'h6612:	data_out=16'h9b5;
17'h6613:	data_out=16'h89f7;
17'h6614:	data_out=16'h89d8;
17'h6615:	data_out=16'h89f3;
17'h6616:	data_out=16'h89f4;
17'h6617:	data_out=16'h89cd;
17'h6618:	data_out=16'h9f4;
17'h6619:	data_out=16'ha00;
17'h661a:	data_out=16'ha00;
17'h661b:	data_out=16'h89e5;
17'h661c:	data_out=16'h89ea;
17'h661d:	data_out=16'h858f;
17'h661e:	data_out=16'h86a7;
17'h661f:	data_out=16'h8837;
17'h6620:	data_out=16'h9ad;
17'h6621:	data_out=16'ha00;
17'h6622:	data_out=16'ha00;
17'h6623:	data_out=16'h8a00;
17'h6624:	data_out=16'h8a00;
17'h6625:	data_out=16'h89d4;
17'h6626:	data_out=16'h8966;
17'h6627:	data_out=16'h669;
17'h6628:	data_out=16'ha00;
17'h6629:	data_out=16'h9e4;
17'h662a:	data_out=16'h9fe;
17'h662b:	data_out=16'ha00;
17'h662c:	data_out=16'h89f4;
17'h662d:	data_out=16'ha00;
17'h662e:	data_out=16'h9e8;
17'h662f:	data_out=16'h95f;
17'h6630:	data_out=16'h22d;
17'h6631:	data_out=16'h89f3;
17'h6632:	data_out=16'h80be;
17'h6633:	data_out=16'h891f;
17'h6634:	data_out=16'h8333;
17'h6635:	data_out=16'h878;
17'h6636:	data_out=16'h9fd;
17'h6637:	data_out=16'h9fa;
17'h6638:	data_out=16'h483;
17'h6639:	data_out=16'h84b9;
17'h663a:	data_out=16'h89fa;
17'h663b:	data_out=16'h86d1;
17'h663c:	data_out=16'h8984;
17'h663d:	data_out=16'h973;
17'h663e:	data_out=16'ha00;
17'h663f:	data_out=16'h872b;
17'h6640:	data_out=16'h8066;
17'h6641:	data_out=16'h88b7;
17'h6642:	data_out=16'h89f1;
17'h6643:	data_out=16'h80c1;
17'h6644:	data_out=16'h870f;
17'h6645:	data_out=16'h89f4;
17'h6646:	data_out=16'ha00;
17'h6647:	data_out=16'h838c;
17'h6648:	data_out=16'h8485;
17'h6649:	data_out=16'h89da;
17'h664a:	data_out=16'h9e6;
17'h664b:	data_out=16'h8a00;
17'h664c:	data_out=16'h89e3;
17'h664d:	data_out=16'ha00;
17'h664e:	data_out=16'ha00;
17'h664f:	data_out=16'h89f2;
17'h6650:	data_out=16'h89f0;
17'h6651:	data_out=16'h89ee;
17'h6652:	data_out=16'h89eb;
17'h6653:	data_out=16'h9e4;
17'h6654:	data_out=16'h9be;
17'h6655:	data_out=16'h89d7;
17'h6656:	data_out=16'h1b3;
17'h6657:	data_out=16'h806f;
17'h6658:	data_out=16'h89f3;
17'h6659:	data_out=16'h911;
17'h665a:	data_out=16'h89ee;
17'h665b:	data_out=16'h9ff;
17'h665c:	data_out=16'h84c4;
17'h665d:	data_out=16'ha00;
17'h665e:	data_out=16'h4ef;
17'h665f:	data_out=16'h9fd;
17'h6660:	data_out=16'h893a;
17'h6661:	data_out=16'h2f;
17'h6662:	data_out=16'h89b6;
17'h6663:	data_out=16'h88d1;
17'h6664:	data_out=16'h89ee;
17'h6665:	data_out=16'h8886;
17'h6666:	data_out=16'ha00;
17'h6667:	data_out=16'ha00;
17'h6668:	data_out=16'ha00;
17'h6669:	data_out=16'h6c7;
17'h666a:	data_out=16'ha00;
17'h666b:	data_out=16'h89c1;
17'h666c:	data_out=16'h9e1;
17'h666d:	data_out=16'h883c;
17'h666e:	data_out=16'ha00;
17'h666f:	data_out=16'h872d;
17'h6670:	data_out=16'ha00;
17'h6671:	data_out=16'h9f0;
17'h6672:	data_out=16'h89c5;
17'h6673:	data_out=16'h895d;
17'h6674:	data_out=16'h149;
17'h6675:	data_out=16'h89f4;
17'h6676:	data_out=16'ha00;
17'h6677:	data_out=16'h89e7;
17'h6678:	data_out=16'ha00;
17'h6679:	data_out=16'h9ff;
17'h667a:	data_out=16'h89ac;
17'h667b:	data_out=16'ha00;
17'h667c:	data_out=16'h9fc;
17'h667d:	data_out=16'h818c;
17'h667e:	data_out=16'h89dc;
17'h667f:	data_out=16'h649;
17'h6680:	data_out=16'h9a5;
17'h6681:	data_out=16'h22d;
17'h6682:	data_out=16'h9fc;
17'h6683:	data_out=16'h89a4;
17'h6684:	data_out=16'h9e5;
17'h6685:	data_out=16'h88d9;
17'h6686:	data_out=16'h8a00;
17'h6687:	data_out=16'h89f5;
17'h6688:	data_out=16'h9e7;
17'h6689:	data_out=16'h89f9;
17'h668a:	data_out=16'h89ed;
17'h668b:	data_out=16'h8737;
17'h668c:	data_out=16'h896f;
17'h668d:	data_out=16'h89fc;
17'h668e:	data_out=16'h9ff;
17'h668f:	data_out=16'h9fc;
17'h6690:	data_out=16'h89e3;
17'h6691:	data_out=16'h8981;
17'h6692:	data_out=16'h3f6;
17'h6693:	data_out=16'h89e1;
17'h6694:	data_out=16'h8901;
17'h6695:	data_out=16'h8892;
17'h6696:	data_out=16'h89a7;
17'h6697:	data_out=16'h8927;
17'h6698:	data_out=16'h9ec;
17'h6699:	data_out=16'h9fe;
17'h669a:	data_out=16'h82c2;
17'h669b:	data_out=16'h8946;
17'h669c:	data_out=16'h897d;
17'h669d:	data_out=16'h88f3;
17'h669e:	data_out=16'h88a2;
17'h669f:	data_out=16'h8826;
17'h66a0:	data_out=16'h9ca;
17'h66a1:	data_out=16'h9ff;
17'h66a2:	data_out=16'h1b6;
17'h66a3:	data_out=16'h8a00;
17'h66a4:	data_out=16'h8a00;
17'h66a5:	data_out=16'h89b4;
17'h66a6:	data_out=16'h82ab;
17'h66a7:	data_out=16'h8138;
17'h66a8:	data_out=16'ha00;
17'h66a9:	data_out=16'h9f7;
17'h66aa:	data_out=16'h9f9;
17'h66ab:	data_out=16'ha00;
17'h66ac:	data_out=16'h89aa;
17'h66ad:	data_out=16'h9ff;
17'h66ae:	data_out=16'h799;
17'h66af:	data_out=16'h895d;
17'h66b0:	data_out=16'h3f;
17'h66b1:	data_out=16'h89a9;
17'h66b2:	data_out=16'h8703;
17'h66b3:	data_out=16'h8938;
17'h66b4:	data_out=16'h840b;
17'h66b5:	data_out=16'h3cd;
17'h66b6:	data_out=16'h9fb;
17'h66b7:	data_out=16'ha00;
17'h66b8:	data_out=16'h89f4;
17'h66b9:	data_out=16'h8962;
17'h66ba:	data_out=16'h89ef;
17'h66bb:	data_out=16'h841c;
17'h66bc:	data_out=16'h8899;
17'h66bd:	data_out=16'h1cd;
17'h66be:	data_out=16'ha00;
17'h66bf:	data_out=16'h88e1;
17'h66c0:	data_out=16'h8505;
17'h66c1:	data_out=16'h8505;
17'h66c2:	data_out=16'h89d7;
17'h66c3:	data_out=16'ha00;
17'h66c4:	data_out=16'h870e;
17'h66c5:	data_out=16'h88f4;
17'h66c6:	data_out=16'ha00;
17'h66c7:	data_out=16'h7d9;
17'h66c8:	data_out=16'h89f8;
17'h66c9:	data_out=16'h89aa;
17'h66ca:	data_out=16'h9e6;
17'h66cb:	data_out=16'h8a00;
17'h66cc:	data_out=16'h89ea;
17'h66cd:	data_out=16'h961;
17'h66ce:	data_out=16'ha00;
17'h66cf:	data_out=16'h89fc;
17'h66d0:	data_out=16'h89a3;
17'h66d1:	data_out=16'h89d5;
17'h66d2:	data_out=16'h89f0;
17'h66d3:	data_out=16'h9b9;
17'h66d4:	data_out=16'h4da;
17'h66d5:	data_out=16'h896a;
17'h66d6:	data_out=16'h81c6;
17'h66d7:	data_out=16'h8336;
17'h66d8:	data_out=16'h89de;
17'h66d9:	data_out=16'h88ee;
17'h66da:	data_out=16'h89d9;
17'h66db:	data_out=16'h80d3;
17'h66dc:	data_out=16'h89f9;
17'h66dd:	data_out=16'ha00;
17'h66de:	data_out=16'h89c4;
17'h66df:	data_out=16'h9f6;
17'h66e0:	data_out=16'h88ce;
17'h66e1:	data_out=16'h864a;
17'h66e2:	data_out=16'h8907;
17'h66e3:	data_out=16'h892f;
17'h66e4:	data_out=16'h899f;
17'h66e5:	data_out=16'h88b5;
17'h66e6:	data_out=16'ha00;
17'h66e7:	data_out=16'ha00;
17'h66e8:	data_out=16'h9ff;
17'h66e9:	data_out=16'h9a6;
17'h66ea:	data_out=16'h9ff;
17'h66eb:	data_out=16'h8928;
17'h66ec:	data_out=16'h9f2;
17'h66ed:	data_out=16'h892b;
17'h66ee:	data_out=16'h9ff;
17'h66ef:	data_out=16'h86d4;
17'h66f0:	data_out=16'h9ff;
17'h66f1:	data_out=16'h9f1;
17'h66f2:	data_out=16'h8995;
17'h66f3:	data_out=16'h891b;
17'h66f4:	data_out=16'h80b4;
17'h66f5:	data_out=16'h89fe;
17'h66f6:	data_out=16'ha00;
17'h66f7:	data_out=16'h89bd;
17'h66f8:	data_out=16'h9ff;
17'h66f9:	data_out=16'h9ff;
17'h66fa:	data_out=16'h890d;
17'h66fb:	data_out=16'ha00;
17'h66fc:	data_out=16'h9f3;
17'h66fd:	data_out=16'h8561;
17'h66fe:	data_out=16'h89d3;
17'h66ff:	data_out=16'h819f;
17'h6700:	data_out=16'h9f6;
17'h6701:	data_out=16'h9af;
17'h6702:	data_out=16'h238;
17'h6703:	data_out=16'h8805;
17'h6704:	data_out=16'h8836;
17'h6705:	data_out=16'h88bc;
17'h6706:	data_out=16'h8a00;
17'h6707:	data_out=16'h8a00;
17'h6708:	data_out=16'h9df;
17'h6709:	data_out=16'h8a00;
17'h670a:	data_out=16'h89f5;
17'h670b:	data_out=16'h885d;
17'h670c:	data_out=16'h8a00;
17'h670d:	data_out=16'h89d9;
17'h670e:	data_out=16'h9ff;
17'h670f:	data_out=16'h2af;
17'h6710:	data_out=16'h89d6;
17'h6711:	data_out=16'h89f6;
17'h6712:	data_out=16'h887e;
17'h6713:	data_out=16'h89b9;
17'h6714:	data_out=16'h8880;
17'h6715:	data_out=16'h3f8;
17'h6716:	data_out=16'h8904;
17'h6717:	data_out=16'h8892;
17'h6718:	data_out=16'h9e3;
17'h6719:	data_out=16'h9f4;
17'h671a:	data_out=16'h86ca;
17'h671b:	data_out=16'h896c;
17'h671c:	data_out=16'h8691;
17'h671d:	data_out=16'h897e;
17'h671e:	data_out=16'h87f6;
17'h671f:	data_out=16'h88f9;
17'h6720:	data_out=16'h9df;
17'h6721:	data_out=16'h9ff;
17'h6722:	data_out=16'h881a;
17'h6723:	data_out=16'h8a00;
17'h6724:	data_out=16'h8a00;
17'h6725:	data_out=16'h89d7;
17'h6726:	data_out=16'h8205;
17'h6727:	data_out=16'h1f8;
17'h6728:	data_out=16'h9ff;
17'h6729:	data_out=16'ha00;
17'h672a:	data_out=16'h9f7;
17'h672b:	data_out=16'ha00;
17'h672c:	data_out=16'h890a;
17'h672d:	data_out=16'h5f8;
17'h672e:	data_out=16'h8966;
17'h672f:	data_out=16'h8295;
17'h6730:	data_out=16'h92;
17'h6731:	data_out=16'h8966;
17'h6732:	data_out=16'h890f;
17'h6733:	data_out=16'h88bd;
17'h6734:	data_out=16'h8f6;
17'h6735:	data_out=16'h899e;
17'h6736:	data_out=16'h9ff;
17'h6737:	data_out=16'h8835;
17'h6738:	data_out=16'h89fb;
17'h6739:	data_out=16'h8884;
17'h673a:	data_out=16'h89f7;
17'h673b:	data_out=16'h899a;
17'h673c:	data_out=16'h86c5;
17'h673d:	data_out=16'h9f7;
17'h673e:	data_out=16'h9ff;
17'h673f:	data_out=16'h88c1;
17'h6740:	data_out=16'h8848;
17'h6741:	data_out=16'ha00;
17'h6742:	data_out=16'h8a00;
17'h6743:	data_out=16'ha00;
17'h6744:	data_out=16'h87ea;
17'h6745:	data_out=16'h31b;
17'h6746:	data_out=16'ha00;
17'h6747:	data_out=16'h89e5;
17'h6748:	data_out=16'h89ff;
17'h6749:	data_out=16'h89cf;
17'h674a:	data_out=16'h9e2;
17'h674b:	data_out=16'h8a00;
17'h674c:	data_out=16'h89f2;
17'h674d:	data_out=16'h867e;
17'h674e:	data_out=16'ha00;
17'h674f:	data_out=16'h8a00;
17'h6750:	data_out=16'h895d;
17'h6751:	data_out=16'h89ae;
17'h6752:	data_out=16'h8a00;
17'h6753:	data_out=16'h891e;
17'h6754:	data_out=16'h9ca;
17'h6755:	data_out=16'h896c;
17'h6756:	data_out=16'h80df;
17'h6757:	data_out=16'h88d9;
17'h6758:	data_out=16'h89bf;
17'h6759:	data_out=16'h8946;
17'h675a:	data_out=16'h89c1;
17'h675b:	data_out=16'h2dd;
17'h675c:	data_out=16'h89d5;
17'h675d:	data_out=16'ha00;
17'h675e:	data_out=16'h8842;
17'h675f:	data_out=16'h9f6;
17'h6760:	data_out=16'h89e7;
17'h6761:	data_out=16'h8881;
17'h6762:	data_out=16'h8893;
17'h6763:	data_out=16'h890b;
17'h6764:	data_out=16'h88bf;
17'h6765:	data_out=16'h89c5;
17'h6766:	data_out=16'h9fd;
17'h6767:	data_out=16'ha00;
17'h6768:	data_out=16'h9ff;
17'h6769:	data_out=16'h950;
17'h676a:	data_out=16'h9ff;
17'h676b:	data_out=16'h890d;
17'h676c:	data_out=16'ha00;
17'h676d:	data_out=16'h88ed;
17'h676e:	data_out=16'h9ff;
17'h676f:	data_out=16'h876b;
17'h6770:	data_out=16'h9ff;
17'h6771:	data_out=16'h2c1;
17'h6772:	data_out=16'h8977;
17'h6773:	data_out=16'h88d2;
17'h6774:	data_out=16'h80d0;
17'h6775:	data_out=16'h89e0;
17'h6776:	data_out=16'h9ff;
17'h6777:	data_out=16'h89cf;
17'h6778:	data_out=16'ha00;
17'h6779:	data_out=16'ha00;
17'h677a:	data_out=16'h88b8;
17'h677b:	data_out=16'h9ff;
17'h677c:	data_out=16'h9ef;
17'h677d:	data_out=16'h8807;
17'h677e:	data_out=16'h89d6;
17'h677f:	data_out=16'h848f;
17'h6780:	data_out=16'h9f1;
17'h6781:	data_out=16'h85b;
17'h6782:	data_out=16'h8962;
17'h6783:	data_out=16'h887d;
17'h6784:	data_out=16'h8916;
17'h6785:	data_out=16'h896e;
17'h6786:	data_out=16'h8a00;
17'h6787:	data_out=16'h8a00;
17'h6788:	data_out=16'h9bc;
17'h6789:	data_out=16'h8a00;
17'h678a:	data_out=16'h8a00;
17'h678b:	data_out=16'h8422;
17'h678c:	data_out=16'h8a00;
17'h678d:	data_out=16'h89ea;
17'h678e:	data_out=16'h9fb;
17'h678f:	data_out=16'h89eb;
17'h6790:	data_out=16'h8922;
17'h6791:	data_out=16'h8a00;
17'h6792:	data_out=16'h89fb;
17'h6793:	data_out=16'h89c1;
17'h6794:	data_out=16'h88dd;
17'h6795:	data_out=16'h85d;
17'h6796:	data_out=16'h896e;
17'h6797:	data_out=16'h8943;
17'h6798:	data_out=16'h835e;
17'h6799:	data_out=16'ha00;
17'h679a:	data_out=16'h8841;
17'h679b:	data_out=16'h8987;
17'h679c:	data_out=16'h216;
17'h679d:	data_out=16'h89f8;
17'h679e:	data_out=16'h88d9;
17'h679f:	data_out=16'h897f;
17'h67a0:	data_out=16'h9e2;
17'h67a1:	data_out=16'h9c3;
17'h67a2:	data_out=16'h8632;
17'h67a3:	data_out=16'h8a00;
17'h67a4:	data_out=16'h8a00;
17'h67a5:	data_out=16'h89dd;
17'h67a6:	data_out=16'h80ea;
17'h67a7:	data_out=16'h43e;
17'h67a8:	data_out=16'h979;
17'h67a9:	data_out=16'h9f5;
17'h67aa:	data_out=16'h86ca;
17'h67ab:	data_out=16'h9da;
17'h67ac:	data_out=16'h8969;
17'h67ad:	data_out=16'h8e;
17'h67ae:	data_out=16'h89ff;
17'h67af:	data_out=16'h948;
17'h67b0:	data_out=16'h681;
17'h67b1:	data_out=16'h89c2;
17'h67b2:	data_out=16'h899e;
17'h67b3:	data_out=16'h88bd;
17'h67b4:	data_out=16'h722;
17'h67b5:	data_out=16'h8550;
17'h67b6:	data_out=16'h9e4;
17'h67b7:	data_out=16'h89d8;
17'h67b8:	data_out=16'h8a00;
17'h67b9:	data_out=16'h87f0;
17'h67ba:	data_out=16'h89fe;
17'h67bb:	data_out=16'h89f6;
17'h67bc:	data_out=16'h59d;
17'h67bd:	data_out=16'h9d9;
17'h67be:	data_out=16'h977;
17'h67bf:	data_out=16'h8970;
17'h67c0:	data_out=16'h8964;
17'h67c1:	data_out=16'h9fe;
17'h67c2:	data_out=16'h8a00;
17'h67c3:	data_out=16'ha00;
17'h67c4:	data_out=16'h614;
17'h67c5:	data_out=16'h7d0;
17'h67c6:	data_out=16'ha00;
17'h67c7:	data_out=16'h89fb;
17'h67c8:	data_out=16'h8a00;
17'h67c9:	data_out=16'h89ae;
17'h67ca:	data_out=16'h218;
17'h67cb:	data_out=16'h8a00;
17'h67cc:	data_out=16'h89ee;
17'h67cd:	data_out=16'h86b1;
17'h67ce:	data_out=16'h6b1;
17'h67cf:	data_out=16'h8a00;
17'h67d0:	data_out=16'h8939;
17'h67d1:	data_out=16'h89ea;
17'h67d2:	data_out=16'h8a00;
17'h67d3:	data_out=16'h831e;
17'h67d4:	data_out=16'h9bc;
17'h67d5:	data_out=16'h89a9;
17'h67d6:	data_out=16'h1b7;
17'h67d7:	data_out=16'h890e;
17'h67d8:	data_out=16'h89f5;
17'h67d9:	data_out=16'h895e;
17'h67da:	data_out=16'h89ec;
17'h67db:	data_out=16'h561;
17'h67dc:	data_out=16'h89fb;
17'h67dd:	data_out=16'ha00;
17'h67de:	data_out=16'h6b;
17'h67df:	data_out=16'h83b6;
17'h67e0:	data_out=16'h8a00;
17'h67e1:	data_out=16'h899f;
17'h67e2:	data_out=16'h8911;
17'h67e3:	data_out=16'h8940;
17'h67e4:	data_out=16'h82ce;
17'h67e5:	data_out=16'h89b8;
17'h67e6:	data_out=16'ha00;
17'h67e7:	data_out=16'ha00;
17'h67e8:	data_out=16'h991;
17'h67e9:	data_out=16'h93e;
17'h67ea:	data_out=16'h9fa;
17'h67eb:	data_out=16'h8931;
17'h67ec:	data_out=16'h9fb;
17'h67ed:	data_out=16'h891e;
17'h67ee:	data_out=16'h9fa;
17'h67ef:	data_out=16'h891d;
17'h67f0:	data_out=16'h9fa;
17'h67f1:	data_out=16'h89e5;
17'h67f2:	data_out=16'h897a;
17'h67f3:	data_out=16'h899b;
17'h67f4:	data_out=16'h45f;
17'h67f5:	data_out=16'h89ff;
17'h67f6:	data_out=16'h9ff;
17'h67f7:	data_out=16'h89ea;
17'h67f8:	data_out=16'h9ff;
17'h67f9:	data_out=16'ha00;
17'h67fa:	data_out=16'h890c;
17'h67fb:	data_out=16'h977;
17'h67fc:	data_out=16'h81fa;
17'h67fd:	data_out=16'h8876;
17'h67fe:	data_out=16'h89e5;
17'h67ff:	data_out=16'h8793;
17'h6800:	data_out=16'h9df;
17'h6801:	data_out=16'h992;
17'h6802:	data_out=16'h89e8;
17'h6803:	data_out=16'h7b;
17'h6804:	data_out=16'h8262;
17'h6805:	data_out=16'h8952;
17'h6806:	data_out=16'h8a00;
17'h6807:	data_out=16'h8a00;
17'h6808:	data_out=16'h9aa;
17'h6809:	data_out=16'h8a00;
17'h680a:	data_out=16'h8a00;
17'h680b:	data_out=16'h9ad;
17'h680c:	data_out=16'h8a00;
17'h680d:	data_out=16'h89d0;
17'h680e:	data_out=16'h94d;
17'h680f:	data_out=16'h89fb;
17'h6810:	data_out=16'h9c9;
17'h6811:	data_out=16'h88fc;
17'h6812:	data_out=16'h8a00;
17'h6813:	data_out=16'h89bc;
17'h6814:	data_out=16'h8780;
17'h6815:	data_out=16'h813c;
17'h6816:	data_out=16'h89aa;
17'h6817:	data_out=16'h881d;
17'h6818:	data_out=16'h8a00;
17'h6819:	data_out=16'h9f3;
17'h681a:	data_out=16'h889e;
17'h681b:	data_out=16'h8046;
17'h681c:	data_out=16'h9f3;
17'h681d:	data_out=16'h899a;
17'h681e:	data_out=16'h88dd;
17'h681f:	data_out=16'h89be;
17'h6820:	data_out=16'h9a9;
17'h6821:	data_out=16'h912;
17'h6822:	data_out=16'h84c8;
17'h6823:	data_out=16'h8a00;
17'h6824:	data_out=16'h8a00;
17'h6825:	data_out=16'h89db;
17'h6826:	data_out=16'h8491;
17'h6827:	data_out=16'h8a9;
17'h6828:	data_out=16'h933;
17'h6829:	data_out=16'h9fa;
17'h682a:	data_out=16'h88b6;
17'h682b:	data_out=16'h96b;
17'h682c:	data_out=16'h899a;
17'h682d:	data_out=16'h86cd;
17'h682e:	data_out=16'h8a00;
17'h682f:	data_out=16'h9cd;
17'h6830:	data_out=16'h8f7;
17'h6831:	data_out=16'h806d;
17'h6832:	data_out=16'h89b1;
17'h6833:	data_out=16'h87d8;
17'h6834:	data_out=16'h885;
17'h6835:	data_out=16'h42b;
17'h6836:	data_out=16'h9cb;
17'h6837:	data_out=16'h8997;
17'h6838:	data_out=16'h8a00;
17'h6839:	data_out=16'h8795;
17'h683a:	data_out=16'h8a00;
17'h683b:	data_out=16'h89df;
17'h683c:	data_out=16'h9f0;
17'h683d:	data_out=16'h9c0;
17'h683e:	data_out=16'h936;
17'h683f:	data_out=16'h8953;
17'h6840:	data_out=16'h8985;
17'h6841:	data_out=16'h9fc;
17'h6842:	data_out=16'h20e;
17'h6843:	data_out=16'ha00;
17'h6844:	data_out=16'h976;
17'h6845:	data_out=16'h8186;
17'h6846:	data_out=16'ha00;
17'h6847:	data_out=16'h8a00;
17'h6848:	data_out=16'h8a00;
17'h6849:	data_out=16'h8984;
17'h684a:	data_out=16'h82ae;
17'h684b:	data_out=16'h8a00;
17'h684c:	data_out=16'h8a00;
17'h684d:	data_out=16'h856e;
17'h684e:	data_out=16'h8155;
17'h684f:	data_out=16'h8a00;
17'h6850:	data_out=16'h8936;
17'h6851:	data_out=16'h89ce;
17'h6852:	data_out=16'h8a00;
17'h6853:	data_out=16'h8ff;
17'h6854:	data_out=16'h8d0;
17'h6855:	data_out=16'h8978;
17'h6856:	data_out=16'h234;
17'h6857:	data_out=16'h8935;
17'h6858:	data_out=16'h83ec;
17'h6859:	data_out=16'h8976;
17'h685a:	data_out=16'h89b5;
17'h685b:	data_out=16'h959;
17'h685c:	data_out=16'h9d6;
17'h685d:	data_out=16'ha00;
17'h685e:	data_out=16'h786;
17'h685f:	data_out=16'h8a00;
17'h6860:	data_out=16'h8a00;
17'h6861:	data_out=16'h89d4;
17'h6862:	data_out=16'h871b;
17'h6863:	data_out=16'h8906;
17'h6864:	data_out=16'h1e8;
17'h6865:	data_out=16'h89c2;
17'h6866:	data_out=16'h9cd;
17'h6867:	data_out=16'ha00;
17'h6868:	data_out=16'h901;
17'h6869:	data_out=16'h915;
17'h686a:	data_out=16'h95e;
17'h686b:	data_out=16'h894c;
17'h686c:	data_out=16'h9d3;
17'h686d:	data_out=16'h88bc;
17'h686e:	data_out=16'h95e;
17'h686f:	data_out=16'h8981;
17'h6870:	data_out=16'h95b;
17'h6871:	data_out=16'h89ff;
17'h6872:	data_out=16'h8993;
17'h6873:	data_out=16'h89c8;
17'h6874:	data_out=16'h61a;
17'h6875:	data_out=16'h899a;
17'h6876:	data_out=16'h9c3;
17'h6877:	data_out=16'h89d9;
17'h6878:	data_out=16'h9ff;
17'h6879:	data_out=16'h9fb;
17'h687a:	data_out=16'h87f4;
17'h687b:	data_out=16'h936;
17'h687c:	data_out=16'h8a00;
17'h687d:	data_out=16'h8924;
17'h687e:	data_out=16'h89a2;
17'h687f:	data_out=16'h89a2;
17'h6880:	data_out=16'h963;
17'h6881:	data_out=16'h839e;
17'h6882:	data_out=16'h208;
17'h6883:	data_out=16'h818b;
17'h6884:	data_out=16'h82f2;
17'h6885:	data_out=16'h89b5;
17'h6886:	data_out=16'h8a00;
17'h6887:	data_out=16'h8a00;
17'h6888:	data_out=16'h97b;
17'h6889:	data_out=16'h89ff;
17'h688a:	data_out=16'h89e9;
17'h688b:	data_out=16'h9e6;
17'h688c:	data_out=16'h8a00;
17'h688d:	data_out=16'h89ef;
17'h688e:	data_out=16'h9fd;
17'h688f:	data_out=16'h89fd;
17'h6890:	data_out=16'h9e1;
17'h6891:	data_out=16'h99b;
17'h6892:	data_out=16'h8a00;
17'h6893:	data_out=16'h89ac;
17'h6894:	data_out=16'h867a;
17'h6895:	data_out=16'h87a1;
17'h6896:	data_out=16'h89cf;
17'h6897:	data_out=16'h884f;
17'h6898:	data_out=16'h8a00;
17'h6899:	data_out=16'h9f0;
17'h689a:	data_out=16'h8926;
17'h689b:	data_out=16'h9fa;
17'h689c:	data_out=16'h9f4;
17'h689d:	data_out=16'h87dd;
17'h689e:	data_out=16'h8975;
17'h689f:	data_out=16'h89c1;
17'h68a0:	data_out=16'h895c;
17'h68a1:	data_out=16'h9fd;
17'h68a2:	data_out=16'h9dc;
17'h68a3:	data_out=16'h8a00;
17'h68a4:	data_out=16'h8a00;
17'h68a5:	data_out=16'h89a3;
17'h68a6:	data_out=16'h968;
17'h68a7:	data_out=16'h8b3;
17'h68a8:	data_out=16'h9fd;
17'h68a9:	data_out=16'ha00;
17'h68aa:	data_out=16'h8949;
17'h68ab:	data_out=16'h7c2;
17'h68ac:	data_out=16'h89be;
17'h68ad:	data_out=16'h18a;
17'h68ae:	data_out=16'h89ff;
17'h68af:	data_out=16'h8605;
17'h68b0:	data_out=16'h30a;
17'h68b1:	data_out=16'h137;
17'h68b2:	data_out=16'h89d3;
17'h68b3:	data_out=16'h8912;
17'h68b4:	data_out=16'h84cc;
17'h68b5:	data_out=16'h837;
17'h68b6:	data_out=16'h98e;
17'h68b7:	data_out=16'h520;
17'h68b8:	data_out=16'h8a00;
17'h68b9:	data_out=16'h89a9;
17'h68ba:	data_out=16'h89fb;
17'h68bb:	data_out=16'h89fd;
17'h68bc:	data_out=16'h9ff;
17'h68bd:	data_out=16'h8201;
17'h68be:	data_out=16'h9fd;
17'h68bf:	data_out=16'h89b3;
17'h68c0:	data_out=16'h899d;
17'h68c1:	data_out=16'h9e7;
17'h68c2:	data_out=16'h901;
17'h68c3:	data_out=16'ha00;
17'h68c4:	data_out=16'h999;
17'h68c5:	data_out=16'h87e9;
17'h68c6:	data_out=16'ha00;
17'h68c7:	data_out=16'h8a00;
17'h68c8:	data_out=16'h8a00;
17'h68c9:	data_out=16'h8897;
17'h68ca:	data_out=16'h89fc;
17'h68cb:	data_out=16'h770;
17'h68cc:	data_out=16'h89fe;
17'h68cd:	data_out=16'h513;
17'h68ce:	data_out=16'h86ea;
17'h68cf:	data_out=16'h89ff;
17'h68d0:	data_out=16'h8965;
17'h68d1:	data_out=16'h89ce;
17'h68d2:	data_out=16'h8a00;
17'h68d3:	data_out=16'h5e1;
17'h68d4:	data_out=16'h89e3;
17'h68d5:	data_out=16'h8821;
17'h68d6:	data_out=16'h9b8;
17'h68d7:	data_out=16'h8894;
17'h68d8:	data_out=16'h837;
17'h68d9:	data_out=16'h8966;
17'h68da:	data_out=16'h898e;
17'h68db:	data_out=16'h533;
17'h68dc:	data_out=16'h9e5;
17'h68dd:	data_out=16'h831d;
17'h68de:	data_out=16'h830b;
17'h68df:	data_out=16'h8a00;
17'h68e0:	data_out=16'h524;
17'h68e1:	data_out=16'h89cb;
17'h68e2:	data_out=16'h80b6;
17'h68e3:	data_out=16'h89d8;
17'h68e4:	data_out=16'h298;
17'h68e5:	data_out=16'h840b;
17'h68e6:	data_out=16'h9c6;
17'h68e7:	data_out=16'ha00;
17'h68e8:	data_out=16'h9fd;
17'h68e9:	data_out=16'h81e;
17'h68ea:	data_out=16'h9fd;
17'h68eb:	data_out=16'h8959;
17'h68ec:	data_out=16'h372;
17'h68ed:	data_out=16'h89d2;
17'h68ee:	data_out=16'h9fd;
17'h68ef:	data_out=16'h89d2;
17'h68f0:	data_out=16'h9fd;
17'h68f1:	data_out=16'h89ff;
17'h68f2:	data_out=16'h8983;
17'h68f3:	data_out=16'h89b3;
17'h68f4:	data_out=16'h4;
17'h68f5:	data_out=16'h837c;
17'h68f6:	data_out=16'h9cc;
17'h68f7:	data_out=16'h8752;
17'h68f8:	data_out=16'h9fb;
17'h68f9:	data_out=16'h9f2;
17'h68fa:	data_out=16'h8836;
17'h68fb:	data_out=16'h9fd;
17'h68fc:	data_out=16'h8a00;
17'h68fd:	data_out=16'h89a6;
17'h68fe:	data_out=16'h351;
17'h68ff:	data_out=16'h89b2;
17'h6900:	data_out=16'h9b8;
17'h6901:	data_out=16'h844a;
17'h6902:	data_out=16'h4a4;
17'h6903:	data_out=16'h96a;
17'h6904:	data_out=16'h9de;
17'h6905:	data_out=16'h87b3;
17'h6906:	data_out=16'h8a00;
17'h6907:	data_out=16'h8a00;
17'h6908:	data_out=16'h9bf;
17'h6909:	data_out=16'h89fc;
17'h690a:	data_out=16'h8726;
17'h690b:	data_out=16'ha00;
17'h690c:	data_out=16'h89ff;
17'h690d:	data_out=16'h8a00;
17'h690e:	data_out=16'h9fb;
17'h690f:	data_out=16'h8a00;
17'h6910:	data_out=16'h9fe;
17'h6911:	data_out=16'h9fc;
17'h6912:	data_out=16'h8a00;
17'h6913:	data_out=16'h89b3;
17'h6914:	data_out=16'h41f;
17'h6915:	data_out=16'h1aa;
17'h6916:	data_out=16'h89e8;
17'h6917:	data_out=16'h80b4;
17'h6918:	data_out=16'h8a00;
17'h6919:	data_out=16'ha00;
17'h691a:	data_out=16'h85fe;
17'h691b:	data_out=16'ha00;
17'h691c:	data_out=16'h9f6;
17'h691d:	data_out=16'h88d;
17'h691e:	data_out=16'h87df;
17'h691f:	data_out=16'h89bf;
17'h6920:	data_out=16'h861c;
17'h6921:	data_out=16'h9fb;
17'h6922:	data_out=16'h9ee;
17'h6923:	data_out=16'h89fb;
17'h6924:	data_out=16'h89fa;
17'h6925:	data_out=16'h8966;
17'h6926:	data_out=16'h9b6;
17'h6927:	data_out=16'h9d4;
17'h6928:	data_out=16'h9fb;
17'h6929:	data_out=16'ha00;
17'h692a:	data_out=16'h8951;
17'h692b:	data_out=16'h90d;
17'h692c:	data_out=16'h89d6;
17'h692d:	data_out=16'h8037;
17'h692e:	data_out=16'h89ca;
17'h692f:	data_out=16'h806b;
17'h6930:	data_out=16'h31e;
17'h6931:	data_out=16'h9e1;
17'h6932:	data_out=16'h8812;
17'h6933:	data_out=16'h8652;
17'h6934:	data_out=16'h89c8;
17'h6935:	data_out=16'h9f2;
17'h6936:	data_out=16'h9b6;
17'h6937:	data_out=16'h9b3;
17'h6938:	data_out=16'h8a00;
17'h6939:	data_out=16'h87a7;
17'h693a:	data_out=16'h89e6;
17'h693b:	data_out=16'h87a8;
17'h693c:	data_out=16'h9ff;
17'h693d:	data_out=16'h9bb;
17'h693e:	data_out=16'h9fb;
17'h693f:	data_out=16'h87bd;
17'h6940:	data_out=16'h865c;
17'h6941:	data_out=16'ha00;
17'h6942:	data_out=16'h9d5;
17'h6943:	data_out=16'ha00;
17'h6944:	data_out=16'h9c8;
17'h6945:	data_out=16'h294;
17'h6946:	data_out=16'ha00;
17'h6947:	data_out=16'h8a00;
17'h6948:	data_out=16'h8a00;
17'h6949:	data_out=16'h22b;
17'h694a:	data_out=16'h869e;
17'h694b:	data_out=16'h98c;
17'h694c:	data_out=16'h8a00;
17'h694d:	data_out=16'h9e4;
17'h694e:	data_out=16'h81ac;
17'h694f:	data_out=16'h8a00;
17'h6950:	data_out=16'h8982;
17'h6951:	data_out=16'h887b;
17'h6952:	data_out=16'h8a00;
17'h6953:	data_out=16'h9d1;
17'h6954:	data_out=16'h8888;
17'h6955:	data_out=16'h9da;
17'h6956:	data_out=16'h9d1;
17'h6957:	data_out=16'h88ff;
17'h6958:	data_out=16'h9da;
17'h6959:	data_out=16'h8920;
17'h695a:	data_out=16'h9c3;
17'h695b:	data_out=16'h9d5;
17'h695c:	data_out=16'h9fa;
17'h695d:	data_out=16'h833c;
17'h695e:	data_out=16'hd1;
17'h695f:	data_out=16'h8a00;
17'h6960:	data_out=16'h935;
17'h6961:	data_out=16'h615;
17'h6962:	data_out=16'h9f6;
17'h6963:	data_out=16'h8706;
17'h6964:	data_out=16'h8a6;
17'h6965:	data_out=16'h9b0;
17'h6966:	data_out=16'h9f5;
17'h6967:	data_out=16'h9e7;
17'h6968:	data_out=16'h9fb;
17'h6969:	data_out=16'h959;
17'h696a:	data_out=16'h9fb;
17'h696b:	data_out=16'h8861;
17'h696c:	data_out=16'h84d5;
17'h696d:	data_out=16'h86dc;
17'h696e:	data_out=16'h9fb;
17'h696f:	data_out=16'h89ff;
17'h6970:	data_out=16'h9fb;
17'h6971:	data_out=16'h8a00;
17'h6972:	data_out=16'h895c;
17'h6973:	data_out=16'h895e;
17'h6974:	data_out=16'heb;
17'h6975:	data_out=16'h9e4;
17'h6976:	data_out=16'h9d9;
17'h6977:	data_out=16'h5b7;
17'h6978:	data_out=16'h9ff;
17'h6979:	data_out=16'h9c6;
17'h697a:	data_out=16'h8361;
17'h697b:	data_out=16'h9fb;
17'h697c:	data_out=16'h8a00;
17'h697d:	data_out=16'h89c2;
17'h697e:	data_out=16'h9fc;
17'h697f:	data_out=16'h89dc;
17'h6980:	data_out=16'h994;
17'h6981:	data_out=16'h876b;
17'h6982:	data_out=16'h80;
17'h6983:	data_out=16'h9af;
17'h6984:	data_out=16'h8b2;
17'h6985:	data_out=16'h89c0;
17'h6986:	data_out=16'h8a00;
17'h6987:	data_out=16'h8a00;
17'h6988:	data_out=16'h9ee;
17'h6989:	data_out=16'h89e1;
17'h698a:	data_out=16'h87c;
17'h698b:	data_out=16'ha00;
17'h698c:	data_out=16'h89ff;
17'h698d:	data_out=16'h8a00;
17'h698e:	data_out=16'h9fe;
17'h698f:	data_out=16'h89ff;
17'h6990:	data_out=16'ha00;
17'h6991:	data_out=16'h9ff;
17'h6992:	data_out=16'h8a00;
17'h6993:	data_out=16'h89d7;
17'h6994:	data_out=16'h433;
17'h6995:	data_out=16'h89e3;
17'h6996:	data_out=16'h8a00;
17'h6997:	data_out=16'h8e7;
17'h6998:	data_out=16'h8a00;
17'h6999:	data_out=16'ha00;
17'h699a:	data_out=16'h89a4;
17'h699b:	data_out=16'ha00;
17'h699c:	data_out=16'h9fc;
17'h699d:	data_out=16'h944;
17'h699e:	data_out=16'h88cb;
17'h699f:	data_out=16'h89fe;
17'h69a0:	data_out=16'h8950;
17'h69a1:	data_out=16'h9fe;
17'h69a2:	data_out=16'h9fd;
17'h69a3:	data_out=16'h8a00;
17'h69a4:	data_out=16'h89ff;
17'h69a5:	data_out=16'h897e;
17'h69a6:	data_out=16'h9b6;
17'h69a7:	data_out=16'h9be;
17'h69a8:	data_out=16'h9ff;
17'h69a9:	data_out=16'ha00;
17'h69aa:	data_out=16'h8985;
17'h69ab:	data_out=16'h9d4;
17'h69ac:	data_out=16'h8a00;
17'h69ad:	data_out=16'h94e;
17'h69ae:	data_out=16'h8926;
17'h69af:	data_out=16'h847f;
17'h69b0:	data_out=16'h81b4;
17'h69b1:	data_out=16'h1b1;
17'h69b2:	data_out=16'h89e6;
17'h69b3:	data_out=16'h85e2;
17'h69b4:	data_out=16'h89f0;
17'h69b5:	data_out=16'h9e1;
17'h69b6:	data_out=16'h9ca;
17'h69b7:	data_out=16'h938;
17'h69b8:	data_out=16'h8886;
17'h69b9:	data_out=16'h8708;
17'h69ba:	data_out=16'h89f6;
17'h69bb:	data_out=16'h89f3;
17'h69bc:	data_out=16'ha00;
17'h69bd:	data_out=16'h6bd;
17'h69be:	data_out=16'h9ff;
17'h69bf:	data_out=16'h89bf;
17'h69c0:	data_out=16'h89c2;
17'h69c1:	data_out=16'ha00;
17'h69c2:	data_out=16'h9b7;
17'h69c3:	data_out=16'ha00;
17'h69c4:	data_out=16'h8e1;
17'h69c5:	data_out=16'h89e5;
17'h69c6:	data_out=16'ha00;
17'h69c7:	data_out=16'h8a00;
17'h69c8:	data_out=16'h8a00;
17'h69c9:	data_out=16'ha6;
17'h69ca:	data_out=16'h89d6;
17'h69cb:	data_out=16'h985;
17'h69cc:	data_out=16'h8a00;
17'h69cd:	data_out=16'h9f0;
17'h69ce:	data_out=16'h877c;
17'h69cf:	data_out=16'h89ff;
17'h69d0:	data_out=16'h89e1;
17'h69d1:	data_out=16'h8a00;
17'h69d2:	data_out=16'h89ff;
17'h69d3:	data_out=16'h9e6;
17'h69d4:	data_out=16'h8966;
17'h69d5:	data_out=16'h863;
17'h69d6:	data_out=16'h9d9;
17'h69d7:	data_out=16'h8957;
17'h69d8:	data_out=16'h9f9;
17'h69d9:	data_out=16'h89bb;
17'h69da:	data_out=16'h9fa;
17'h69db:	data_out=16'h7b;
17'h69dc:	data_out=16'h9e7;
17'h69dd:	data_out=16'h8598;
17'h69de:	data_out=16'h8233;
17'h69df:	data_out=16'h8a00;
17'h69e0:	data_out=16'h95a;
17'h69e1:	data_out=16'h8835;
17'h69e2:	data_out=16'h9f7;
17'h69e3:	data_out=16'h8696;
17'h69e4:	data_out=16'h96d;
17'h69e5:	data_out=16'h89c2;
17'h69e6:	data_out=16'h9f6;
17'h69e7:	data_out=16'h108;
17'h69e8:	data_out=16'h9ff;
17'h69e9:	data_out=16'h9a6;
17'h69ea:	data_out=16'h9fe;
17'h69eb:	data_out=16'h8991;
17'h69ec:	data_out=16'h89b2;
17'h69ed:	data_out=16'h8675;
17'h69ee:	data_out=16'h9fe;
17'h69ef:	data_out=16'h8a00;
17'h69f0:	data_out=16'h9fe;
17'h69f1:	data_out=16'h8a00;
17'h69f2:	data_out=16'h89b6;
17'h69f3:	data_out=16'h89bc;
17'h69f4:	data_out=16'h8368;
17'h69f5:	data_out=16'h9e3;
17'h69f6:	data_out=16'h9e9;
17'h69f7:	data_out=16'h394;
17'h69f8:	data_out=16'ha00;
17'h69f9:	data_out=16'h9c1;
17'h69fa:	data_out=16'h830e;
17'h69fb:	data_out=16'h9ff;
17'h69fc:	data_out=16'h8a00;
17'h69fd:	data_out=16'h89fa;
17'h69fe:	data_out=16'h9fe;
17'h69ff:	data_out=16'h8a00;
17'h6a00:	data_out=16'h992;
17'h6a01:	data_out=16'h29b;
17'h6a02:	data_out=16'hd6;
17'h6a03:	data_out=16'h9bd;
17'h6a04:	data_out=16'h85e5;
17'h6a05:	data_out=16'h8a00;
17'h6a06:	data_out=16'h8a00;
17'h6a07:	data_out=16'h8a00;
17'h6a08:	data_out=16'h9e9;
17'h6a09:	data_out=16'h89cb;
17'h6a0a:	data_out=16'h9ae;
17'h6a0b:	data_out=16'ha00;
17'h6a0c:	data_out=16'h844f;
17'h6a0d:	data_out=16'h8a00;
17'h6a0e:	data_out=16'ha00;
17'h6a0f:	data_out=16'h89ac;
17'h6a10:	data_out=16'h9e4;
17'h6a11:	data_out=16'ha00;
17'h6a12:	data_out=16'h8a00;
17'h6a13:	data_out=16'h89ed;
17'h6a14:	data_out=16'h81fc;
17'h6a15:	data_out=16'h89f9;
17'h6a16:	data_out=16'h8a00;
17'h6a17:	data_out=16'h835a;
17'h6a18:	data_out=16'h8a00;
17'h6a19:	data_out=16'ha00;
17'h6a1a:	data_out=16'h8a00;
17'h6a1b:	data_out=16'ha00;
17'h6a1c:	data_out=16'h9fc;
17'h6a1d:	data_out=16'h9b6;
17'h6a1e:	data_out=16'h87f7;
17'h6a1f:	data_out=16'h89cc;
17'h6a20:	data_out=16'h892e;
17'h6a21:	data_out=16'ha00;
17'h6a22:	data_out=16'h9ee;
17'h6a23:	data_out=16'h89fa;
17'h6a24:	data_out=16'h89fa;
17'h6a25:	data_out=16'h87b1;
17'h6a26:	data_out=16'h9c0;
17'h6a27:	data_out=16'h9a6;
17'h6a28:	data_out=16'ha00;
17'h6a29:	data_out=16'h9ec;
17'h6a2a:	data_out=16'h864c;
17'h6a2b:	data_out=16'h9f0;
17'h6a2c:	data_out=16'h8a00;
17'h6a2d:	data_out=16'h9b3;
17'h6a2e:	data_out=16'h84ae;
17'h6a2f:	data_out=16'h85d6;
17'h6a30:	data_out=16'h88c0;
17'h6a31:	data_out=16'h49a;
17'h6a32:	data_out=16'h8a00;
17'h6a33:	data_out=16'h870b;
17'h6a34:	data_out=16'h8559;
17'h6a35:	data_out=16'h9c4;
17'h6a36:	data_out=16'h9c1;
17'h6a37:	data_out=16'h9ce;
17'h6a38:	data_out=16'h837f;
17'h6a39:	data_out=16'h87a8;
17'h6a3a:	data_out=16'h89e7;
17'h6a3b:	data_out=16'h89ab;
17'h6a3c:	data_out=16'h9de;
17'h6a3d:	data_out=16'h7a3;
17'h6a3e:	data_out=16'ha00;
17'h6a3f:	data_out=16'h8a00;
17'h6a40:	data_out=16'h8a00;
17'h6a41:	data_out=16'ha00;
17'h6a42:	data_out=16'h93d;
17'h6a43:	data_out=16'ha00;
17'h6a44:	data_out=16'h59d;
17'h6a45:	data_out=16'h89fd;
17'h6a46:	data_out=16'h9d3;
17'h6a47:	data_out=16'h8a00;
17'h6a48:	data_out=16'h8a00;
17'h6a49:	data_out=16'h289;
17'h6a4a:	data_out=16'h89eb;
17'h6a4b:	data_out=16'h921;
17'h6a4c:	data_out=16'h89ff;
17'h6a4d:	data_out=16'h6fc;
17'h6a4e:	data_out=16'h8572;
17'h6a4f:	data_out=16'h89f9;
17'h6a50:	data_out=16'h8a00;
17'h6a51:	data_out=16'h89f6;
17'h6a52:	data_out=16'h89e5;
17'h6a53:	data_out=16'h5f4;
17'h6a54:	data_out=16'h8964;
17'h6a55:	data_out=16'h7bf;
17'h6a56:	data_out=16'h9df;
17'h6a57:	data_out=16'h8131;
17'h6a58:	data_out=16'h9fd;
17'h6a59:	data_out=16'h8a00;
17'h6a5a:	data_out=16'h9fa;
17'h6a5b:	data_out=16'h4ca;
17'h6a5c:	data_out=16'h5ef;
17'h6a5d:	data_out=16'h845c;
17'h6a5e:	data_out=16'h83a9;
17'h6a5f:	data_out=16'h89ff;
17'h6a60:	data_out=16'h995;
17'h6a61:	data_out=16'h89b0;
17'h6a62:	data_out=16'h9ff;
17'h6a63:	data_out=16'h881f;
17'h6a64:	data_out=16'h9aa;
17'h6a65:	data_out=16'h89fd;
17'h6a66:	data_out=16'h9e7;
17'h6a67:	data_out=16'h89b6;
17'h6a68:	data_out=16'ha00;
17'h6a69:	data_out=16'h9d4;
17'h6a6a:	data_out=16'ha00;
17'h6a6b:	data_out=16'h89ff;
17'h6a6c:	data_out=16'h83ee;
17'h6a6d:	data_out=16'h87d6;
17'h6a6e:	data_out=16'ha00;
17'h6a6f:	data_out=16'h8a00;
17'h6a70:	data_out=16'ha00;
17'h6a71:	data_out=16'h8a00;
17'h6a72:	data_out=16'h8a00;
17'h6a73:	data_out=16'h8a00;
17'h6a74:	data_out=16'h8a00;
17'h6a75:	data_out=16'h952;
17'h6a76:	data_out=16'h9f7;
17'h6a77:	data_out=16'h402;
17'h6a78:	data_out=16'h9fe;
17'h6a79:	data_out=16'h8b9;
17'h6a7a:	data_out=16'h84e2;
17'h6a7b:	data_out=16'ha00;
17'h6a7c:	data_out=16'h8a00;
17'h6a7d:	data_out=16'h89dc;
17'h6a7e:	data_out=16'ha00;
17'h6a7f:	data_out=16'h8a00;
17'h6a80:	data_out=16'h973;
17'h6a81:	data_out=16'h9d2;
17'h6a82:	data_out=16'h9d2;
17'h6a83:	data_out=16'h76d;
17'h6a84:	data_out=16'h855c;
17'h6a85:	data_out=16'h89fe;
17'h6a86:	data_out=16'h8a00;
17'h6a87:	data_out=16'h8a00;
17'h6a88:	data_out=16'h9ef;
17'h6a89:	data_out=16'h8839;
17'h6a8a:	data_out=16'h9c6;
17'h6a8b:	data_out=16'ha00;
17'h6a8c:	data_out=16'h90d;
17'h6a8d:	data_out=16'h8a00;
17'h6a8e:	data_out=16'ha00;
17'h6a8f:	data_out=16'h81f1;
17'h6a90:	data_out=16'h930;
17'h6a91:	data_out=16'ha00;
17'h6a92:	data_out=16'h81b2;
17'h6a93:	data_out=16'h89d8;
17'h6a94:	data_out=16'h830a;
17'h6a95:	data_out=16'h8955;
17'h6a96:	data_out=16'h8922;
17'h6a97:	data_out=16'h8399;
17'h6a98:	data_out=16'h8a00;
17'h6a99:	data_out=16'h9d7;
17'h6a9a:	data_out=16'h89fe;
17'h6a9b:	data_out=16'ha00;
17'h6a9c:	data_out=16'h9fd;
17'h6a9d:	data_out=16'h9bd;
17'h6a9e:	data_out=16'h83db;
17'h6a9f:	data_out=16'h89d6;
17'h6aa0:	data_out=16'h856b;
17'h6aa1:	data_out=16'h9ff;
17'h6aa2:	data_out=16'h83a0;
17'h6aa3:	data_out=16'h46f;
17'h6aa4:	data_out=16'h466;
17'h6aa5:	data_out=16'h8561;
17'h6aa6:	data_out=16'h9e9;
17'h6aa7:	data_out=16'h98d;
17'h6aa8:	data_out=16'h9fe;
17'h6aa9:	data_out=16'h9dd;
17'h6aaa:	data_out=16'h9aa;
17'h6aab:	data_out=16'h953;
17'h6aac:	data_out=16'h89e9;
17'h6aad:	data_out=16'h9df;
17'h6aae:	data_out=16'h2d7;
17'h6aaf:	data_out=16'h83b9;
17'h6ab0:	data_out=16'h8a00;
17'h6ab1:	data_out=16'h9b9;
17'h6ab2:	data_out=16'h89fd;
17'h6ab3:	data_out=16'h8838;
17'h6ab4:	data_out=16'h7e2;
17'h6ab5:	data_out=16'h9ad;
17'h6ab6:	data_out=16'h9e0;
17'h6ab7:	data_out=16'h9ed;
17'h6ab8:	data_out=16'h8156;
17'h6ab9:	data_out=16'h88cd;
17'h6aba:	data_out=16'h87cf;
17'h6abb:	data_out=16'h97c;
17'h6abc:	data_out=16'h9f9;
17'h6abd:	data_out=16'h70d;
17'h6abe:	data_out=16'h9fe;
17'h6abf:	data_out=16'h89fe;
17'h6ac0:	data_out=16'h89fa;
17'h6ac1:	data_out=16'h9fa;
17'h6ac2:	data_out=16'h968;
17'h6ac3:	data_out=16'ha00;
17'h6ac4:	data_out=16'h934;
17'h6ac5:	data_out=16'h8967;
17'h6ac6:	data_out=16'h8242;
17'h6ac7:	data_out=16'h807c;
17'h6ac8:	data_out=16'h89ff;
17'h6ac9:	data_out=16'h8343;
17'h6aca:	data_out=16'h8953;
17'h6acb:	data_out=16'h95f;
17'h6acc:	data_out=16'h89fe;
17'h6acd:	data_out=16'h8833;
17'h6ace:	data_out=16'h412;
17'h6acf:	data_out=16'h86dd;
17'h6ad0:	data_out=16'h89ff;
17'h6ad1:	data_out=16'h8911;
17'h6ad2:	data_out=16'h8281;
17'h6ad3:	data_out=16'h994;
17'h6ad4:	data_out=16'h8613;
17'h6ad5:	data_out=16'h9fb;
17'h6ad6:	data_out=16'h538;
17'h6ad7:	data_out=16'h18c;
17'h6ad8:	data_out=16'h9b1;
17'h6ad9:	data_out=16'h89fc;
17'h6ada:	data_out=16'h9ee;
17'h6adb:	data_out=16'h8ca;
17'h6adc:	data_out=16'h873b;
17'h6add:	data_out=16'h8129;
17'h6ade:	data_out=16'h8137;
17'h6adf:	data_out=16'h89fe;
17'h6ae0:	data_out=16'h9d7;
17'h6ae1:	data_out=16'h89eb;
17'h6ae2:	data_out=16'ha00;
17'h6ae3:	data_out=16'h88e6;
17'h6ae4:	data_out=16'h8ae;
17'h6ae5:	data_out=16'h89ff;
17'h6ae6:	data_out=16'h9d6;
17'h6ae7:	data_out=16'h89e8;
17'h6ae8:	data_out=16'h9fe;
17'h6ae9:	data_out=16'h9f3;
17'h6aea:	data_out=16'ha00;
17'h6aeb:	data_out=16'h89f4;
17'h6aec:	data_out=16'h46e;
17'h6aed:	data_out=16'h8893;
17'h6aee:	data_out=16'ha00;
17'h6aef:	data_out=16'h8a00;
17'h6af0:	data_out=16'ha00;
17'h6af1:	data_out=16'h89ff;
17'h6af2:	data_out=16'h8a00;
17'h6af3:	data_out=16'h89ff;
17'h6af4:	data_out=16'h8a00;
17'h6af5:	data_out=16'h8897;
17'h6af6:	data_out=16'h9c8;
17'h6af7:	data_out=16'h83ea;
17'h6af8:	data_out=16'h9f2;
17'h6af9:	data_out=16'h24;
17'h6afa:	data_out=16'h8348;
17'h6afb:	data_out=16'h9fe;
17'h6afc:	data_out=16'h8a00;
17'h6afd:	data_out=16'h89fc;
17'h6afe:	data_out=16'ha00;
17'h6aff:	data_out=16'h8a00;
17'h6b00:	data_out=16'h6ab;
17'h6b01:	data_out=16'h9d0;
17'h6b02:	data_out=16'h96d;
17'h6b03:	data_out=16'h284;
17'h6b04:	data_out=16'h841c;
17'h6b05:	data_out=16'h89fc;
17'h6b06:	data_out=16'h8a00;
17'h6b07:	data_out=16'h8a00;
17'h6b08:	data_out=16'h76;
17'h6b09:	data_out=16'h89ef;
17'h6b0a:	data_out=16'h9f8;
17'h6b0b:	data_out=16'ha00;
17'h6b0c:	data_out=16'h89ff;
17'h6b0d:	data_out=16'h8a00;
17'h6b0e:	data_out=16'h9fd;
17'h6b0f:	data_out=16'h30f;
17'h6b10:	data_out=16'h8888;
17'h6b11:	data_out=16'ha00;
17'h6b12:	data_out=16'h5a;
17'h6b13:	data_out=16'h8725;
17'h6b14:	data_out=16'h8290;
17'h6b15:	data_out=16'h894d;
17'h6b16:	data_out=16'h89eb;
17'h6b17:	data_out=16'h8646;
17'h6b18:	data_out=16'h8a00;
17'h6b19:	data_out=16'h31a;
17'h6b1a:	data_out=16'h89f8;
17'h6b1b:	data_out=16'h9fa;
17'h6b1c:	data_out=16'h8ec;
17'h6b1d:	data_out=16'h9f2;
17'h6b1e:	data_out=16'h92;
17'h6b1f:	data_out=16'h89f9;
17'h6b20:	data_out=16'h8232;
17'h6b21:	data_out=16'h9fc;
17'h6b22:	data_out=16'h867e;
17'h6b23:	data_out=16'h9fa;
17'h6b24:	data_out=16'h9f7;
17'h6b25:	data_out=16'h86a8;
17'h6b26:	data_out=16'h9f4;
17'h6b27:	data_out=16'h927;
17'h6b28:	data_out=16'h9fb;
17'h6b29:	data_out=16'h9e8;
17'h6b2a:	data_out=16'h9a9;
17'h6b2b:	data_out=16'h660;
17'h6b2c:	data_out=16'h89e9;
17'h6b2d:	data_out=16'h9f1;
17'h6b2e:	data_out=16'h9e9;
17'h6b2f:	data_out=16'h836d;
17'h6b30:	data_out=16'h8a00;
17'h6b31:	data_out=16'h9db;
17'h6b32:	data_out=16'h89f2;
17'h6b33:	data_out=16'h84c2;
17'h6b34:	data_out=16'h8ba;
17'h6b35:	data_out=16'h39b;
17'h6b36:	data_out=16'h8ee;
17'h6b37:	data_out=16'h9ec;
17'h6b38:	data_out=16'h94a;
17'h6b39:	data_out=16'h8965;
17'h6b3a:	data_out=16'h89e9;
17'h6b3b:	data_out=16'h760;
17'h6b3c:	data_out=16'h9ff;
17'h6b3d:	data_out=16'h279;
17'h6b3e:	data_out=16'h9fb;
17'h6b3f:	data_out=16'h89fc;
17'h6b40:	data_out=16'h89ee;
17'h6b41:	data_out=16'h8c4;
17'h6b42:	data_out=16'h871b;
17'h6b43:	data_out=16'ha00;
17'h6b44:	data_out=16'h977;
17'h6b45:	data_out=16'h895f;
17'h6b46:	data_out=16'h9e1;
17'h6b47:	data_out=16'h89e7;
17'h6b48:	data_out=16'h89fd;
17'h6b49:	data_out=16'h8468;
17'h6b4a:	data_out=16'h89ff;
17'h6b4b:	data_out=16'h64;
17'h6b4c:	data_out=16'h89f7;
17'h6b4d:	data_out=16'h8974;
17'h6b4e:	data_out=16'h10d;
17'h6b4f:	data_out=16'h8831;
17'h6b50:	data_out=16'h89f9;
17'h6b51:	data_out=16'h8498;
17'h6b52:	data_out=16'h217;
17'h6b53:	data_out=16'h528;
17'h6b54:	data_out=16'h83b7;
17'h6b55:	data_out=16'h9e5;
17'h6b56:	data_out=16'h8024;
17'h6b57:	data_out=16'h9c8;
17'h6b58:	data_out=16'h8473;
17'h6b59:	data_out=16'h899f;
17'h6b5a:	data_out=16'h8e7;
17'h6b5b:	data_out=16'h9ce;
17'h6b5c:	data_out=16'h8d7;
17'h6b5d:	data_out=16'h828f;
17'h6b5e:	data_out=16'h8063;
17'h6b5f:	data_out=16'h89ff;
17'h6b60:	data_out=16'h9e1;
17'h6b61:	data_out=16'h832a;
17'h6b62:	data_out=16'ha00;
17'h6b63:	data_out=16'h83cc;
17'h6b64:	data_out=16'h90b;
17'h6b65:	data_out=16'h8a00;
17'h6b66:	data_out=16'h9c5;
17'h6b67:	data_out=16'h89cc;
17'h6b68:	data_out=16'h9fb;
17'h6b69:	data_out=16'h240;
17'h6b6a:	data_out=16'h9fe;
17'h6b6b:	data_out=16'h89f4;
17'h6b6c:	data_out=16'had;
17'h6b6d:	data_out=16'h8351;
17'h6b6e:	data_out=16'h9fe;
17'h6b6f:	data_out=16'h8a00;
17'h6b70:	data_out=16'h9fe;
17'h6b71:	data_out=16'h89ff;
17'h6b72:	data_out=16'h89e7;
17'h6b73:	data_out=16'h8911;
17'h6b74:	data_out=16'h8a00;
17'h6b75:	data_out=16'h976;
17'h6b76:	data_out=16'h9df;
17'h6b77:	data_out=16'h895e;
17'h6b78:	data_out=16'h9cd;
17'h6b79:	data_out=16'h8a00;
17'h6b7a:	data_out=16'h8000;
17'h6b7b:	data_out=16'h9fb;
17'h6b7c:	data_out=16'h8a00;
17'h6b7d:	data_out=16'h89fc;
17'h6b7e:	data_out=16'ha00;
17'h6b7f:	data_out=16'h8a00;
17'h6b80:	data_out=16'h82b8;
17'h6b81:	data_out=16'h9c6;
17'h6b82:	data_out=16'h830;
17'h6b83:	data_out=16'h85e0;
17'h6b84:	data_out=16'h83c1;
17'h6b85:	data_out=16'h89f6;
17'h6b86:	data_out=16'h8a00;
17'h6b87:	data_out=16'h8a00;
17'h6b88:	data_out=16'h85c2;
17'h6b89:	data_out=16'h89f0;
17'h6b8a:	data_out=16'h9ff;
17'h6b8b:	data_out=16'h9f9;
17'h6b8c:	data_out=16'h89c3;
17'h6b8d:	data_out=16'h8a00;
17'h6b8e:	data_out=16'h9fc;
17'h6b8f:	data_out=16'h8b8;
17'h6b90:	data_out=16'h89b5;
17'h6b91:	data_out=16'ha00;
17'h6b92:	data_out=16'h370;
17'h6b93:	data_out=16'h41c;
17'h6b94:	data_out=16'h82f7;
17'h6b95:	data_out=16'h8962;
17'h6b96:	data_out=16'h89f4;
17'h6b97:	data_out=16'h88af;
17'h6b98:	data_out=16'h8a00;
17'h6b99:	data_out=16'h8982;
17'h6b9a:	data_out=16'h89f5;
17'h6b9b:	data_out=16'h9f3;
17'h6b9c:	data_out=16'h6ee;
17'h6b9d:	data_out=16'h9a5;
17'h6b9e:	data_out=16'h69b;
17'h6b9f:	data_out=16'h89fd;
17'h6ba0:	data_out=16'h8043;
17'h6ba1:	data_out=16'h9fa;
17'h6ba2:	data_out=16'h89ad;
17'h6ba3:	data_out=16'ha00;
17'h6ba4:	data_out=16'ha00;
17'h6ba5:	data_out=16'h8934;
17'h6ba6:	data_out=16'h9f3;
17'h6ba7:	data_out=16'h36d;
17'h6ba8:	data_out=16'h9f9;
17'h6ba9:	data_out=16'h9f6;
17'h6baa:	data_out=16'h96a;
17'h6bab:	data_out=16'h8985;
17'h6bac:	data_out=16'h89f4;
17'h6bad:	data_out=16'h9fd;
17'h6bae:	data_out=16'h445;
17'h6baf:	data_out=16'h869c;
17'h6bb0:	data_out=16'h8a00;
17'h6bb1:	data_out=16'h9f6;
17'h6bb2:	data_out=16'h89f2;
17'h6bb3:	data_out=16'h235;
17'h6bb4:	data_out=16'h525;
17'h6bb5:	data_out=16'h611;
17'h6bb6:	data_out=16'h19c;
17'h6bb7:	data_out=16'h9eb;
17'h6bb8:	data_out=16'h578;
17'h6bb9:	data_out=16'h84a0;
17'h6bba:	data_out=16'h89ef;
17'h6bbb:	data_out=16'h194;
17'h6bbc:	data_out=16'ha00;
17'h6bbd:	data_out=16'h8098;
17'h6bbe:	data_out=16'h9f9;
17'h6bbf:	data_out=16'h89f6;
17'h6bc0:	data_out=16'h88d1;
17'h6bc1:	data_out=16'h8990;
17'h6bc2:	data_out=16'h89c6;
17'h6bc3:	data_out=16'ha00;
17'h6bc4:	data_out=16'h9aa;
17'h6bc5:	data_out=16'h8971;
17'h6bc6:	data_out=16'h9ec;
17'h6bc7:	data_out=16'h89ad;
17'h6bc8:	data_out=16'h89fb;
17'h6bc9:	data_out=16'h87eb;
17'h6bca:	data_out=16'h8a00;
17'h6bcb:	data_out=16'h89b3;
17'h6bcc:	data_out=16'h89e3;
17'h6bcd:	data_out=16'h89b9;
17'h6bce:	data_out=16'h8131;
17'h6bcf:	data_out=16'h89d3;
17'h6bd0:	data_out=16'h89f3;
17'h6bd1:	data_out=16'h721;
17'h6bd2:	data_out=16'h8303;
17'h6bd3:	data_out=16'h409;
17'h6bd4:	data_out=16'h85df;
17'h6bd5:	data_out=16'h9d1;
17'h6bd6:	data_out=16'h8950;
17'h6bd7:	data_out=16'h450;
17'h6bd8:	data_out=16'h875b;
17'h6bd9:	data_out=16'h89b8;
17'h6bda:	data_out=16'h847;
17'h6bdb:	data_out=16'h9d3;
17'h6bdc:	data_out=16'h9d3;
17'h6bdd:	data_out=16'h885e;
17'h6bde:	data_out=16'h841e;
17'h6bdf:	data_out=16'h89fb;
17'h6be0:	data_out=16'h9de;
17'h6be1:	data_out=16'h8f2;
17'h6be2:	data_out=16'h9f9;
17'h6be3:	data_out=16'h3df;
17'h6be4:	data_out=16'h2d8;
17'h6be5:	data_out=16'h8a00;
17'h6be6:	data_out=16'h87b1;
17'h6be7:	data_out=16'h89ad;
17'h6be8:	data_out=16'h9f9;
17'h6be9:	data_out=16'h8848;
17'h6bea:	data_out=16'h9fc;
17'h6beb:	data_out=16'h89ec;
17'h6bec:	data_out=16'h87e5;
17'h6bed:	data_out=16'h3c9;
17'h6bee:	data_out=16'h9fc;
17'h6bef:	data_out=16'h89fe;
17'h6bf0:	data_out=16'h9fc;
17'h6bf1:	data_out=16'h4ce;
17'h6bf2:	data_out=16'h89d9;
17'h6bf3:	data_out=16'h89e9;
17'h6bf4:	data_out=16'h8a00;
17'h6bf5:	data_out=16'h98d;
17'h6bf6:	data_out=16'h363;
17'h6bf7:	data_out=16'h89d0;
17'h6bf8:	data_out=16'h991;
17'h6bf9:	data_out=16'h8a00;
17'h6bfa:	data_out=16'h309;
17'h6bfb:	data_out=16'h9f8;
17'h6bfc:	data_out=16'h8a00;
17'h6bfd:	data_out=16'h89fa;
17'h6bfe:	data_out=16'ha00;
17'h6bff:	data_out=16'h89fd;
17'h6c00:	data_out=16'h81c2;
17'h6c01:	data_out=16'h9db;
17'h6c02:	data_out=16'h849e;
17'h6c03:	data_out=16'h88be;
17'h6c04:	data_out=16'hf1;
17'h6c05:	data_out=16'h89fa;
17'h6c06:	data_out=16'h8a00;
17'h6c07:	data_out=16'h8a00;
17'h6c08:	data_out=16'h8335;
17'h6c09:	data_out=16'h89fc;
17'h6c0a:	data_out=16'h9ff;
17'h6c0b:	data_out=16'h9e8;
17'h6c0c:	data_out=16'h89d6;
17'h6c0d:	data_out=16'h89ff;
17'h6c0e:	data_out=16'h9fc;
17'h6c0f:	data_out=16'h8b9;
17'h6c10:	data_out=16'h89eb;
17'h6c11:	data_out=16'ha00;
17'h6c12:	data_out=16'h750;
17'h6c13:	data_out=16'hfe;
17'h6c14:	data_out=16'h8966;
17'h6c15:	data_out=16'h899d;
17'h6c16:	data_out=16'h89f7;
17'h6c17:	data_out=16'h89d1;
17'h6c18:	data_out=16'h89f4;
17'h6c19:	data_out=16'h8860;
17'h6c1a:	data_out=16'h89fd;
17'h6c1b:	data_out=16'h9f1;
17'h6c1c:	data_out=16'h154;
17'h6c1d:	data_out=16'h7dc;
17'h6c1e:	data_out=16'h80e4;
17'h6c1f:	data_out=16'h8a00;
17'h6c20:	data_out=16'h51;
17'h6c21:	data_out=16'h9fb;
17'h6c22:	data_out=16'h89eb;
17'h6c23:	data_out=16'ha00;
17'h6c24:	data_out=16'ha00;
17'h6c25:	data_out=16'h89d5;
17'h6c26:	data_out=16'h86b1;
17'h6c27:	data_out=16'h9af;
17'h6c28:	data_out=16'h9f8;
17'h6c29:	data_out=16'h927;
17'h6c2a:	data_out=16'h9eb;
17'h6c2b:	data_out=16'h89aa;
17'h6c2c:	data_out=16'h89f6;
17'h6c2d:	data_out=16'ha00;
17'h6c2e:	data_out=16'h8289;
17'h6c2f:	data_out=16'h87d1;
17'h6c30:	data_out=16'h8a00;
17'h6c31:	data_out=16'h9fc;
17'h6c32:	data_out=16'h89f7;
17'h6c33:	data_out=16'h89d0;
17'h6c34:	data_out=16'h6ab;
17'h6c35:	data_out=16'h47e;
17'h6c36:	data_out=16'h280;
17'h6c37:	data_out=16'h9b9;
17'h6c38:	data_out=16'h184;
17'h6c39:	data_out=16'h89c8;
17'h6c3a:	data_out=16'h89f6;
17'h6c3b:	data_out=16'h88ce;
17'h6c3c:	data_out=16'h9fd;
17'h6c3d:	data_out=16'h8457;
17'h6c3e:	data_out=16'h9f8;
17'h6c3f:	data_out=16'h89fa;
17'h6c40:	data_out=16'h8878;
17'h6c41:	data_out=16'h89d9;
17'h6c42:	data_out=16'h89c6;
17'h6c43:	data_out=16'h9db;
17'h6c44:	data_out=16'h9c4;
17'h6c45:	data_out=16'h89a1;
17'h6c46:	data_out=16'h9f6;
17'h6c47:	data_out=16'h89de;
17'h6c48:	data_out=16'h89fe;
17'h6c49:	data_out=16'h899e;
17'h6c4a:	data_out=16'h8933;
17'h6c4b:	data_out=16'h89bd;
17'h6c4c:	data_out=16'h89d7;
17'h6c4d:	data_out=16'h89ec;
17'h6c4e:	data_out=16'h38;
17'h6c4f:	data_out=16'h89e0;
17'h6c50:	data_out=16'h89f9;
17'h6c51:	data_out=16'h84c2;
17'h6c52:	data_out=16'h815b;
17'h6c53:	data_out=16'h594;
17'h6c54:	data_out=16'h81bd;
17'h6c55:	data_out=16'h46a;
17'h6c56:	data_out=16'h891c;
17'h6c57:	data_out=16'h85a4;
17'h6c58:	data_out=16'h893a;
17'h6c59:	data_out=16'h89bf;
17'h6c5a:	data_out=16'h87b;
17'h6c5b:	data_out=16'h9ce;
17'h6c5c:	data_out=16'h9dd;
17'h6c5d:	data_out=16'h8907;
17'h6c5e:	data_out=16'h86d9;
17'h6c5f:	data_out=16'h895e;
17'h6c60:	data_out=16'h5bc;
17'h6c61:	data_out=16'h5bf;
17'h6c62:	data_out=16'h3ba;
17'h6c63:	data_out=16'h8903;
17'h6c64:	data_out=16'h704;
17'h6c65:	data_out=16'h8a00;
17'h6c66:	data_out=16'h89b2;
17'h6c67:	data_out=16'h873a;
17'h6c68:	data_out=16'h9f9;
17'h6c69:	data_out=16'h874f;
17'h6c6a:	data_out=16'h9fd;
17'h6c6b:	data_out=16'h89f3;
17'h6c6c:	data_out=16'h877f;
17'h6c6d:	data_out=16'h88cc;
17'h6c6e:	data_out=16'h9fd;
17'h6c6f:	data_out=16'h89fe;
17'h6c70:	data_out=16'h9fd;
17'h6c71:	data_out=16'h65e;
17'h6c72:	data_out=16'h89ed;
17'h6c73:	data_out=16'h89f1;
17'h6c74:	data_out=16'h8a00;
17'h6c75:	data_out=16'h8083;
17'h6c76:	data_out=16'h87a9;
17'h6c77:	data_out=16'h89f9;
17'h6c78:	data_out=16'h8a00;
17'h6c79:	data_out=16'h89fe;
17'h6c7a:	data_out=16'h88f1;
17'h6c7b:	data_out=16'h9f8;
17'h6c7c:	data_out=16'h899b;
17'h6c7d:	data_out=16'h8a00;
17'h6c7e:	data_out=16'ha00;
17'h6c7f:	data_out=16'h89fe;
17'h6c80:	data_out=16'h8688;
17'h6c81:	data_out=16'h802a;
17'h6c82:	data_out=16'h888f;
17'h6c83:	data_out=16'h89c9;
17'h6c84:	data_out=16'h10;
17'h6c85:	data_out=16'h89fb;
17'h6c86:	data_out=16'h8089;
17'h6c87:	data_out=16'h89f5;
17'h6c88:	data_out=16'h85f1;
17'h6c89:	data_out=16'h89fb;
17'h6c8a:	data_out=16'h516;
17'h6c8b:	data_out=16'h872e;
17'h6c8c:	data_out=16'h89bc;
17'h6c8d:	data_out=16'h89fd;
17'h6c8e:	data_out=16'h9fc;
17'h6c8f:	data_out=16'h614;
17'h6c90:	data_out=16'h89ed;
17'h6c91:	data_out=16'ha00;
17'h6c92:	data_out=16'h9ea;
17'h6c93:	data_out=16'h8018;
17'h6c94:	data_out=16'h899c;
17'h6c95:	data_out=16'h89b1;
17'h6c96:	data_out=16'h89de;
17'h6c97:	data_out=16'h89c3;
17'h6c98:	data_out=16'h9fb;
17'h6c99:	data_out=16'h89e6;
17'h6c9a:	data_out=16'h89fe;
17'h6c9b:	data_out=16'h881e;
17'h6c9c:	data_out=16'h899c;
17'h6c9d:	data_out=16'h814a;
17'h6c9e:	data_out=16'h889a;
17'h6c9f:	data_out=16'h89ec;
17'h6ca0:	data_out=16'h86f1;
17'h6ca1:	data_out=16'h9fb;
17'h6ca2:	data_out=16'h89fa;
17'h6ca3:	data_out=16'ha00;
17'h6ca4:	data_out=16'ha00;
17'h6ca5:	data_out=16'h89df;
17'h6ca6:	data_out=16'h889f;
17'h6ca7:	data_out=16'h8681;
17'h6ca8:	data_out=16'h9f8;
17'h6ca9:	data_out=16'h80cc;
17'h6caa:	data_out=16'h9f7;
17'h6cab:	data_out=16'h89c2;
17'h6cac:	data_out=16'h89e1;
17'h6cad:	data_out=16'ha00;
17'h6cae:	data_out=16'h853e;
17'h6caf:	data_out=16'h889f;
17'h6cb0:	data_out=16'h8a00;
17'h6cb1:	data_out=16'h9e8;
17'h6cb2:	data_out=16'h89fa;
17'h6cb3:	data_out=16'h89b7;
17'h6cb4:	data_out=16'h8544;
17'h6cb5:	data_out=16'h883f;
17'h6cb6:	data_out=16'h8508;
17'h6cb7:	data_out=16'h88b9;
17'h6cb8:	data_out=16'h2dd;
17'h6cb9:	data_out=16'h8997;
17'h6cba:	data_out=16'h8959;
17'h6cbb:	data_out=16'h89e2;
17'h6cbc:	data_out=16'h890a;
17'h6cbd:	data_out=16'h86b9;
17'h6cbe:	data_out=16'h9f8;
17'h6cbf:	data_out=16'h89fb;
17'h6cc0:	data_out=16'h8988;
17'h6cc1:	data_out=16'h89d4;
17'h6cc2:	data_out=16'h89a2;
17'h6cc3:	data_out=16'h806d;
17'h6cc4:	data_out=16'h87b0;
17'h6cc5:	data_out=16'h89b6;
17'h6cc6:	data_out=16'h8aa;
17'h6cc7:	data_out=16'h8768;
17'h6cc8:	data_out=16'h8871;
17'h6cc9:	data_out=16'h89b3;
17'h6cca:	data_out=16'h888c;
17'h6ccb:	data_out=16'h8929;
17'h6ccc:	data_out=16'h89dd;
17'h6ccd:	data_out=16'h89f6;
17'h6cce:	data_out=16'h820b;
17'h6ccf:	data_out=16'h89d6;
17'h6cd0:	data_out=16'h89f8;
17'h6cd1:	data_out=16'h89bd;
17'h6cd2:	data_out=16'h511;
17'h6cd3:	data_out=16'h88de;
17'h6cd4:	data_out=16'h86b9;
17'h6cd5:	data_out=16'h8869;
17'h6cd6:	data_out=16'h8918;
17'h6cd7:	data_out=16'h8242;
17'h6cd8:	data_out=16'h8984;
17'h6cd9:	data_out=16'h89d4;
17'h6cda:	data_out=16'h896b;
17'h6cdb:	data_out=16'h9dd;
17'h6cdc:	data_out=16'h8ce;
17'h6cdd:	data_out=16'h897a;
17'h6cde:	data_out=16'h882e;
17'h6cdf:	data_out=16'h6a3;
17'h6ce0:	data_out=16'h34a;
17'h6ce1:	data_out=16'h30;
17'h6ce2:	data_out=16'h88d5;
17'h6ce3:	data_out=16'h89b9;
17'h6ce4:	data_out=16'h31f;
17'h6ce5:	data_out=16'h8a00;
17'h6ce6:	data_out=16'h89cf;
17'h6ce7:	data_out=16'hf9;
17'h6ce8:	data_out=16'h9fa;
17'h6ce9:	data_out=16'h86c6;
17'h6cea:	data_out=16'h9fd;
17'h6ceb:	data_out=16'h89f3;
17'h6cec:	data_out=16'h8829;
17'h6ced:	data_out=16'h89b6;
17'h6cee:	data_out=16'h9fd;
17'h6cef:	data_out=16'h89f8;
17'h6cf0:	data_out=16'h9fd;
17'h6cf1:	data_out=16'h9ee;
17'h6cf2:	data_out=16'h89f3;
17'h6cf3:	data_out=16'h89f8;
17'h6cf4:	data_out=16'h8a00;
17'h6cf5:	data_out=16'h89fa;
17'h6cf6:	data_out=16'h88be;
17'h6cf7:	data_out=16'h89f6;
17'h6cf8:	data_out=16'h8a00;
17'h6cf9:	data_out=16'h89b2;
17'h6cfa:	data_out=16'h8977;
17'h6cfb:	data_out=16'h9f8;
17'h6cfc:	data_out=16'h9fb;
17'h6cfd:	data_out=16'h89fd;
17'h6cfe:	data_out=16'h630;
17'h6cff:	data_out=16'h89fd;
17'h6d00:	data_out=16'ha00;
17'h6d01:	data_out=16'h9d5;
17'h6d02:	data_out=16'h867;
17'h6d03:	data_out=16'h89de;
17'h6d04:	data_out=16'h9f5;
17'h6d05:	data_out=16'h8818;
17'h6d06:	data_out=16'h836;
17'h6d07:	data_out=16'h89df;
17'h6d08:	data_out=16'h4ca;
17'h6d09:	data_out=16'h89fb;
17'h6d0a:	data_out=16'h9e2;
17'h6d0b:	data_out=16'h896d;
17'h6d0c:	data_out=16'h89da;
17'h6d0d:	data_out=16'h89f3;
17'h6d0e:	data_out=16'ha00;
17'h6d0f:	data_out=16'h9fd;
17'h6d10:	data_out=16'h89f9;
17'h6d11:	data_out=16'ha00;
17'h6d12:	data_out=16'h9fb;
17'h6d13:	data_out=16'h64;
17'h6d14:	data_out=16'h8992;
17'h6d15:	data_out=16'h9f7;
17'h6d16:	data_out=16'h822f;
17'h6d17:	data_out=16'h89b7;
17'h6d18:	data_out=16'h9ff;
17'h6d19:	data_out=16'h89fe;
17'h6d1a:	data_out=16'h89fc;
17'h6d1b:	data_out=16'h8972;
17'h6d1c:	data_out=16'h89c0;
17'h6d1d:	data_out=16'h734;
17'h6d1e:	data_out=16'h50e;
17'h6d1f:	data_out=16'h7d0;
17'h6d20:	data_out=16'h8599;
17'h6d21:	data_out=16'h9ff;
17'h6d22:	data_out=16'h89fe;
17'h6d23:	data_out=16'ha00;
17'h6d24:	data_out=16'ha00;
17'h6d25:	data_out=16'h89bd;
17'h6d26:	data_out=16'h73f;
17'h6d27:	data_out=16'h93f;
17'h6d28:	data_out=16'h9fd;
17'h6d29:	data_out=16'h8872;
17'h6d2a:	data_out=16'h9fb;
17'h6d2b:	data_out=16'h89e3;
17'h6d2c:	data_out=16'h53;
17'h6d2d:	data_out=16'ha00;
17'h6d2e:	data_out=16'h9fe;
17'h6d2f:	data_out=16'h8917;
17'h6d30:	data_out=16'h8a00;
17'h6d31:	data_out=16'h9e6;
17'h6d32:	data_out=16'h89fd;
17'h6d33:	data_out=16'h8995;
17'h6d34:	data_out=16'h8217;
17'h6d35:	data_out=16'h9dd;
17'h6d36:	data_out=16'h408;
17'h6d37:	data_out=16'h5bb;
17'h6d38:	data_out=16'h875;
17'h6d39:	data_out=16'h8865;
17'h6d3a:	data_out=16'h306;
17'h6d3b:	data_out=16'h8488;
17'h6d3c:	data_out=16'h89e0;
17'h6d3d:	data_out=16'ha00;
17'h6d3e:	data_out=16'h9fd;
17'h6d3f:	data_out=16'h87c7;
17'h6d40:	data_out=16'h862e;
17'h6d41:	data_out=16'h89e7;
17'h6d42:	data_out=16'h89aa;
17'h6d43:	data_out=16'h898f;
17'h6d44:	data_out=16'h637;
17'h6d45:	data_out=16'h9f7;
17'h6d46:	data_out=16'hc2;
17'h6d47:	data_out=16'h9fa;
17'h6d48:	data_out=16'h862b;
17'h6d49:	data_out=16'h8997;
17'h6d4a:	data_out=16'h803d;
17'h6d4b:	data_out=16'h88ab;
17'h6d4c:	data_out=16'h9e5;
17'h6d4d:	data_out=16'h89fd;
17'h6d4e:	data_out=16'h337;
17'h6d4f:	data_out=16'h9cb;
17'h6d50:	data_out=16'h89fc;
17'h6d51:	data_out=16'h88e1;
17'h6d52:	data_out=16'h9ed;
17'h6d53:	data_out=16'h8978;
17'h6d54:	data_out=16'h8721;
17'h6d55:	data_out=16'h87c0;
17'h6d56:	data_out=16'h9ff;
17'h6d57:	data_out=16'h9fd;
17'h6d58:	data_out=16'h89a5;
17'h6d59:	data_out=16'h9c6;
17'h6d5a:	data_out=16'h89a1;
17'h6d5b:	data_out=16'h9f7;
17'h6d5c:	data_out=16'h8573;
17'h6d5d:	data_out=16'h4c0;
17'h6d5e:	data_out=16'h88d7;
17'h6d5f:	data_out=16'h9ff;
17'h6d60:	data_out=16'h9f7;
17'h6d61:	data_out=16'h8c2;
17'h6d62:	data_out=16'h8974;
17'h6d63:	data_out=16'h898e;
17'h6d64:	data_out=16'h8381;
17'h6d65:	data_out=16'h8a00;
17'h6d66:	data_out=16'h89f0;
17'h6d67:	data_out=16'h8103;
17'h6d68:	data_out=16'h9fe;
17'h6d69:	data_out=16'h26a;
17'h6d6a:	data_out=16'ha00;
17'h6d6b:	data_out=16'h899d;
17'h6d6c:	data_out=16'h9ff;
17'h6d6d:	data_out=16'h8988;
17'h6d6e:	data_out=16'ha00;
17'h6d6f:	data_out=16'h89f9;
17'h6d70:	data_out=16'ha00;
17'h6d71:	data_out=16'h9fe;
17'h6d72:	data_out=16'h618;
17'h6d73:	data_out=16'h822b;
17'h6d74:	data_out=16'h89fe;
17'h6d75:	data_out=16'h89ee;
17'h6d76:	data_out=16'h89c0;
17'h6d77:	data_out=16'h89e4;
17'h6d78:	data_out=16'h8a00;
17'h6d79:	data_out=16'h896b;
17'h6d7a:	data_out=16'h896a;
17'h6d7b:	data_out=16'h9fd;
17'h6d7c:	data_out=16'h9ff;
17'h6d7d:	data_out=16'h8890;
17'h6d7e:	data_out=16'h244;
17'h6d7f:	data_out=16'h8828;
17'h6d80:	data_out=16'ha00;
17'h6d81:	data_out=16'h9ff;
17'h6d82:	data_out=16'ha00;
17'h6d83:	data_out=16'h89c6;
17'h6d84:	data_out=16'ha00;
17'h6d85:	data_out=16'h670;
17'h6d86:	data_out=16'h87b7;
17'h6d87:	data_out=16'h957;
17'h6d88:	data_out=16'h9fc;
17'h6d89:	data_out=16'h8a00;
17'h6d8a:	data_out=16'ha00;
17'h6d8b:	data_out=16'h89d4;
17'h6d8c:	data_out=16'h830a;
17'h6d8d:	data_out=16'h9e1;
17'h6d8e:	data_out=16'ha00;
17'h6d8f:	data_out=16'h9fe;
17'h6d90:	data_out=16'h8a00;
17'h6d91:	data_out=16'h9fc;
17'h6d92:	data_out=16'h9fe;
17'h6d93:	data_out=16'h87;
17'h6d94:	data_out=16'h89df;
17'h6d95:	data_out=16'ha00;
17'h6d96:	data_out=16'h9fe;
17'h6d97:	data_out=16'h89ed;
17'h6d98:	data_out=16'ha00;
17'h6d99:	data_out=16'h8a00;
17'h6d9a:	data_out=16'h8410;
17'h6d9b:	data_out=16'h8989;
17'h6d9c:	data_out=16'h864d;
17'h6d9d:	data_out=16'h6bc;
17'h6d9e:	data_out=16'h7b0;
17'h6d9f:	data_out=16'h3d4;
17'h6da0:	data_out=16'h89b0;
17'h6da1:	data_out=16'ha00;
17'h6da2:	data_out=16'h89f9;
17'h6da3:	data_out=16'ha00;
17'h6da4:	data_out=16'ha00;
17'h6da5:	data_out=16'h808f;
17'h6da6:	data_out=16'ha00;
17'h6da7:	data_out=16'h89bf;
17'h6da8:	data_out=16'ha00;
17'h6da9:	data_out=16'h86ed;
17'h6daa:	data_out=16'h9fd;
17'h6dab:	data_out=16'h8a00;
17'h6dac:	data_out=16'h9fc;
17'h6dad:	data_out=16'ha00;
17'h6dae:	data_out=16'h9fd;
17'h6daf:	data_out=16'h89c8;
17'h6db0:	data_out=16'h8e4;
17'h6db1:	data_out=16'h8d5;
17'h6db2:	data_out=16'h954;
17'h6db3:	data_out=16'h89f6;
17'h6db4:	data_out=16'h816c;
17'h6db5:	data_out=16'h9fd;
17'h6db6:	data_out=16'h9fc;
17'h6db7:	data_out=16'h9ff;
17'h6db8:	data_out=16'h2e3;
17'h6db9:	data_out=16'h89ef;
17'h6dba:	data_out=16'h2cc;
17'h6dbb:	data_out=16'h953;
17'h6dbc:	data_out=16'h89e3;
17'h6dbd:	data_out=16'ha00;
17'h6dbe:	data_out=16'ha00;
17'h6dbf:	data_out=16'h709;
17'h6dc0:	data_out=16'h88e;
17'h6dc1:	data_out=16'h89a6;
17'h6dc2:	data_out=16'h9ff;
17'h6dc3:	data_out=16'h89fd;
17'h6dc4:	data_out=16'h355;
17'h6dc5:	data_out=16'ha00;
17'h6dc6:	data_out=16'h9fe;
17'h6dc7:	data_out=16'h9e4;
17'h6dc8:	data_out=16'h88c0;
17'h6dc9:	data_out=16'h43e;
17'h6dca:	data_out=16'h85cb;
17'h6dcb:	data_out=16'h87e7;
17'h6dcc:	data_out=16'ha00;
17'h6dcd:	data_out=16'h8a00;
17'h6dce:	data_out=16'h968;
17'h6dcf:	data_out=16'h9fd;
17'h6dd0:	data_out=16'h89fe;
17'h6dd1:	data_out=16'h9f9;
17'h6dd2:	data_out=16'ha00;
17'h6dd3:	data_out=16'h89c4;
17'h6dd4:	data_out=16'h899e;
17'h6dd5:	data_out=16'ha00;
17'h6dd6:	data_out=16'ha00;
17'h6dd7:	data_out=16'ha00;
17'h6dd8:	data_out=16'h9e6;
17'h6dd9:	data_out=16'ha00;
17'h6dda:	data_out=16'h89cf;
17'h6ddb:	data_out=16'ha00;
17'h6ddc:	data_out=16'h89ce;
17'h6ddd:	data_out=16'h9c6;
17'h6dde:	data_out=16'h89b9;
17'h6ddf:	data_out=16'h9ff;
17'h6de0:	data_out=16'ha00;
17'h6de1:	data_out=16'ha00;
17'h6de2:	data_out=16'h89be;
17'h6de3:	data_out=16'h89f5;
17'h6de4:	data_out=16'h89ea;
17'h6de5:	data_out=16'h8a00;
17'h6de6:	data_out=16'h8a00;
17'h6de7:	data_out=16'h89d9;
17'h6de8:	data_out=16'ha00;
17'h6de9:	data_out=16'h9fd;
17'h6dea:	data_out=16'ha00;
17'h6deb:	data_out=16'h8754;
17'h6dec:	data_out=16'ha00;
17'h6ded:	data_out=16'h89f3;
17'h6dee:	data_out=16'ha00;
17'h6def:	data_out=16'h89fc;
17'h6df0:	data_out=16'ha00;
17'h6df1:	data_out=16'ha00;
17'h6df2:	data_out=16'h973;
17'h6df3:	data_out=16'h9ee;
17'h6df4:	data_out=16'h9ec;
17'h6df5:	data_out=16'h7c3;
17'h6df6:	data_out=16'h89ee;
17'h6df7:	data_out=16'h840d;
17'h6df8:	data_out=16'h8a00;
17'h6df9:	data_out=16'h9ff;
17'h6dfa:	data_out=16'h89da;
17'h6dfb:	data_out=16'ha00;
17'h6dfc:	data_out=16'ha00;
17'h6dfd:	data_out=16'h89e1;
17'h6dfe:	data_out=16'h841c;
17'h6dff:	data_out=16'h62a;
17'h6e00:	data_out=16'ha00;
17'h6e01:	data_out=16'ha00;
17'h6e02:	data_out=16'ha00;
17'h6e03:	data_out=16'h899d;
17'h6e04:	data_out=16'ha00;
17'h6e05:	data_out=16'ha00;
17'h6e06:	data_out=16'h8a00;
17'h6e07:	data_out=16'h9bd;
17'h6e08:	data_out=16'ha00;
17'h6e09:	data_out=16'h8a00;
17'h6e0a:	data_out=16'ha00;
17'h6e0b:	data_out=16'h8a00;
17'h6e0c:	data_out=16'h2b7;
17'h6e0d:	data_out=16'h9ff;
17'h6e0e:	data_out=16'ha00;
17'h6e0f:	data_out=16'ha00;
17'h6e10:	data_out=16'h8a00;
17'h6e11:	data_out=16'h9a4;
17'h6e12:	data_out=16'ha00;
17'h6e13:	data_out=16'h8286;
17'h6e14:	data_out=16'h8a00;
17'h6e15:	data_out=16'ha00;
17'h6e16:	data_out=16'ha00;
17'h6e17:	data_out=16'h8a00;
17'h6e18:	data_out=16'ha00;
17'h6e19:	data_out=16'h8a00;
17'h6e1a:	data_out=16'ha00;
17'h6e1b:	data_out=16'h8785;
17'h6e1c:	data_out=16'h9f3;
17'h6e1d:	data_out=16'h5e5;
17'h6e1e:	data_out=16'ha00;
17'h6e1f:	data_out=16'h6fd;
17'h6e20:	data_out=16'h976;
17'h6e21:	data_out=16'ha00;
17'h6e22:	data_out=16'h895e;
17'h6e23:	data_out=16'ha00;
17'h6e24:	data_out=16'ha00;
17'h6e25:	data_out=16'ha00;
17'h6e26:	data_out=16'ha00;
17'h6e27:	data_out=16'h51f;
17'h6e28:	data_out=16'ha00;
17'h6e29:	data_out=16'h88c2;
17'h6e2a:	data_out=16'ha00;
17'h6e2b:	data_out=16'h8a00;
17'h6e2c:	data_out=16'ha00;
17'h6e2d:	data_out=16'h89f5;
17'h6e2e:	data_out=16'h9ff;
17'h6e2f:	data_out=16'h8879;
17'h6e30:	data_out=16'ha00;
17'h6e31:	data_out=16'h8701;
17'h6e32:	data_out=16'ha00;
17'h6e33:	data_out=16'h8a00;
17'h6e34:	data_out=16'h89d8;
17'h6e35:	data_out=16'ha00;
17'h6e36:	data_out=16'ha00;
17'h6e37:	data_out=16'ha00;
17'h6e38:	data_out=16'h5b;
17'h6e39:	data_out=16'h87b0;
17'h6e3a:	data_out=16'h22c;
17'h6e3b:	data_out=16'h9ef;
17'h6e3c:	data_out=16'h4a8;
17'h6e3d:	data_out=16'ha00;
17'h6e3e:	data_out=16'ha00;
17'h6e3f:	data_out=16'ha00;
17'h6e40:	data_out=16'ha00;
17'h6e41:	data_out=16'ha00;
17'h6e42:	data_out=16'ha00;
17'h6e43:	data_out=16'h8a00;
17'h6e44:	data_out=16'h804;
17'h6e45:	data_out=16'ha00;
17'h6e46:	data_out=16'ha00;
17'h6e47:	data_out=16'h9c9;
17'h6e48:	data_out=16'h88fa;
17'h6e49:	data_out=16'ha00;
17'h6e4a:	data_out=16'h80db;
17'h6e4b:	data_out=16'h87c7;
17'h6e4c:	data_out=16'ha00;
17'h6e4d:	data_out=16'h89f9;
17'h6e4e:	data_out=16'h9ff;
17'h6e4f:	data_out=16'ha00;
17'h6e50:	data_out=16'h82e6;
17'h6e51:	data_out=16'ha00;
17'h6e52:	data_out=16'ha00;
17'h6e53:	data_out=16'h89ec;
17'h6e54:	data_out=16'h9e8;
17'h6e55:	data_out=16'ha00;
17'h6e56:	data_out=16'ha00;
17'h6e57:	data_out=16'ha00;
17'h6e58:	data_out=16'ha00;
17'h6e59:	data_out=16'ha00;
17'h6e5a:	data_out=16'h8a00;
17'h6e5b:	data_out=16'ha00;
17'h6e5c:	data_out=16'h89e8;
17'h6e5d:	data_out=16'ha00;
17'h6e5e:	data_out=16'h898f;
17'h6e5f:	data_out=16'ha00;
17'h6e60:	data_out=16'ha00;
17'h6e61:	data_out=16'ha00;
17'h6e62:	data_out=16'h89fc;
17'h6e63:	data_out=16'h8a00;
17'h6e64:	data_out=16'h89ff;
17'h6e65:	data_out=16'h8a00;
17'h6e66:	data_out=16'h8a00;
17'h6e67:	data_out=16'h89f1;
17'h6e68:	data_out=16'ha00;
17'h6e69:	data_out=16'h9ff;
17'h6e6a:	data_out=16'ha00;
17'h6e6b:	data_out=16'h9af;
17'h6e6c:	data_out=16'ha00;
17'h6e6d:	data_out=16'h8a00;
17'h6e6e:	data_out=16'ha00;
17'h6e6f:	data_out=16'h755;
17'h6e70:	data_out=16'ha00;
17'h6e71:	data_out=16'ha00;
17'h6e72:	data_out=16'ha00;
17'h6e73:	data_out=16'ha00;
17'h6e74:	data_out=16'ha00;
17'h6e75:	data_out=16'ha00;
17'h6e76:	data_out=16'h8a00;
17'h6e77:	data_out=16'h9fa;
17'h6e78:	data_out=16'h8a00;
17'h6e79:	data_out=16'ha00;
17'h6e7a:	data_out=16'h8a00;
17'h6e7b:	data_out=16'ha00;
17'h6e7c:	data_out=16'ha00;
17'h6e7d:	data_out=16'h87ec;
17'h6e7e:	data_out=16'h87b3;
17'h6e7f:	data_out=16'h9f8;
17'h6e80:	data_out=16'ha00;
17'h6e81:	data_out=16'h9e0;
17'h6e82:	data_out=16'ha00;
17'h6e83:	data_out=16'h931;
17'h6e84:	data_out=16'ha00;
17'h6e85:	data_out=16'ha00;
17'h6e86:	data_out=16'h130;
17'h6e87:	data_out=16'h9f0;
17'h6e88:	data_out=16'ha00;
17'h6e89:	data_out=16'h42e;
17'h6e8a:	data_out=16'ha00;
17'h6e8b:	data_out=16'h8a00;
17'h6e8c:	data_out=16'h6ea;
17'h6e8d:	data_out=16'ha00;
17'h6e8e:	data_out=16'ha00;
17'h6e8f:	data_out=16'ha00;
17'h6e90:	data_out=16'h185;
17'h6e91:	data_out=16'ha00;
17'h6e92:	data_out=16'h82d3;
17'h6e93:	data_out=16'h92c;
17'h6e94:	data_out=16'h61f;
17'h6e95:	data_out=16'ha00;
17'h6e96:	data_out=16'ha00;
17'h6e97:	data_out=16'h8a00;
17'h6e98:	data_out=16'ha00;
17'h6e99:	data_out=16'h8a00;
17'h6e9a:	data_out=16'ha00;
17'h6e9b:	data_out=16'h8118;
17'h6e9c:	data_out=16'ha00;
17'h6e9d:	data_out=16'h693;
17'h6e9e:	data_out=16'h9ff;
17'h6e9f:	data_out=16'h9ed;
17'h6ea0:	data_out=16'ha00;
17'h6ea1:	data_out=16'ha00;
17'h6ea2:	data_out=16'h8914;
17'h6ea3:	data_out=16'ha00;
17'h6ea4:	data_out=16'ha00;
17'h6ea5:	data_out=16'ha00;
17'h6ea6:	data_out=16'ha00;
17'h6ea7:	data_out=16'h9ff;
17'h6ea8:	data_out=16'ha00;
17'h6ea9:	data_out=16'h8a00;
17'h6eaa:	data_out=16'ha00;
17'h6eab:	data_out=16'h8a00;
17'h6eac:	data_out=16'ha00;
17'h6ead:	data_out=16'h8a00;
17'h6eae:	data_out=16'h9ee;
17'h6eaf:	data_out=16'h9f2;
17'h6eb0:	data_out=16'ha00;
17'h6eb1:	data_out=16'h88cb;
17'h6eb2:	data_out=16'ha00;
17'h6eb3:	data_out=16'h726;
17'h6eb4:	data_out=16'h85f7;
17'h6eb5:	data_out=16'ha00;
17'h6eb6:	data_out=16'ha00;
17'h6eb7:	data_out=16'ha00;
17'h6eb8:	data_out=16'h362;
17'h6eb9:	data_out=16'h90b;
17'h6eba:	data_out=16'hc8;
17'h6ebb:	data_out=16'h9ff;
17'h6ebc:	data_out=16'h900;
17'h6ebd:	data_out=16'ha00;
17'h6ebe:	data_out=16'ha00;
17'h6ebf:	data_out=16'ha00;
17'h6ec0:	data_out=16'ha00;
17'h6ec1:	data_out=16'ha00;
17'h6ec2:	data_out=16'h815b;
17'h6ec3:	data_out=16'h8a00;
17'h6ec4:	data_out=16'ha00;
17'h6ec5:	data_out=16'ha00;
17'h6ec6:	data_out=16'h1d2;
17'h6ec7:	data_out=16'h9e3;
17'h6ec8:	data_out=16'h80d1;
17'h6ec9:	data_out=16'ha00;
17'h6eca:	data_out=16'h7d2;
17'h6ecb:	data_out=16'h8965;
17'h6ecc:	data_out=16'ha00;
17'h6ecd:	data_out=16'h8999;
17'h6ece:	data_out=16'ha00;
17'h6ecf:	data_out=16'ha00;
17'h6ed0:	data_out=16'h86d;
17'h6ed1:	data_out=16'ha00;
17'h6ed2:	data_out=16'ha00;
17'h6ed3:	data_out=16'h8506;
17'h6ed4:	data_out=16'ha00;
17'h6ed5:	data_out=16'ha00;
17'h6ed6:	data_out=16'ha00;
17'h6ed7:	data_out=16'ha00;
17'h6ed8:	data_out=16'ha00;
17'h6ed9:	data_out=16'ha00;
17'h6eda:	data_out=16'h8a00;
17'h6edb:	data_out=16'ha00;
17'h6edc:	data_out=16'h480;
17'h6edd:	data_out=16'ha00;
17'h6ede:	data_out=16'h7b4;
17'h6edf:	data_out=16'ha00;
17'h6ee0:	data_out=16'ha00;
17'h6ee1:	data_out=16'ha00;
17'h6ee2:	data_out=16'h8a00;
17'h6ee3:	data_out=16'h5bb;
17'h6ee4:	data_out=16'h89ff;
17'h6ee5:	data_out=16'h8a00;
17'h6ee6:	data_out=16'h8a00;
17'h6ee7:	data_out=16'h8a00;
17'h6ee8:	data_out=16'ha00;
17'h6ee9:	data_out=16'ha00;
17'h6eea:	data_out=16'ha00;
17'h6eeb:	data_out=16'ha00;
17'h6eec:	data_out=16'ha00;
17'h6eed:	data_out=16'h677;
17'h6eee:	data_out=16'ha00;
17'h6eef:	data_out=16'h9f6;
17'h6ef0:	data_out=16'ha00;
17'h6ef1:	data_out=16'ha00;
17'h6ef2:	data_out=16'ha00;
17'h6ef3:	data_out=16'ha00;
17'h6ef4:	data_out=16'ha00;
17'h6ef5:	data_out=16'ha00;
17'h6ef6:	data_out=16'h8a00;
17'h6ef7:	data_out=16'h9fc;
17'h6ef8:	data_out=16'h8a00;
17'h6ef9:	data_out=16'ha00;
17'h6efa:	data_out=16'h878;
17'h6efb:	data_out=16'ha00;
17'h6efc:	data_out=16'ha00;
17'h6efd:	data_out=16'h9f9;
17'h6efe:	data_out=16'h86dc;
17'h6eff:	data_out=16'ha00;
17'h6f00:	data_out=16'hc7;
17'h6f01:	data_out=16'h359;
17'h6f02:	data_out=16'ha00;
17'h6f03:	data_out=16'h4a3;
17'h6f04:	data_out=16'ha00;
17'h6f05:	data_out=16'ha00;
17'h6f06:	data_out=16'h845;
17'h6f07:	data_out=16'h972;
17'h6f08:	data_out=16'ha00;
17'h6f09:	data_out=16'h8424;
17'h6f0a:	data_out=16'h698;
17'h6f0b:	data_out=16'h8a00;
17'h6f0c:	data_out=16'h8df;
17'h6f0d:	data_out=16'h822;
17'h6f0e:	data_out=16'h731;
17'h6f0f:	data_out=16'ha00;
17'h6f10:	data_out=16'h82da;
17'h6f11:	data_out=16'h9cd;
17'h6f12:	data_out=16'h1a5;
17'h6f13:	data_out=16'h5bb;
17'h6f14:	data_out=16'h3ee;
17'h6f15:	data_out=16'ha00;
17'h6f16:	data_out=16'ha00;
17'h6f17:	data_out=16'h8175;
17'h6f18:	data_out=16'ha00;
17'h6f19:	data_out=16'h8a00;
17'h6f1a:	data_out=16'ha00;
17'h6f1b:	data_out=16'h87b7;
17'h6f1c:	data_out=16'h9fd;
17'h6f1d:	data_out=16'h21d;
17'h6f1e:	data_out=16'h766;
17'h6f1f:	data_out=16'h9fa;
17'h6f20:	data_out=16'h5d6;
17'h6f21:	data_out=16'h716;
17'h6f22:	data_out=16'h868a;
17'h6f23:	data_out=16'h90e;
17'h6f24:	data_out=16'h916;
17'h6f25:	data_out=16'h1d8;
17'h6f26:	data_out=16'h830d;
17'h6f27:	data_out=16'h19d;
17'h6f28:	data_out=16'h6f8;
17'h6f29:	data_out=16'h842b;
17'h6f2a:	data_out=16'h90e;
17'h6f2b:	data_out=16'h8a00;
17'h6f2c:	data_out=16'ha00;
17'h6f2d:	data_out=16'h8a00;
17'h6f2e:	data_out=16'h9f1;
17'h6f2f:	data_out=16'h34;
17'h6f30:	data_out=16'ha00;
17'h6f31:	data_out=16'h878f;
17'h6f32:	data_out=16'ha00;
17'h6f33:	data_out=16'h50f;
17'h6f34:	data_out=16'h830f;
17'h6f35:	data_out=16'ha00;
17'h6f36:	data_out=16'ha00;
17'h6f37:	data_out=16'ha00;
17'h6f38:	data_out=16'h96d;
17'h6f39:	data_out=16'h61d;
17'h6f3a:	data_out=16'h17;
17'h6f3b:	data_out=16'h9d7;
17'h6f3c:	data_out=16'h64d;
17'h6f3d:	data_out=16'ha00;
17'h6f3e:	data_out=16'h6f8;
17'h6f3f:	data_out=16'ha00;
17'h6f40:	data_out=16'ha00;
17'h6f41:	data_out=16'ha00;
17'h6f42:	data_out=16'h20b;
17'h6f43:	data_out=16'h522;
17'h6f44:	data_out=16'h9cb;
17'h6f45:	data_out=16'ha00;
17'h6f46:	data_out=16'h86b2;
17'h6f47:	data_out=16'h38b;
17'h6f48:	data_out=16'h19a;
17'h6f49:	data_out=16'h2ab;
17'h6f4a:	data_out=16'h974;
17'h6f4b:	data_out=16'h8594;
17'h6f4c:	data_out=16'h767;
17'h6f4d:	data_out=16'h86cf;
17'h6f4e:	data_out=16'ha00;
17'h6f4f:	data_out=16'h7b9;
17'h6f50:	data_out=16'h9f5;
17'h6f51:	data_out=16'ha00;
17'h6f52:	data_out=16'ha00;
17'h6f53:	data_out=16'h84a5;
17'h6f54:	data_out=16'h709;
17'h6f55:	data_out=16'h9fe;
17'h6f56:	data_out=16'ha00;
17'h6f57:	data_out=16'ha00;
17'h6f58:	data_out=16'ha00;
17'h6f59:	data_out=16'ha00;
17'h6f5a:	data_out=16'h8841;
17'h6f5b:	data_out=16'ha00;
17'h6f5c:	data_out=16'h27e;
17'h6f5d:	data_out=16'ha00;
17'h6f5e:	data_out=16'h80af;
17'h6f5f:	data_out=16'h587;
17'h6f60:	data_out=16'h81e3;
17'h6f61:	data_out=16'ha00;
17'h6f62:	data_out=16'h840c;
17'h6f63:	data_out=16'h494;
17'h6f64:	data_out=16'h88a4;
17'h6f65:	data_out=16'h89bd;
17'h6f66:	data_out=16'h8a00;
17'h6f67:	data_out=16'h841c;
17'h6f68:	data_out=16'h704;
17'h6f69:	data_out=16'h9fc;
17'h6f6a:	data_out=16'h748;
17'h6f6b:	data_out=16'ha00;
17'h6f6c:	data_out=16'h6f0;
17'h6f6d:	data_out=16'h4bf;
17'h6f6e:	data_out=16'h748;
17'h6f6f:	data_out=16'h9fe;
17'h6f70:	data_out=16'h73c;
17'h6f71:	data_out=16'ha00;
17'h6f72:	data_out=16'ha00;
17'h6f73:	data_out=16'ha00;
17'h6f74:	data_out=16'ha00;
17'h6f75:	data_out=16'ha00;
17'h6f76:	data_out=16'h8a00;
17'h6f77:	data_out=16'h9fe;
17'h6f78:	data_out=16'h44b;
17'h6f79:	data_out=16'ha00;
17'h6f7a:	data_out=16'h494;
17'h6f7b:	data_out=16'h6f8;
17'h6f7c:	data_out=16'h855;
17'h6f7d:	data_out=16'ha00;
17'h6f7e:	data_out=16'h85dc;
17'h6f7f:	data_out=16'ha00;
17'h6f80:	data_out=16'h8155;
17'h6f81:	data_out=16'h2d;
17'h6f82:	data_out=16'h40;
17'h6f83:	data_out=16'h1a;
17'h6f84:	data_out=16'h2ef;
17'h6f85:	data_out=16'h165;
17'h6f86:	data_out=16'h1b8;
17'h6f87:	data_out=16'hca;
17'h6f88:	data_out=16'h8177;
17'h6f89:	data_out=16'h80e0;
17'h6f8a:	data_out=16'h9c;
17'h6f8b:	data_out=16'h81d2;
17'h6f8c:	data_out=16'h2d9;
17'h6f8d:	data_out=16'h805c;
17'h6f8e:	data_out=16'h5e;
17'h6f8f:	data_out=16'h802c;
17'h6f90:	data_out=16'h80b5;
17'h6f91:	data_out=16'h157;
17'h6f92:	data_out=16'h8106;
17'h6f93:	data_out=16'h65;
17'h6f94:	data_out=16'h8130;
17'h6f95:	data_out=16'h26;
17'h6f96:	data_out=16'h8006;
17'h6f97:	data_out=16'h8146;
17'h6f98:	data_out=16'h24;
17'h6f99:	data_out=16'hfa;
17'h6f9a:	data_out=16'h28e;
17'h6f9b:	data_out=16'h8135;
17'h6f9c:	data_out=16'h1;
17'h6f9d:	data_out=16'h8116;
17'h6f9e:	data_out=16'h815b;
17'h6f9f:	data_out=16'had;
17'h6fa0:	data_out=16'h813d;
17'h6fa1:	data_out=16'h56;
17'h6fa2:	data_out=16'h805f;
17'h6fa3:	data_out=16'h137;
17'h6fa4:	data_out=16'h137;
17'h6fa5:	data_out=16'h137;
17'h6fa6:	data_out=16'h825b;
17'h6fa7:	data_out=16'h81d5;
17'h6fa8:	data_out=16'h5f;
17'h6fa9:	data_out=16'h8014;
17'h6faa:	data_out=16'h815c;
17'h6fab:	data_out=16'h82b1;
17'h6fac:	data_out=16'h801f;
17'h6fad:	data_out=16'h96;
17'h6fae:	data_out=16'h813d;
17'h6faf:	data_out=16'h802a;
17'h6fb0:	data_out=16'h184;
17'h6fb1:	data_out=16'h8090;
17'h6fb2:	data_out=16'h198;
17'h6fb3:	data_out=16'h817d;
17'h6fb4:	data_out=16'h804e;
17'h6fb5:	data_out=16'h27c;
17'h6fb6:	data_out=16'h8040;
17'h6fb7:	data_out=16'h8002;
17'h6fb8:	data_out=16'h22b;
17'h6fb9:	data_out=16'h811f;
17'h6fba:	data_out=16'h36;
17'h6fbb:	data_out=16'h22;
17'h6fbc:	data_out=16'h80a3;
17'h6fbd:	data_out=16'h807d;
17'h6fbe:	data_out=16'h5d;
17'h6fbf:	data_out=16'h27b;
17'h6fc0:	data_out=16'h30a;
17'h6fc1:	data_out=16'h80e1;
17'h6fc2:	data_out=16'h293;
17'h6fc3:	data_out=16'h1e5;
17'h6fc4:	data_out=16'h4a;
17'h6fc5:	data_out=16'hc;
17'h6fc6:	data_out=16'h81d4;
17'h6fc7:	data_out=16'h80;
17'h6fc8:	data_out=16'h80e1;
17'h6fc9:	data_out=16'h153;
17'h6fca:	data_out=16'h20b;
17'h6fcb:	data_out=16'h2ad;
17'h6fcc:	data_out=16'h1e3;
17'h6fcd:	data_out=16'h8050;
17'h6fce:	data_out=16'h30;
17'h6fcf:	data_out=16'h1cf;
17'h6fd0:	data_out=16'h2ad;
17'h6fd1:	data_out=16'h17;
17'h6fd2:	data_out=16'h148;
17'h6fd3:	data_out=16'h81f7;
17'h6fd4:	data_out=16'h8045;
17'h6fd5:	data_out=16'h804e;
17'h6fd6:	data_out=16'h8043;
17'h6fd7:	data_out=16'h138;
17'h6fd8:	data_out=16'h8082;
17'h6fd9:	data_out=16'h27e;
17'h6fda:	data_out=16'h81a9;
17'h6fdb:	data_out=16'h14f;
17'h6fdc:	data_out=16'hb;
17'h6fdd:	data_out=16'h807e;
17'h6fde:	data_out=16'h8034;
17'h6fdf:	data_out=16'h8034;
17'h6fe0:	data_out=16'h810c;
17'h6fe1:	data_out=16'he6;
17'h6fe2:	data_out=16'h8169;
17'h6fe3:	data_out=16'h8164;
17'h6fe4:	data_out=16'h80f4;
17'h6fe5:	data_out=16'h1cb;
17'h6fe6:	data_out=16'h111;
17'h6fe7:	data_out=16'h8136;
17'h6fe8:	data_out=16'h57;
17'h6fe9:	data_out=16'h8108;
17'h6fea:	data_out=16'h66;
17'h6feb:	data_out=16'h1d8;
17'h6fec:	data_out=16'h803d;
17'h6fed:	data_out=16'h8173;
17'h6fee:	data_out=16'h5d;
17'h6fef:	data_out=16'he0;
17'h6ff0:	data_out=16'h5f;
17'h6ff1:	data_out=16'h8160;
17'h6ff2:	data_out=16'h12f;
17'h6ff3:	data_out=16'h196;
17'h6ff4:	data_out=16'h188;
17'h6ff5:	data_out=16'h161;
17'h6ff6:	data_out=16'h82df;
17'h6ff7:	data_out=16'h2a7;
17'h6ff8:	data_out=16'h149;
17'h6ff9:	data_out=16'h815c;
17'h6ffa:	data_out=16'h813b;
17'h6ffb:	data_out=16'h5c;
17'h6ffc:	data_out=16'h8002;
17'h6ffd:	data_out=16'h1a5;
17'h6ffe:	data_out=16'h80c3;
17'h6fff:	data_out=16'h21f;
17'h7000:	data_out=16'hc7;
17'h7001:	data_out=16'h32;
17'h7002:	data_out=16'h808f;
17'h7003:	data_out=16'h80c6;
17'h7004:	data_out=16'h8016;
17'h7005:	data_out=16'h80ec;
17'h7006:	data_out=16'h80c0;
17'h7007:	data_out=16'h3d;
17'h7008:	data_out=16'h77;
17'h7009:	data_out=16'h4e;
17'h700a:	data_out=16'h115;
17'h700b:	data_out=16'h8015;
17'h700c:	data_out=16'h170;
17'h700d:	data_out=16'h80ba;
17'h700e:	data_out=16'h803d;
17'h700f:	data_out=16'h80e7;
17'h7010:	data_out=16'h8014;
17'h7011:	data_out=16'h78;
17'h7012:	data_out=16'h804c;
17'h7013:	data_out=16'h80a9;
17'h7014:	data_out=16'h8127;
17'h7015:	data_out=16'h803b;
17'h7016:	data_out=16'h805f;
17'h7017:	data_out=16'h8127;
17'h7018:	data_out=16'h802e;
17'h7019:	data_out=16'h169;
17'h701a:	data_out=16'h8033;
17'h701b:	data_out=16'h80ba;
17'h701c:	data_out=16'h810b;
17'h701d:	data_out=16'h74;
17'h701e:	data_out=16'h8125;
17'h701f:	data_out=16'h8112;
17'h7020:	data_out=16'h80bf;
17'h7021:	data_out=16'h8031;
17'h7022:	data_out=16'h8055;
17'h7023:	data_out=16'hdb;
17'h7024:	data_out=16'hd9;
17'h7025:	data_out=16'ha;
17'h7026:	data_out=16'hd4;
17'h7027:	data_out=16'h42;
17'h7028:	data_out=16'h802e;
17'h7029:	data_out=16'h80a8;
17'h702a:	data_out=16'h8040;
17'h702b:	data_out=16'h11a;
17'h702c:	data_out=16'h8050;
17'h702d:	data_out=16'ha1;
17'h702e:	data_out=16'h80f2;
17'h702f:	data_out=16'h80b5;
17'h7030:	data_out=16'h8029;
17'h7031:	data_out=16'h125;
17'h7032:	data_out=16'h802f;
17'h7033:	data_out=16'h8129;
17'h7034:	data_out=16'he8;
17'h7035:	data_out=16'ha3;
17'h7036:	data_out=16'h8040;
17'h7037:	data_out=16'h80b7;
17'h7038:	data_out=16'h8072;
17'h7039:	data_out=16'h80f5;
17'h703a:	data_out=16'h8001;
17'h703b:	data_out=16'h102;
17'h703c:	data_out=16'h807c;
17'h703d:	data_out=16'h8016;
17'h703e:	data_out=16'h803c;
17'h703f:	data_out=16'h80ca;
17'h7040:	data_out=16'h80cf;
17'h7041:	data_out=16'h80bd;
17'h7042:	data_out=16'hbb;
17'h7043:	data_out=16'h811d;
17'h7044:	data_out=16'h3a;
17'h7045:	data_out=16'h8040;
17'h7046:	data_out=16'h8064;
17'h7047:	data_out=16'h802a;
17'h7048:	data_out=16'h80c3;
17'h7049:	data_out=16'h8009;
17'h704a:	data_out=16'h8021;
17'h704b:	data_out=16'h15a;
17'h704c:	data_out=16'h8031;
17'h704d:	data_out=16'h8058;
17'h704e:	data_out=16'h8052;
17'h704f:	data_out=16'h8010;
17'h7050:	data_out=16'h810e;
17'h7051:	data_out=16'h80c9;
17'h7052:	data_out=16'hae;
17'h7053:	data_out=16'h809a;
17'h7054:	data_out=16'h80ba;
17'h7055:	data_out=16'h80a3;
17'h7056:	data_out=16'h80a1;
17'h7057:	data_out=16'h8071;
17'h7058:	data_out=16'h807a;
17'h7059:	data_out=16'h807f;
17'h705a:	data_out=16'h80bf;
17'h705b:	data_out=16'h8091;
17'h705c:	data_out=16'h801a;
17'h705d:	data_out=16'h80a3;
17'h705e:	data_out=16'h80be;
17'h705f:	data_out=16'h8046;
17'h7060:	data_out=16'h88;
17'h7061:	data_out=16'h805f;
17'h7062:	data_out=16'h8088;
17'h7063:	data_out=16'h812c;
17'h7064:	data_out=16'haa;
17'h7065:	data_out=16'h2f;
17'h7066:	data_out=16'h14a;
17'h7067:	data_out=16'h80e5;
17'h7068:	data_out=16'h8030;
17'h7069:	data_out=16'h53;
17'h706a:	data_out=16'h8033;
17'h706b:	data_out=16'h808b;
17'h706c:	data_out=16'hc0;
17'h706d:	data_out=16'h8126;
17'h706e:	data_out=16'h803c;
17'h706f:	data_out=16'h80d7;
17'h7070:	data_out=16'h8034;
17'h7071:	data_out=16'h80ac;
17'h7072:	data_out=16'h80ef;
17'h7073:	data_out=16'h80e5;
17'h7074:	data_out=16'h8022;
17'h7075:	data_out=16'h80cc;
17'h7076:	data_out=16'hb7;
17'h7077:	data_out=16'h807d;
17'h7078:	data_out=16'h80c4;
17'h7079:	data_out=16'h80f6;
17'h707a:	data_out=16'h8135;
17'h707b:	data_out=16'h8032;
17'h707c:	data_out=16'h8067;
17'h707d:	data_out=16'h811a;
17'h707e:	data_out=16'h4d;
17'h707f:	data_out=16'h80b5;
17'h7080:	data_out=16'h3d5;
17'h7081:	data_out=16'h3ce;
17'h7082:	data_out=16'h153;
17'h7083:	data_out=16'h1e3;
17'h7084:	data_out=16'h8035;
17'h7085:	data_out=16'h8063;
17'h7086:	data_out=16'h8231;
17'h7087:	data_out=16'h89;
17'h7088:	data_out=16'h25b;
17'h7089:	data_out=16'had;
17'h708a:	data_out=16'h1cc;
17'h708b:	data_out=16'hf;
17'h708c:	data_out=16'h8068;
17'h708d:	data_out=16'h1ef;
17'h708e:	data_out=16'h8015;
17'h708f:	data_out=16'h1d5;
17'h7090:	data_out=16'h1cb;
17'h7091:	data_out=16'h8059;
17'h7092:	data_out=16'h242;
17'h7093:	data_out=16'h177;
17'h7094:	data_out=16'h1a0;
17'h7095:	data_out=16'hcd;
17'h7096:	data_out=16'h10f;
17'h7097:	data_out=16'h1f3;
17'h7098:	data_out=16'h7a;
17'h7099:	data_out=16'h16;
17'h709a:	data_out=16'h80bd;
17'h709b:	data_out=16'h2af;
17'h709c:	data_out=16'hb;
17'h709d:	data_out=16'h364;
17'h709e:	data_out=16'h280;
17'h709f:	data_out=16'h81db;
17'h70a0:	data_out=16'h575;
17'h70a1:	data_out=16'h8012;
17'h70a2:	data_out=16'h302;
17'h70a3:	data_out=16'h8072;
17'h70a4:	data_out=16'h8070;
17'h70a5:	data_out=16'h197;
17'h70a6:	data_out=16'h8064;
17'h70a7:	data_out=16'h3a3;
17'h70a8:	data_out=16'h8006;
17'h70a9:	data_out=16'h23a;
17'h70aa:	data_out=16'h350;
17'h70ab:	data_out=16'h19c;
17'h70ac:	data_out=16'ha9;
17'h70ad:	data_out=16'h3ed;
17'h70ae:	data_out=16'h28e;
17'h70af:	data_out=16'h53a;
17'h70b0:	data_out=16'h8087;
17'h70b1:	data_out=16'h1d0;
17'h70b2:	data_out=16'h806c;
17'h70b3:	data_out=16'h1e8;
17'h70b4:	data_out=16'h1ac;
17'h70b5:	data_out=16'h80c5;
17'h70b6:	data_out=16'h32f;
17'h70b7:	data_out=16'h14d;
17'h70b8:	data_out=16'h8013;
17'h70b9:	data_out=16'h222;
17'h70ba:	data_out=16'h412;
17'h70bb:	data_out=16'h807a;
17'h70bc:	data_out=16'h280;
17'h70bd:	data_out=16'h169;
17'h70be:	data_out=16'h800a;
17'h70bf:	data_out=16'h808f;
17'h70c0:	data_out=16'h8011;
17'h70c1:	data_out=16'h149;
17'h70c2:	data_out=16'h483;
17'h70c3:	data_out=16'h82d1;
17'h70c4:	data_out=16'h8063;
17'h70c5:	data_out=16'hf;
17'h70c6:	data_out=16'h224;
17'h70c7:	data_out=16'h1e4;
17'h70c8:	data_out=16'h1e0;
17'h70c9:	data_out=16'h14e;
17'h70ca:	data_out=16'h14d;
17'h70cb:	data_out=16'h3d7;
17'h70cc:	data_out=16'h2e5;
17'h70cd:	data_out=16'h345;
17'h70ce:	data_out=16'h332;
17'h70cf:	data_out=16'h23f;
17'h70d0:	data_out=16'h80b6;
17'h70d1:	data_out=16'h8081;
17'h70d2:	data_out=16'h809b;
17'h70d3:	data_out=16'h4ee;
17'h70d4:	data_out=16'h542;
17'h70d5:	data_out=16'hf;
17'h70d6:	data_out=16'h56;
17'h70d7:	data_out=16'h4e;
17'h70d8:	data_out=16'h8d;
17'h70d9:	data_out=16'ha4;
17'h70da:	data_out=16'h1c2;
17'h70db:	data_out=16'h81d4;
17'h70dc:	data_out=16'h1dc;
17'h70dd:	data_out=16'h3d3;
17'h70de:	data_out=16'h50a;
17'h70df:	data_out=16'h274;
17'h70e0:	data_out=16'ha4;
17'h70e1:	data_out=16'h80ac;
17'h70e2:	data_out=16'h7d;
17'h70e3:	data_out=16'h1e6;
17'h70e4:	data_out=16'hb3;
17'h70e5:	data_out=16'hd2;
17'h70e6:	data_out=16'h8067;
17'h70e7:	data_out=16'h1e6;
17'h70e8:	data_out=16'h8015;
17'h70e9:	data_out=16'h1fd;
17'h70ea:	data_out=16'h8011;
17'h70eb:	data_out=16'h8038;
17'h70ec:	data_out=16'h6fc;
17'h70ed:	data_out=16'h1f2;
17'h70ee:	data_out=16'h8019;
17'h70ef:	data_out=16'he1;
17'h70f0:	data_out=16'h800e;
17'h70f1:	data_out=16'h55;
17'h70f2:	data_out=16'h80bc;
17'h70f3:	data_out=16'h8052;
17'h70f4:	data_out=16'h808b;
17'h70f5:	data_out=16'h820e;
17'h70f6:	data_out=16'h10f;
17'h70f7:	data_out=16'h80f1;
17'h70f8:	data_out=16'h8238;
17'h70f9:	data_out=16'h2b2;
17'h70fa:	data_out=16'h1cf;
17'h70fb:	data_out=16'h800d;
17'h70fc:	data_out=16'h8a;
17'h70fd:	data_out=16'h82c1;
17'h70fe:	data_out=16'h805a;
17'h70ff:	data_out=16'h80aa;
17'h7100:	data_out=16'h9dc;
17'h7101:	data_out=16'ha00;
17'h7102:	data_out=16'h40c;
17'h7103:	data_out=16'h83e;
17'h7104:	data_out=16'h2a5;
17'h7105:	data_out=16'h1fd;
17'h7106:	data_out=16'h8338;
17'h7107:	data_out=16'h81d;
17'h7108:	data_out=16'h49a;
17'h7109:	data_out=16'h6cf;
17'h710a:	data_out=16'h7a7;
17'h710b:	data_out=16'h805c;
17'h710c:	data_out=16'h83e6;
17'h710d:	data_out=16'h576;
17'h710e:	data_out=16'h6e;
17'h710f:	data_out=16'h779;
17'h7110:	data_out=16'h820;
17'h7111:	data_out=16'h5b;
17'h7112:	data_out=16'h9aa;
17'h7113:	data_out=16'h81f;
17'h7114:	data_out=16'h491;
17'h7115:	data_out=16'h1df;
17'h7116:	data_out=16'h4b8;
17'h7117:	data_out=16'h51b;
17'h7118:	data_out=16'h9a;
17'h7119:	data_out=16'hc9;
17'h711a:	data_out=16'h164;
17'h711b:	data_out=16'h95e;
17'h711c:	data_out=16'h37;
17'h711d:	data_out=16'ha00;
17'h711e:	data_out=16'h89a;
17'h711f:	data_out=16'h6d;
17'h7120:	data_out=16'ha00;
17'h7121:	data_out=16'h6d;
17'h7122:	data_out=16'ha00;
17'h7123:	data_out=16'h845a;
17'h7124:	data_out=16'h845b;
17'h7125:	data_out=16'h8ad;
17'h7126:	data_out=16'h1bd;
17'h7127:	data_out=16'ha00;
17'h7128:	data_out=16'h6c;
17'h7129:	data_out=16'ha00;
17'h712a:	data_out=16'ha00;
17'h712b:	data_out=16'h4dc;
17'h712c:	data_out=16'h3b2;
17'h712d:	data_out=16'h8ac;
17'h712e:	data_out=16'h879;
17'h712f:	data_out=16'ha00;
17'h7130:	data_out=16'h8042;
17'h7131:	data_out=16'h72e;
17'h7132:	data_out=16'h7d;
17'h7133:	data_out=16'h63d;
17'h7134:	data_out=16'h386;
17'h7135:	data_out=16'h8141;
17'h7136:	data_out=16'h73c;
17'h7137:	data_out=16'h418;
17'h7138:	data_out=16'ha5;
17'h7139:	data_out=16'h6f3;
17'h713a:	data_out=16'ha00;
17'h713b:	data_out=16'h6a;
17'h713c:	data_out=16'h4ae;
17'h713d:	data_out=16'h917;
17'h713e:	data_out=16'h6c;
17'h713f:	data_out=16'h19a;
17'h7140:	data_out=16'h578;
17'h7141:	data_out=16'h8141;
17'h7142:	data_out=16'ha00;
17'h7143:	data_out=16'h857b;
17'h7144:	data_out=16'h2e0;
17'h7145:	data_out=16'h1d9;
17'h7146:	data_out=16'h38f;
17'h7147:	data_out=16'ha00;
17'h7148:	data_out=16'h85a;
17'h7149:	data_out=16'h860;
17'h714a:	data_out=16'h77f;
17'h714b:	data_out=16'h98e;
17'h714c:	data_out=16'ha00;
17'h714d:	data_out=16'ha00;
17'h714e:	data_out=16'h9e9;
17'h714f:	data_out=16'ha00;
17'h7150:	data_out=16'h193;
17'h7151:	data_out=16'h84ec;
17'h7152:	data_out=16'h83e5;
17'h7153:	data_out=16'ha00;
17'h7154:	data_out=16'ha00;
17'h7155:	data_out=16'h8367;
17'h7156:	data_out=16'h70f;
17'h7157:	data_out=16'h7ff;
17'h7158:	data_out=16'h8051;
17'h7159:	data_out=16'h805;
17'h715a:	data_out=16'h5a4;
17'h715b:	data_out=16'h858a;
17'h715c:	data_out=16'h714;
17'h715d:	data_out=16'ha00;
17'h715e:	data_out=16'ha00;
17'h715f:	data_out=16'h732;
17'h7160:	data_out=16'h334;
17'h7161:	data_out=16'h8103;
17'h7162:	data_out=16'h815d;
17'h7163:	data_out=16'h5ef;
17'h7164:	data_out=16'h268;
17'h7165:	data_out=16'h96f;
17'h7166:	data_out=16'h3a;
17'h7167:	data_out=16'h64f;
17'h7168:	data_out=16'h6c;
17'h7169:	data_out=16'h401;
17'h716a:	data_out=16'h6c;
17'h716b:	data_out=16'h315;
17'h716c:	data_out=16'ha00;
17'h716d:	data_out=16'h635;
17'h716e:	data_out=16'h6c;
17'h716f:	data_out=16'h82f;
17'h7170:	data_out=16'h6d;
17'h7171:	data_out=16'h3ca;
17'h7172:	data_out=16'h3c3;
17'h7173:	data_out=16'h4bd;
17'h7174:	data_out=16'h8060;
17'h7175:	data_out=16'h877f;
17'h7176:	data_out=16'h294;
17'h7177:	data_out=16'h1e2;
17'h7178:	data_out=16'h848f;
17'h7179:	data_out=16'h9e0;
17'h717a:	data_out=16'h529;
17'h717b:	data_out=16'h6c;
17'h717c:	data_out=16'h1ea;
17'h717d:	data_out=16'h8411;
17'h717e:	data_out=16'h442;
17'h717f:	data_out=16'h502;
17'h7180:	data_out=16'h840b;
17'h7181:	data_out=16'ha00;
17'h7182:	data_out=16'h9f6;
17'h7183:	data_out=16'h99b;
17'h7184:	data_out=16'h8463;
17'h7185:	data_out=16'h6f3;
17'h7186:	data_out=16'h8221;
17'h7187:	data_out=16'h9fa;
17'h7188:	data_out=16'h33a;
17'h7189:	data_out=16'h888b;
17'h718a:	data_out=16'h4a5;
17'h718b:	data_out=16'ha00;
17'h718c:	data_out=16'h82c2;
17'h718d:	data_out=16'h748;
17'h718e:	data_out=16'h8126;
17'h718f:	data_out=16'h9fe;
17'h7190:	data_out=16'h41e;
17'h7191:	data_out=16'h20f;
17'h7192:	data_out=16'h9ff;
17'h7193:	data_out=16'h7a1;
17'h7194:	data_out=16'h9fd;
17'h7195:	data_out=16'h875d;
17'h7196:	data_out=16'h83ec;
17'h7197:	data_out=16'h9fb;
17'h7198:	data_out=16'h80f7;
17'h7199:	data_out=16'h27c;
17'h719a:	data_out=16'h81ed;
17'h719b:	data_out=16'h9f9;
17'h719c:	data_out=16'h4f3;
17'h719d:	data_out=16'ha00;
17'h719e:	data_out=16'ha00;
17'h719f:	data_out=16'h8736;
17'h71a0:	data_out=16'ha00;
17'h71a1:	data_out=16'h810e;
17'h71a2:	data_out=16'h9e0;
17'h71a3:	data_out=16'h8a00;
17'h71a4:	data_out=16'h8a00;
17'h71a5:	data_out=16'h1dc;
17'h71a6:	data_out=16'h8a00;
17'h71a7:	data_out=16'ha00;
17'h71a8:	data_out=16'h80d4;
17'h71a9:	data_out=16'h9ff;
17'h71aa:	data_out=16'ha00;
17'h71ab:	data_out=16'ha00;
17'h71ac:	data_out=16'h8593;
17'h71ad:	data_out=16'h5ee;
17'h71ae:	data_out=16'ha00;
17'h71af:	data_out=16'ha00;
17'h71b0:	data_out=16'h831b;
17'h71b1:	data_out=16'h9fd;
17'h71b2:	data_out=16'h82aa;
17'h71b3:	data_out=16'ha00;
17'h71b4:	data_out=16'h6ac;
17'h71b5:	data_out=16'h8197;
17'h71b6:	data_out=16'ha00;
17'h71b7:	data_out=16'h9fb;
17'h71b8:	data_out=16'ha00;
17'h71b9:	data_out=16'ha00;
17'h71ba:	data_out=16'h9f1;
17'h71bb:	data_out=16'h8607;
17'h71bc:	data_out=16'h9fb;
17'h71bd:	data_out=16'ha1;
17'h71be:	data_out=16'h80d1;
17'h71bf:	data_out=16'h6c8;
17'h71c0:	data_out=16'h87f6;
17'h71c1:	data_out=16'h385;
17'h71c2:	data_out=16'h935;
17'h71c3:	data_out=16'h8809;
17'h71c4:	data_out=16'ha0;
17'h71c5:	data_out=16'h876e;
17'h71c6:	data_out=16'h9a4;
17'h71c7:	data_out=16'h5d5;
17'h71c8:	data_out=16'ha00;
17'h71c9:	data_out=16'h16;
17'h71ca:	data_out=16'ha00;
17'h71cb:	data_out=16'h9fe;
17'h71cc:	data_out=16'h8fb;
17'h71cd:	data_out=16'h9ff;
17'h71ce:	data_out=16'ha00;
17'h71cf:	data_out=16'h65c;
17'h71d0:	data_out=16'h890d;
17'h71d1:	data_out=16'h8a00;
17'h71d2:	data_out=16'h8a00;
17'h71d3:	data_out=16'ha00;
17'h71d4:	data_out=16'ha00;
17'h71d5:	data_out=16'h8872;
17'h71d6:	data_out=16'h856f;
17'h71d7:	data_out=16'h8435;
17'h71d8:	data_out=16'h825b;
17'h71d9:	data_out=16'h84de;
17'h71da:	data_out=16'h9fc;
17'h71db:	data_out=16'h80ad;
17'h71dc:	data_out=16'h9ff;
17'h71dd:	data_out=16'h9ff;
17'h71de:	data_out=16'ha00;
17'h71df:	data_out=16'ha00;
17'h71e0:	data_out=16'h89fd;
17'h71e1:	data_out=16'h82aa;
17'h71e2:	data_out=16'h9fe;
17'h71e3:	data_out=16'ha00;
17'h71e4:	data_out=16'h3ce;
17'h71e5:	data_out=16'ha00;
17'h71e6:	data_out=16'h303;
17'h71e7:	data_out=16'ha00;
17'h71e8:	data_out=16'h8103;
17'h71e9:	data_out=16'h98;
17'h71ea:	data_out=16'h813d;
17'h71eb:	data_out=16'h137;
17'h71ec:	data_out=16'h9dc;
17'h71ed:	data_out=16'ha00;
17'h71ee:	data_out=16'h813d;
17'h71ef:	data_out=16'h980;
17'h71f0:	data_out=16'h8131;
17'h71f1:	data_out=16'ha00;
17'h71f2:	data_out=16'h848f;
17'h71f3:	data_out=16'h16f;
17'h71f4:	data_out=16'h834d;
17'h71f5:	data_out=16'h872;
17'h71f6:	data_out=16'h603;
17'h71f7:	data_out=16'h8893;
17'h71f8:	data_out=16'h885a;
17'h71f9:	data_out=16'h9fe;
17'h71fa:	data_out=16'ha00;
17'h71fb:	data_out=16'h80d0;
17'h71fc:	data_out=16'h599;
17'h71fd:	data_out=16'h12b;
17'h71fe:	data_out=16'h8996;
17'h71ff:	data_out=16'h89eb;
17'h7200:	data_out=16'h8a00;
17'h7201:	data_out=16'h9f2;
17'h7202:	data_out=16'h90c;
17'h7203:	data_out=16'h89ff;
17'h7204:	data_out=16'h899e;
17'h7205:	data_out=16'h9fc;
17'h7206:	data_out=16'ha00;
17'h7207:	data_out=16'h87a;
17'h7208:	data_out=16'h87cb;
17'h7209:	data_out=16'h8930;
17'h720a:	data_out=16'h8a00;
17'h720b:	data_out=16'h9fb;
17'h720c:	data_out=16'h847c;
17'h720d:	data_out=16'h8390;
17'h720e:	data_out=16'h84fb;
17'h720f:	data_out=16'h9dc;
17'h7210:	data_out=16'h8985;
17'h7211:	data_out=16'h95d;
17'h7212:	data_out=16'h9f1;
17'h7213:	data_out=16'h8630;
17'h7214:	data_out=16'h9f9;
17'h7215:	data_out=16'h8a00;
17'h7216:	data_out=16'h89ff;
17'h7217:	data_out=16'h9f2;
17'h7218:	data_out=16'h86de;
17'h7219:	data_out=16'ha00;
17'h721a:	data_out=16'h518;
17'h721b:	data_out=16'h9c1;
17'h721c:	data_out=16'h666;
17'h721d:	data_out=16'h9fb;
17'h721e:	data_out=16'h9e4;
17'h721f:	data_out=16'h8031;
17'h7220:	data_out=16'h9eb;
17'h7221:	data_out=16'h8411;
17'h7222:	data_out=16'h2a2;
17'h7223:	data_out=16'h8a00;
17'h7224:	data_out=16'h8a00;
17'h7225:	data_out=16'h89f3;
17'h7226:	data_out=16'h8a00;
17'h7227:	data_out=16'h9f8;
17'h7228:	data_out=16'h8293;
17'h7229:	data_out=16'h3bb;
17'h722a:	data_out=16'h8076;
17'h722b:	data_out=16'ha00;
17'h722c:	data_out=16'h89ff;
17'h722d:	data_out=16'h87b2;
17'h722e:	data_out=16'ha00;
17'h722f:	data_out=16'h9f3;
17'h7230:	data_out=16'h862d;
17'h7231:	data_out=16'h9e1;
17'h7232:	data_out=16'h85f8;
17'h7233:	data_out=16'ha00;
17'h7234:	data_out=16'h83ef;
17'h7235:	data_out=16'h533;
17'h7236:	data_out=16'h8097;
17'h7237:	data_out=16'h9d8;
17'h7238:	data_out=16'ha00;
17'h7239:	data_out=16'h9fc;
17'h723a:	data_out=16'h386;
17'h723b:	data_out=16'h89d8;
17'h723c:	data_out=16'h88a;
17'h723d:	data_out=16'h89fe;
17'h723e:	data_out=16'h828a;
17'h723f:	data_out=16'h9fc;
17'h7240:	data_out=16'h884a;
17'h7241:	data_out=16'h530;
17'h7242:	data_out=16'h8a00;
17'h7243:	data_out=16'ha00;
17'h7244:	data_out=16'h86c5;
17'h7245:	data_out=16'h8a00;
17'h7246:	data_out=16'h6e4;
17'h7247:	data_out=16'h8831;
17'h7248:	data_out=16'ha00;
17'h7249:	data_out=16'h89fd;
17'h724a:	data_out=16'ha00;
17'h724b:	data_out=16'h672;
17'h724c:	data_out=16'h8994;
17'h724d:	data_out=16'h640;
17'h724e:	data_out=16'h9fa;
17'h724f:	data_out=16'h89f7;
17'h7250:	data_out=16'h86be;
17'h7251:	data_out=16'h89f8;
17'h7252:	data_out=16'h8a00;
17'h7253:	data_out=16'ha00;
17'h7254:	data_out=16'h9e8;
17'h7255:	data_out=16'h89f0;
17'h7256:	data_out=16'h8a00;
17'h7257:	data_out=16'h89fd;
17'h7258:	data_out=16'h89fa;
17'h7259:	data_out=16'h89da;
17'h725a:	data_out=16'h9f5;
17'h725b:	data_out=16'h245;
17'h725c:	data_out=16'h9f6;
17'h725d:	data_out=16'h5b4;
17'h725e:	data_out=16'h9f2;
17'h725f:	data_out=16'h9fd;
17'h7260:	data_out=16'h8a00;
17'h7261:	data_out=16'h8701;
17'h7262:	data_out=16'h9e3;
17'h7263:	data_out=16'ha00;
17'h7264:	data_out=16'h379;
17'h7265:	data_out=16'ha00;
17'h7266:	data_out=16'ha00;
17'h7267:	data_out=16'ha00;
17'h7268:	data_out=16'h836b;
17'h7269:	data_out=16'h8a00;
17'h726a:	data_out=16'h864c;
17'h726b:	data_out=16'h601;
17'h726c:	data_out=16'h8a00;
17'h726d:	data_out=16'ha00;
17'h726e:	data_out=16'h864d;
17'h726f:	data_out=16'h4e5;
17'h7270:	data_out=16'h854d;
17'h7271:	data_out=16'h9f2;
17'h7272:	data_out=16'h89e4;
17'h7273:	data_out=16'h8696;
17'h7274:	data_out=16'h86d5;
17'h7275:	data_out=16'h7e7;
17'h7276:	data_out=16'ha00;
17'h7277:	data_out=16'h89f3;
17'h7278:	data_out=16'h9f4;
17'h7279:	data_out=16'h945;
17'h727a:	data_out=16'ha00;
17'h727b:	data_out=16'h8287;
17'h727c:	data_out=16'ha00;
17'h727d:	data_out=16'ha00;
17'h727e:	data_out=16'h89ac;
17'h727f:	data_out=16'h8894;
17'h7280:	data_out=16'h8a00;
17'h7281:	data_out=16'h9eb;
17'h7282:	data_out=16'h96c;
17'h7283:	data_out=16'h8a00;
17'h7284:	data_out=16'h85;
17'h7285:	data_out=16'h9f4;
17'h7286:	data_out=16'h8313;
17'h7287:	data_out=16'h95e;
17'h7288:	data_out=16'h8067;
17'h7289:	data_out=16'h89b4;
17'h728a:	data_out=16'h8a00;
17'h728b:	data_out=16'h9f5;
17'h728c:	data_out=16'h89e5;
17'h728d:	data_out=16'h8992;
17'h728e:	data_out=16'h80a8;
17'h728f:	data_out=16'h9fa;
17'h7290:	data_out=16'h8929;
17'h7291:	data_out=16'h9e9;
17'h7292:	data_out=16'ha00;
17'h7293:	data_out=16'h89f7;
17'h7294:	data_out=16'h887;
17'h7295:	data_out=16'h89ff;
17'h7296:	data_out=16'h89fc;
17'h7297:	data_out=16'h823;
17'h7298:	data_out=16'h733;
17'h7299:	data_out=16'h9fc;
17'h729a:	data_out=16'h9f9;
17'h729b:	data_out=16'h810;
17'h729c:	data_out=16'h46;
17'h729d:	data_out=16'h9e7;
17'h729e:	data_out=16'h9b2;
17'h729f:	data_out=16'h829a;
17'h72a0:	data_out=16'h9e6;
17'h72a1:	data_out=16'hc;
17'h72a2:	data_out=16'ha00;
17'h72a3:	data_out=16'h8a00;
17'h72a4:	data_out=16'h8a00;
17'h72a5:	data_out=16'h89ec;
17'h72a6:	data_out=16'h8a00;
17'h72a7:	data_out=16'h9f8;
17'h72a8:	data_out=16'h12b;
17'h72a9:	data_out=16'h80c6;
17'h72aa:	data_out=16'h9e2;
17'h72ab:	data_out=16'ha00;
17'h72ac:	data_out=16'h89fd;
17'h72ad:	data_out=16'h843c;
17'h72ae:	data_out=16'ha00;
17'h72af:	data_out=16'h9f2;
17'h72b0:	data_out=16'h825f;
17'h72b1:	data_out=16'h5a1;
17'h72b2:	data_out=16'h80da;
17'h72b3:	data_out=16'ha00;
17'h72b4:	data_out=16'h82db;
17'h72b5:	data_out=16'h67c;
17'h72b6:	data_out=16'h9f9;
17'h72b7:	data_out=16'h9ea;
17'h72b8:	data_out=16'h9ee;
17'h72b9:	data_out=16'ha00;
17'h72ba:	data_out=16'h8bd;
17'h72bb:	data_out=16'h8942;
17'h72bc:	data_out=16'h559;
17'h72bd:	data_out=16'h82d9;
17'h72be:	data_out=16'h132;
17'h72bf:	data_out=16'h9f3;
17'h72c0:	data_out=16'h82c2;
17'h72c1:	data_out=16'h58b;
17'h72c2:	data_out=16'h8a00;
17'h72c3:	data_out=16'h870c;
17'h72c4:	data_out=16'h84a8;
17'h72c5:	data_out=16'h89ff;
17'h72c6:	data_out=16'h6bf;
17'h72c7:	data_out=16'h8401;
17'h72c8:	data_out=16'ha00;
17'h72c9:	data_out=16'h89f9;
17'h72ca:	data_out=16'ha00;
17'h72cb:	data_out=16'h6;
17'h72cc:	data_out=16'h8672;
17'h72cd:	data_out=16'ha00;
17'h72ce:	data_out=16'ha00;
17'h72cf:	data_out=16'h8899;
17'h72d0:	data_out=16'h3e1;
17'h72d1:	data_out=16'h89f2;
17'h72d2:	data_out=16'h8a00;
17'h72d3:	data_out=16'ha00;
17'h72d4:	data_out=16'h9e9;
17'h72d5:	data_out=16'h89ea;
17'h72d6:	data_out=16'h8a00;
17'h72d7:	data_out=16'h89eb;
17'h72d8:	data_out=16'h89f0;
17'h72d9:	data_out=16'h879b;
17'h72da:	data_out=16'ha00;
17'h72db:	data_out=16'h7e4;
17'h72dc:	data_out=16'h9f1;
17'h72dd:	data_out=16'h951;
17'h72de:	data_out=16'h9d7;
17'h72df:	data_out=16'ha00;
17'h72e0:	data_out=16'h8a00;
17'h72e1:	data_out=16'h63;
17'h72e2:	data_out=16'h8ef;
17'h72e3:	data_out=16'ha00;
17'h72e4:	data_out=16'h112;
17'h72e5:	data_out=16'h9ef;
17'h72e6:	data_out=16'ha00;
17'h72e7:	data_out=16'h9ff;
17'h72e8:	data_out=16'h85;
17'h72e9:	data_out=16'h89f9;
17'h72ea:	data_out=16'h8143;
17'h72eb:	data_out=16'h872;
17'h72ec:	data_out=16'h8a00;
17'h72ed:	data_out=16'ha00;
17'h72ee:	data_out=16'h8140;
17'h72ef:	data_out=16'h801b;
17'h72f0:	data_out=16'h80e8;
17'h72f1:	data_out=16'ha00;
17'h72f2:	data_out=16'h886f;
17'h72f3:	data_out=16'h84b9;
17'h72f4:	data_out=16'h834a;
17'h72f5:	data_out=16'h3b6;
17'h72f6:	data_out=16'ha00;
17'h72f7:	data_out=16'h8943;
17'h72f8:	data_out=16'hc1;
17'h72f9:	data_out=16'ha00;
17'h72fa:	data_out=16'ha00;
17'h72fb:	data_out=16'h136;
17'h72fc:	data_out=16'ha00;
17'h72fd:	data_out=16'ha00;
17'h72fe:	data_out=16'h89cb;
17'h72ff:	data_out=16'h1da;
17'h7300:	data_out=16'h88b4;
17'h7301:	data_out=16'h9df;
17'h7302:	data_out=16'h9ee;
17'h7303:	data_out=16'h89ff;
17'h7304:	data_out=16'h4f5;
17'h7305:	data_out=16'h810c;
17'h7306:	data_out=16'h891e;
17'h7307:	data_out=16'h116;
17'h7308:	data_out=16'h9ef;
17'h7309:	data_out=16'h89eb;
17'h730a:	data_out=16'h8a00;
17'h730b:	data_out=16'h8790;
17'h730c:	data_out=16'h89d0;
17'h730d:	data_out=16'h89ff;
17'h730e:	data_out=16'h9fe;
17'h730f:	data_out=16'h9fe;
17'h7310:	data_out=16'h89ff;
17'h7311:	data_out=16'h9e8;
17'h7312:	data_out=16'h9f3;
17'h7313:	data_out=16'h89ff;
17'h7314:	data_out=16'hb;
17'h7315:	data_out=16'h89ff;
17'h7316:	data_out=16'h89ff;
17'h7317:	data_out=16'h82dc;
17'h7318:	data_out=16'ha00;
17'h7319:	data_out=16'h9f9;
17'h731a:	data_out=16'h9ff;
17'h731b:	data_out=16'h58f;
17'h731c:	data_out=16'h8a00;
17'h731d:	data_out=16'h9d7;
17'h731e:	data_out=16'h72a;
17'h731f:	data_out=16'h879f;
17'h7320:	data_out=16'h9be;
17'h7321:	data_out=16'h9ff;
17'h7322:	data_out=16'ha00;
17'h7323:	data_out=16'h89ff;
17'h7324:	data_out=16'h89ff;
17'h7325:	data_out=16'h89e6;
17'h7326:	data_out=16'h89fd;
17'h7327:	data_out=16'h9cc;
17'h7328:	data_out=16'ha00;
17'h7329:	data_out=16'h963;
17'h732a:	data_out=16'h9db;
17'h732b:	data_out=16'ha00;
17'h732c:	data_out=16'h89ff;
17'h732d:	data_out=16'h9e3;
17'h732e:	data_out=16'ha00;
17'h732f:	data_out=16'h9c4;
17'h7330:	data_out=16'h2a4;
17'h7331:	data_out=16'h81f7;
17'h7332:	data_out=16'h48f;
17'h7333:	data_out=16'h97d;
17'h7334:	data_out=16'h4cb;
17'h7335:	data_out=16'h6b9;
17'h7336:	data_out=16'h9f1;
17'h7337:	data_out=16'ha00;
17'h7338:	data_out=16'h9e5;
17'h7339:	data_out=16'h91b;
17'h733a:	data_out=16'h32;
17'h733b:	data_out=16'h898b;
17'h733c:	data_out=16'h72e;
17'h733d:	data_out=16'h93;
17'h733e:	data_out=16'ha00;
17'h733f:	data_out=16'h813a;
17'h7340:	data_out=16'h8035;
17'h7341:	data_out=16'h89fa;
17'h7342:	data_out=16'h89fd;
17'h7343:	data_out=16'h89ea;
17'h7344:	data_out=16'h859d;
17'h7345:	data_out=16'h89ff;
17'h7346:	data_out=16'h9e7;
17'h7347:	data_out=16'h85ad;
17'h7348:	data_out=16'h9b0;
17'h7349:	data_out=16'h89f3;
17'h734a:	data_out=16'h9fb;
17'h734b:	data_out=16'h87cf;
17'h734c:	data_out=16'h80ae;
17'h734d:	data_out=16'ha00;
17'h734e:	data_out=16'ha00;
17'h734f:	data_out=16'h83e8;
17'h7350:	data_out=16'h2e2;
17'h7351:	data_out=16'h89f3;
17'h7352:	data_out=16'h8a00;
17'h7353:	data_out=16'ha00;
17'h7354:	data_out=16'h9c3;
17'h7355:	data_out=16'h89e9;
17'h7356:	data_out=16'h89fd;
17'h7357:	data_out=16'h89d2;
17'h7358:	data_out=16'h89ef;
17'h7359:	data_out=16'h816e;
17'h735a:	data_out=16'h93f;
17'h735b:	data_out=16'h9ea;
17'h735c:	data_out=16'h9b5;
17'h735d:	data_out=16'h93f;
17'h735e:	data_out=16'h950;
17'h735f:	data_out=16'h9fd;
17'h7360:	data_out=16'h89fc;
17'h7361:	data_out=16'h175;
17'h7362:	data_out=16'h8227;
17'h7363:	data_out=16'h9f0;
17'h7364:	data_out=16'h60;
17'h7365:	data_out=16'h84d0;
17'h7366:	data_out=16'h9fa;
17'h7367:	data_out=16'ha00;
17'h7368:	data_out=16'ha00;
17'h7369:	data_out=16'h80ae;
17'h736a:	data_out=16'h9f2;
17'h736b:	data_out=16'h8418;
17'h736c:	data_out=16'h847;
17'h736d:	data_out=16'h9ef;
17'h736e:	data_out=16'h9f2;
17'h736f:	data_out=16'h85a7;
17'h7370:	data_out=16'h9f9;
17'h7371:	data_out=16'ha00;
17'h7372:	data_out=16'h834f;
17'h7373:	data_out=16'h4c9;
17'h7374:	data_out=16'h1a2;
17'h7375:	data_out=16'h8580;
17'h7376:	data_out=16'ha00;
17'h7377:	data_out=16'h89f3;
17'h7378:	data_out=16'h1be;
17'h7379:	data_out=16'ha00;
17'h737a:	data_out=16'h6ed;
17'h737b:	data_out=16'ha00;
17'h737c:	data_out=16'ha00;
17'h737d:	data_out=16'h82ec;
17'h737e:	data_out=16'h89d7;
17'h737f:	data_out=16'h908;
17'h7380:	data_out=16'h8e;
17'h7381:	data_out=16'h9e3;
17'h7382:	data_out=16'h947;
17'h7383:	data_out=16'h89fe;
17'h7384:	data_out=16'h917;
17'h7385:	data_out=16'h89e4;
17'h7386:	data_out=16'h89f0;
17'h7387:	data_out=16'h8886;
17'h7388:	data_out=16'h9c9;
17'h7389:	data_out=16'h89f7;
17'h738a:	data_out=16'h89ea;
17'h738b:	data_out=16'h88a9;
17'h738c:	data_out=16'h88e2;
17'h738d:	data_out=16'h8a00;
17'h738e:	data_out=16'h9fc;
17'h738f:	data_out=16'h9ec;
17'h7390:	data_out=16'h89fb;
17'h7391:	data_out=16'h808d;
17'h7392:	data_out=16'h995;
17'h7393:	data_out=16'h8a00;
17'h7394:	data_out=16'h89fd;
17'h7395:	data_out=16'h89fe;
17'h7396:	data_out=16'h89ff;
17'h7397:	data_out=16'h89fc;
17'h7398:	data_out=16'h408;
17'h7399:	data_out=16'h9fe;
17'h739a:	data_out=16'h7e7;
17'h739b:	data_out=16'h89fa;
17'h739c:	data_out=16'h89ff;
17'h739d:	data_out=16'h147;
17'h739e:	data_out=16'h89f4;
17'h739f:	data_out=16'h89ba;
17'h73a0:	data_out=16'h96b;
17'h73a1:	data_out=16'h9ff;
17'h73a2:	data_out=16'ha00;
17'h73a3:	data_out=16'h89fc;
17'h73a4:	data_out=16'h89fd;
17'h73a5:	data_out=16'h89e3;
17'h73a6:	data_out=16'h89e3;
17'h73a7:	data_out=16'h20e;
17'h73a8:	data_out=16'h9ff;
17'h73a9:	data_out=16'h181;
17'h73aa:	data_out=16'h9cb;
17'h73ab:	data_out=16'ha00;
17'h73ac:	data_out=16'h89ff;
17'h73ad:	data_out=16'h9fc;
17'h73ae:	data_out=16'h9ec;
17'h73af:	data_out=16'h84d;
17'h73b0:	data_out=16'h18a;
17'h73b1:	data_out=16'h89fc;
17'h73b2:	data_out=16'h86;
17'h73b3:	data_out=16'h89f7;
17'h73b4:	data_out=16'h9d9;
17'h73b5:	data_out=16'h82b4;
17'h73b6:	data_out=16'h9d2;
17'h73b7:	data_out=16'h938;
17'h73b8:	data_out=16'h9b0;
17'h73b9:	data_out=16'h89f7;
17'h73ba:	data_out=16'h86cd;
17'h73bb:	data_out=16'h89f7;
17'h73bc:	data_out=16'h89f5;
17'h73bd:	data_out=16'h82aa;
17'h73be:	data_out=16'h9ff;
17'h73bf:	data_out=16'h89e5;
17'h73c0:	data_out=16'h8275;
17'h73c1:	data_out=16'h89f9;
17'h73c2:	data_out=16'h89fc;
17'h73c3:	data_out=16'h8944;
17'h73c4:	data_out=16'h8926;
17'h73c5:	data_out=16'h89fe;
17'h73c6:	data_out=16'ha00;
17'h73c7:	data_out=16'h80ef;
17'h73c8:	data_out=16'h1d7;
17'h73c9:	data_out=16'h89f0;
17'h73ca:	data_out=16'h9d2;
17'h73cb:	data_out=16'h89fd;
17'h73cc:	data_out=16'h10e;
17'h73cd:	data_out=16'h9f6;
17'h73ce:	data_out=16'ha00;
17'h73cf:	data_out=16'h81c4;
17'h73d0:	data_out=16'h89fd;
17'h73d1:	data_out=16'h8a00;
17'h73d2:	data_out=16'h89e7;
17'h73d3:	data_out=16'h9cd;
17'h73d4:	data_out=16'h987;
17'h73d5:	data_out=16'h89ff;
17'h73d6:	data_out=16'h8a00;
17'h73d7:	data_out=16'h89cb;
17'h73d8:	data_out=16'h89ff;
17'h73d9:	data_out=16'h8183;
17'h73da:	data_out=16'h89f6;
17'h73db:	data_out=16'h1c9;
17'h73dc:	data_out=16'h1ce;
17'h73dd:	data_out=16'h861;
17'h73de:	data_out=16'h6d3;
17'h73df:	data_out=16'h9fc;
17'h73e0:	data_out=16'h89d1;
17'h73e1:	data_out=16'h80b2;
17'h73e2:	data_out=16'h89fa;
17'h73e3:	data_out=16'h89f6;
17'h73e4:	data_out=16'h84cf;
17'h73e5:	data_out=16'h8936;
17'h73e6:	data_out=16'h9f7;
17'h73e7:	data_out=16'ha00;
17'h73e8:	data_out=16'h9ff;
17'h73e9:	data_out=16'h80af;
17'h73ea:	data_out=16'h9fb;
17'h73eb:	data_out=16'h89ed;
17'h73ec:	data_out=16'h99f;
17'h73ed:	data_out=16'h89f6;
17'h73ee:	data_out=16'h9fb;
17'h73ef:	data_out=16'h898f;
17'h73f0:	data_out=16'h9fc;
17'h73f1:	data_out=16'h9f8;
17'h73f2:	data_out=16'h89ec;
17'h73f3:	data_out=16'h81af;
17'h73f4:	data_out=16'h11;
17'h73f5:	data_out=16'h8a00;
17'h73f6:	data_out=16'ha00;
17'h73f7:	data_out=16'h89f2;
17'h73f8:	data_out=16'h64b;
17'h73f9:	data_out=16'ha00;
17'h73fa:	data_out=16'h89fa;
17'h73fb:	data_out=16'h9ff;
17'h73fc:	data_out=16'ha00;
17'h73fd:	data_out=16'h88c4;
17'h73fe:	data_out=16'h89e5;
17'h73ff:	data_out=16'h3c0;
17'h7400:	data_out=16'h9a6;
17'h7401:	data_out=16'h580;
17'h7402:	data_out=16'h958;
17'h7403:	data_out=16'h89d6;
17'h7404:	data_out=16'h429;
17'h7405:	data_out=16'h89f4;
17'h7406:	data_out=16'h89ff;
17'h7407:	data_out=16'h89ff;
17'h7408:	data_out=16'h9a3;
17'h7409:	data_out=16'h89ed;
17'h740a:	data_out=16'h8a00;
17'h740b:	data_out=16'h86f8;
17'h740c:	data_out=16'h8928;
17'h740d:	data_out=16'h8a00;
17'h740e:	data_out=16'h9ff;
17'h740f:	data_out=16'h9cb;
17'h7410:	data_out=16'h89d6;
17'h7411:	data_out=16'h8978;
17'h7412:	data_out=16'h873;
17'h7413:	data_out=16'h89e3;
17'h7414:	data_out=16'h89e3;
17'h7415:	data_out=16'h89f0;
17'h7416:	data_out=16'h89e8;
17'h7417:	data_out=16'h89e5;
17'h7418:	data_out=16'h9e7;
17'h7419:	data_out=16'h9ff;
17'h741a:	data_out=16'h84ca;
17'h741b:	data_out=16'h89ee;
17'h741c:	data_out=16'h89ed;
17'h741d:	data_out=16'h88e4;
17'h741e:	data_out=16'h89dc;
17'h741f:	data_out=16'h89de;
17'h7420:	data_out=16'h964;
17'h7421:	data_out=16'h9ff;
17'h7422:	data_out=16'ha00;
17'h7423:	data_out=16'h89f7;
17'h7424:	data_out=16'h89f7;
17'h7425:	data_out=16'h89b6;
17'h7426:	data_out=16'h266;
17'h7427:	data_out=16'h8349;
17'h7428:	data_out=16'h9ff;
17'h7429:	data_out=16'h215;
17'h742a:	data_out=16'h9d1;
17'h742b:	data_out=16'ha00;
17'h742c:	data_out=16'h89eb;
17'h742d:	data_out=16'ha00;
17'h742e:	data_out=16'h3e8;
17'h742f:	data_out=16'h68;
17'h7430:	data_out=16'h21b;
17'h7431:	data_out=16'h89f8;
17'h7432:	data_out=16'h86b9;
17'h7433:	data_out=16'h89e6;
17'h7434:	data_out=16'h80f4;
17'h7435:	data_out=16'h83df;
17'h7436:	data_out=16'h9c0;
17'h7437:	data_out=16'h7fd;
17'h7438:	data_out=16'h89f6;
17'h7439:	data_out=16'h89df;
17'h743a:	data_out=16'h8752;
17'h743b:	data_out=16'h89f1;
17'h743c:	data_out=16'h89db;
17'h743d:	data_out=16'h302;
17'h743e:	data_out=16'h9ff;
17'h743f:	data_out=16'h89f4;
17'h7440:	data_out=16'h85ad;
17'h7441:	data_out=16'h89eb;
17'h7442:	data_out=16'h89ef;
17'h7443:	data_out=16'h4fa;
17'h7444:	data_out=16'h89bb;
17'h7445:	data_out=16'h89f1;
17'h7446:	data_out=16'ha00;
17'h7447:	data_out=16'ha00;
17'h7448:	data_out=16'h89fc;
17'h7449:	data_out=16'h89bb;
17'h744a:	data_out=16'h9b5;
17'h744b:	data_out=16'h89fc;
17'h744c:	data_out=16'h846b;
17'h744d:	data_out=16'ha00;
17'h744e:	data_out=16'h9fe;
17'h744f:	data_out=16'h879a;
17'h7450:	data_out=16'h89f4;
17'h7451:	data_out=16'h89f7;
17'h7452:	data_out=16'h89d7;
17'h7453:	data_out=16'h954;
17'h7454:	data_out=16'h95c;
17'h7455:	data_out=16'h89e2;
17'h7456:	data_out=16'h8181;
17'h7457:	data_out=16'h8992;
17'h7458:	data_out=16'h89ff;
17'h7459:	data_out=16'h82d0;
17'h745a:	data_out=16'h89f7;
17'h745b:	data_out=16'h893a;
17'h745c:	data_out=16'h89fc;
17'h745d:	data_out=16'h90b;
17'h745e:	data_out=16'h896d;
17'h745f:	data_out=16'h9f9;
17'h7460:	data_out=16'h892a;
17'h7461:	data_out=16'h871b;
17'h7462:	data_out=16'h89ee;
17'h7463:	data_out=16'h89f2;
17'h7464:	data_out=16'h880a;
17'h7465:	data_out=16'h89c5;
17'h7466:	data_out=16'h9f3;
17'h7467:	data_out=16'ha00;
17'h7468:	data_out=16'h9ff;
17'h7469:	data_out=16'h978;
17'h746a:	data_out=16'h9ff;
17'h746b:	data_out=16'h89eb;
17'h746c:	data_out=16'h9eb;
17'h746d:	data_out=16'h89f2;
17'h746e:	data_out=16'h9ff;
17'h746f:	data_out=16'h89a9;
17'h7470:	data_out=16'h9ff;
17'h7471:	data_out=16'h9c3;
17'h7472:	data_out=16'h89d8;
17'h7473:	data_out=16'h89e2;
17'h7474:	data_out=16'h10a;
17'h7475:	data_out=16'h8a00;
17'h7476:	data_out=16'ha00;
17'h7477:	data_out=16'h8998;
17'h7478:	data_out=16'h9ed;
17'h7479:	data_out=16'h9f0;
17'h747a:	data_out=16'h89f5;
17'h747b:	data_out=16'h9ff;
17'h747c:	data_out=16'h9f3;
17'h747d:	data_out=16'h89b4;
17'h747e:	data_out=16'h89cd;
17'h747f:	data_out=16'h805e;
17'h7480:	data_out=16'h9c4;
17'h7481:	data_out=16'h8f2;
17'h7482:	data_out=16'h85d;
17'h7483:	data_out=16'h8984;
17'h7484:	data_out=16'h6a3;
17'h7485:	data_out=16'h89f2;
17'h7486:	data_out=16'h8a00;
17'h7487:	data_out=16'h8a00;
17'h7488:	data_out=16'h9b1;
17'h7489:	data_out=16'h89c9;
17'h748a:	data_out=16'h89f1;
17'h748b:	data_out=16'h866a;
17'h748c:	data_out=16'h89ee;
17'h748d:	data_out=16'h89f6;
17'h748e:	data_out=16'ha00;
17'h748f:	data_out=16'h9f0;
17'h7490:	data_out=16'h89ba;
17'h7491:	data_out=16'h896e;
17'h7492:	data_out=16'h89d9;
17'h7493:	data_out=16'h89c8;
17'h7494:	data_out=16'h89bb;
17'h7495:	data_out=16'h89d1;
17'h7496:	data_out=16'h89cc;
17'h7497:	data_out=16'h89b9;
17'h7498:	data_out=16'h9ca;
17'h7499:	data_out=16'ha00;
17'h749a:	data_out=16'h8897;
17'h749b:	data_out=16'h89db;
17'h749c:	data_out=16'h89bd;
17'h749d:	data_out=16'h8357;
17'h749e:	data_out=16'h89b6;
17'h749f:	data_out=16'h89b5;
17'h74a0:	data_out=16'h8db;
17'h74a1:	data_out=16'ha00;
17'h74a2:	data_out=16'ha00;
17'h74a3:	data_out=16'h8a00;
17'h74a4:	data_out=16'h8a00;
17'h74a5:	data_out=16'h897d;
17'h74a6:	data_out=16'h9ff;
17'h74a7:	data_out=16'h5b0;
17'h74a8:	data_out=16'ha00;
17'h74a9:	data_out=16'h314;
17'h74aa:	data_out=16'h9f7;
17'h74ab:	data_out=16'ha00;
17'h74ac:	data_out=16'h89d5;
17'h74ad:	data_out=16'ha00;
17'h74ae:	data_out=16'h8179;
17'h74af:	data_out=16'h87dd;
17'h74b0:	data_out=16'h888;
17'h74b1:	data_out=16'h89f5;
17'h74b2:	data_out=16'h87e1;
17'h74b3:	data_out=16'h89c6;
17'h74b4:	data_out=16'h99b;
17'h74b5:	data_out=16'h80cb;
17'h74b6:	data_out=16'h9e9;
17'h74b7:	data_out=16'h841d;
17'h74b8:	data_out=16'h89f8;
17'h74b9:	data_out=16'h89c3;
17'h74ba:	data_out=16'h83e1;
17'h74bb:	data_out=16'h89e7;
17'h74bc:	data_out=16'h8927;
17'h74bd:	data_out=16'h9fb;
17'h74be:	data_out=16'ha00;
17'h74bf:	data_out=16'h89f2;
17'h74c0:	data_out=16'h86d2;
17'h74c1:	data_out=16'h8411;
17'h74c2:	data_out=16'h8932;
17'h74c3:	data_out=16'ha00;
17'h74c4:	data_out=16'h8986;
17'h74c5:	data_out=16'h89e6;
17'h74c6:	data_out=16'ha00;
17'h74c7:	data_out=16'h9ff;
17'h74c8:	data_out=16'h89fa;
17'h74c9:	data_out=16'h8946;
17'h74ca:	data_out=16'h9ae;
17'h74cb:	data_out=16'h89f4;
17'h74cc:	data_out=16'h81bd;
17'h74cd:	data_out=16'ha00;
17'h74ce:	data_out=16'h9fa;
17'h74cf:	data_out=16'h8205;
17'h74d0:	data_out=16'h89d8;
17'h74d1:	data_out=16'h89e3;
17'h74d2:	data_out=16'h89e4;
17'h74d3:	data_out=16'h89c1;
17'h74d4:	data_out=16'h997;
17'h74d5:	data_out=16'h89b2;
17'h74d6:	data_out=16'h8a5;
17'h74d7:	data_out=16'h871a;
17'h74d8:	data_out=16'h89fb;
17'h74d9:	data_out=16'h8838;
17'h74da:	data_out=16'h89fa;
17'h74db:	data_out=16'h88e2;
17'h74dc:	data_out=16'h89fe;
17'h74dd:	data_out=16'ha00;
17'h74de:	data_out=16'h89e8;
17'h74df:	data_out=16'h9fc;
17'h74e0:	data_out=16'h517;
17'h74e1:	data_out=16'h88b0;
17'h74e2:	data_out=16'h89cd;
17'h74e3:	data_out=16'h89d7;
17'h74e4:	data_out=16'h8558;
17'h74e5:	data_out=16'h8960;
17'h74e6:	data_out=16'ha00;
17'h74e7:	data_out=16'ha00;
17'h74e8:	data_out=16'ha00;
17'h74e9:	data_out=16'h944;
17'h74ea:	data_out=16'ha00;
17'h74eb:	data_out=16'h89e1;
17'h74ec:	data_out=16'ha00;
17'h74ed:	data_out=16'h89d4;
17'h74ee:	data_out=16'ha00;
17'h74ef:	data_out=16'h8945;
17'h74f0:	data_out=16'ha00;
17'h74f1:	data_out=16'h9b9;
17'h74f2:	data_out=16'h8976;
17'h74f3:	data_out=16'h8942;
17'h74f4:	data_out=16'h722;
17'h74f5:	data_out=16'h8a00;
17'h74f6:	data_out=16'ha00;
17'h74f7:	data_out=16'h8909;
17'h74f8:	data_out=16'ha00;
17'h74f9:	data_out=16'h9ed;
17'h74fa:	data_out=16'h89d0;
17'h74fb:	data_out=16'ha00;
17'h74fc:	data_out=16'h9e0;
17'h74fd:	data_out=16'h89b1;
17'h74fe:	data_out=16'h89b9;
17'h74ff:	data_out=16'h89a1;
17'h7500:	data_out=16'h9ff;
17'h7501:	data_out=16'h8a5;
17'h7502:	data_out=16'h896e;
17'h7503:	data_out=16'h8986;
17'h7504:	data_out=16'h44d;
17'h7505:	data_out=16'h89ea;
17'h7506:	data_out=16'h8a00;
17'h7507:	data_out=16'h8a00;
17'h7508:	data_out=16'h930;
17'h7509:	data_out=16'h89ec;
17'h750a:	data_out=16'h89f4;
17'h750b:	data_out=16'h895a;
17'h750c:	data_out=16'h8a00;
17'h750d:	data_out=16'h8a00;
17'h750e:	data_out=16'h9ff;
17'h750f:	data_out=16'h38e;
17'h7510:	data_out=16'h899c;
17'h7511:	data_out=16'h89e4;
17'h7512:	data_out=16'h89f0;
17'h7513:	data_out=16'h89d1;
17'h7514:	data_out=16'h89d3;
17'h7515:	data_out=16'h5ae;
17'h7516:	data_out=16'h89ca;
17'h7517:	data_out=16'h89d3;
17'h7518:	data_out=16'h507;
17'h7519:	data_out=16'ha00;
17'h751a:	data_out=16'h8909;
17'h751b:	data_out=16'h89f3;
17'h751c:	data_out=16'h891c;
17'h751d:	data_out=16'h2b1;
17'h751e:	data_out=16'h89c7;
17'h751f:	data_out=16'h89d0;
17'h7520:	data_out=16'h9bf;
17'h7521:	data_out=16'h9ff;
17'h7522:	data_out=16'h344;
17'h7523:	data_out=16'h8a00;
17'h7524:	data_out=16'h8a00;
17'h7525:	data_out=16'h89d1;
17'h7526:	data_out=16'h664;
17'h7527:	data_out=16'h232;
17'h7528:	data_out=16'h9ff;
17'h7529:	data_out=16'h112;
17'h752a:	data_out=16'h80a;
17'h752b:	data_out=16'h9e7;
17'h752c:	data_out=16'h89cf;
17'h752d:	data_out=16'h9d8;
17'h752e:	data_out=16'h8a00;
17'h752f:	data_out=16'h576;
17'h7530:	data_out=16'ha00;
17'h7531:	data_out=16'h89f9;
17'h7532:	data_out=16'h8924;
17'h7533:	data_out=16'h89d3;
17'h7534:	data_out=16'h8a7;
17'h7535:	data_out=16'h8741;
17'h7536:	data_out=16'h9b3;
17'h7537:	data_out=16'h89ef;
17'h7538:	data_out=16'h89fd;
17'h7539:	data_out=16'h89cf;
17'h753a:	data_out=16'h89e2;
17'h753b:	data_out=16'h89f7;
17'h753c:	data_out=16'h88ff;
17'h753d:	data_out=16'h9f9;
17'h753e:	data_out=16'h9ff;
17'h753f:	data_out=16'h89ea;
17'h7540:	data_out=16'h88b8;
17'h7541:	data_out=16'h9e6;
17'h7542:	data_out=16'h827a;
17'h7543:	data_out=16'ha00;
17'h7544:	data_out=16'h8990;
17'h7545:	data_out=16'h561;
17'h7546:	data_out=16'ha00;
17'h7547:	data_out=16'h829b;
17'h7548:	data_out=16'h89ff;
17'h7549:	data_out=16'h8930;
17'h754a:	data_out=16'h77d;
17'h754b:	data_out=16'h89f1;
17'h754c:	data_out=16'h8889;
17'h754d:	data_out=16'h9fc;
17'h754e:	data_out=16'h9c2;
17'h754f:	data_out=16'h89d9;
17'h7550:	data_out=16'h89ba;
17'h7551:	data_out=16'h8a00;
17'h7552:	data_out=16'h8a00;
17'h7553:	data_out=16'h89e4;
17'h7554:	data_out=16'h998;
17'h7555:	data_out=16'h89d3;
17'h7556:	data_out=16'h857;
17'h7557:	data_out=16'h88a3;
17'h7558:	data_out=16'h89fc;
17'h7559:	data_out=16'h825a;
17'h755a:	data_out=16'h8a00;
17'h755b:	data_out=16'h3d4;
17'h755c:	data_out=16'h89ff;
17'h755d:	data_out=16'ha00;
17'h755e:	data_out=16'h5f2;
17'h755f:	data_out=16'h9f7;
17'h7560:	data_out=16'h89eb;
17'h7561:	data_out=16'h891a;
17'h7562:	data_out=16'h89f3;
17'h7563:	data_out=16'h89e4;
17'h7564:	data_out=16'h5d3;
17'h7565:	data_out=16'h89ca;
17'h7566:	data_out=16'ha00;
17'h7567:	data_out=16'ha00;
17'h7568:	data_out=16'h9ff;
17'h7569:	data_out=16'h7df;
17'h756a:	data_out=16'h9ff;
17'h756b:	data_out=16'h89c0;
17'h756c:	data_out=16'ha00;
17'h756d:	data_out=16'h89e1;
17'h756e:	data_out=16'h9ff;
17'h756f:	data_out=16'h89b6;
17'h7570:	data_out=16'h9ff;
17'h7571:	data_out=16'h89e0;
17'h7572:	data_out=16'h8916;
17'h7573:	data_out=16'h8914;
17'h7574:	data_out=16'h7f9;
17'h7575:	data_out=16'h8a00;
17'h7576:	data_out=16'ha00;
17'h7577:	data_out=16'h89c4;
17'h7578:	data_out=16'h9ff;
17'h7579:	data_out=16'h9fc;
17'h757a:	data_out=16'h89df;
17'h757b:	data_out=16'h9ff;
17'h757c:	data_out=16'h8d8;
17'h757d:	data_out=16'h89c1;
17'h757e:	data_out=16'h89e7;
17'h757f:	data_out=16'h886a;
17'h7580:	data_out=16'h9eb;
17'h7581:	data_out=16'h951;
17'h7582:	data_out=16'h8659;
17'h7583:	data_out=16'h46e;
17'h7584:	data_out=16'h667;
17'h7585:	data_out=16'h89ff;
17'h7586:	data_out=16'h8a00;
17'h7587:	data_out=16'h8a00;
17'h7588:	data_out=16'h878;
17'h7589:	data_out=16'h8a00;
17'h758a:	data_out=16'h8a00;
17'h758b:	data_out=16'h89c2;
17'h758c:	data_out=16'h89ff;
17'h758d:	data_out=16'h89c4;
17'h758e:	data_out=16'h9fd;
17'h758f:	data_out=16'h806f;
17'h7590:	data_out=16'h8036;
17'h7591:	data_out=16'h8029;
17'h7592:	data_out=16'h89fb;
17'h7593:	data_out=16'h89bc;
17'h7594:	data_out=16'h89fc;
17'h7595:	data_out=16'h9e6;
17'h7596:	data_out=16'h628;
17'h7597:	data_out=16'h8a00;
17'h7598:	data_out=16'h83ea;
17'h7599:	data_out=16'h9f2;
17'h759a:	data_out=16'h839c;
17'h759b:	data_out=16'h89f7;
17'h759c:	data_out=16'h9d8;
17'h759d:	data_out=16'h3fb;
17'h759e:	data_out=16'h89d3;
17'h759f:	data_out=16'h89f9;
17'h75a0:	data_out=16'h981;
17'h75a1:	data_out=16'h9fd;
17'h75a2:	data_out=16'h84fd;
17'h75a3:	data_out=16'h8a00;
17'h75a4:	data_out=16'h8a00;
17'h75a5:	data_out=16'h89c1;
17'h75a6:	data_out=16'h815e;
17'h75a7:	data_out=16'h711;
17'h75a8:	data_out=16'h9fd;
17'h75a9:	data_out=16'h9f4;
17'h75aa:	data_out=16'h967;
17'h75ab:	data_out=16'h7c2;
17'h75ac:	data_out=16'h595;
17'h75ad:	data_out=16'h81b5;
17'h75ae:	data_out=16'h8a00;
17'h75af:	data_out=16'h8e6;
17'h75b0:	data_out=16'ha00;
17'h75b1:	data_out=16'h1e2;
17'h75b2:	data_out=16'h89c0;
17'h75b3:	data_out=16'h89fa;
17'h75b4:	data_out=16'h8cf;
17'h75b5:	data_out=16'hb2;
17'h75b6:	data_out=16'h95d;
17'h75b7:	data_out=16'h89f8;
17'h75b8:	data_out=16'h8a00;
17'h75b9:	data_out=16'h89ee;
17'h75ba:	data_out=16'h89e6;
17'h75bb:	data_out=16'h8a00;
17'h75bc:	data_out=16'h801b;
17'h75bd:	data_out=16'h9d8;
17'h75be:	data_out=16'h9fd;
17'h75bf:	data_out=16'h89fd;
17'h75c0:	data_out=16'heb;
17'h75c1:	data_out=16'h9d5;
17'h75c2:	data_out=16'h85b;
17'h75c3:	data_out=16'h9ff;
17'h75c4:	data_out=16'h71d;
17'h75c5:	data_out=16'h9d7;
17'h75c6:	data_out=16'h9fe;
17'h75c7:	data_out=16'h89da;
17'h75c8:	data_out=16'h8a00;
17'h75c9:	data_out=16'h893b;
17'h75ca:	data_out=16'h83df;
17'h75cb:	data_out=16'h514;
17'h75cc:	data_out=16'h8966;
17'h75cd:	data_out=16'h851f;
17'h75ce:	data_out=16'h774;
17'h75cf:	data_out=16'h89dd;
17'h75d0:	data_out=16'h89a6;
17'h75d1:	data_out=16'h8a00;
17'h75d2:	data_out=16'h8a00;
17'h75d3:	data_out=16'h89fa;
17'h75d4:	data_out=16'h807;
17'h75d5:	data_out=16'h89e8;
17'h75d6:	data_out=16'h9cd;
17'h75d7:	data_out=16'h88c4;
17'h75d8:	data_out=16'h89fc;
17'h75d9:	data_out=16'h6a5;
17'h75da:	data_out=16'h8a00;
17'h75db:	data_out=16'h96b;
17'h75dc:	data_out=16'h8a00;
17'h75dd:	data_out=16'ha00;
17'h75de:	data_out=16'h9fe;
17'h75df:	data_out=16'h9de;
17'h75e0:	data_out=16'h8a00;
17'h75e1:	data_out=16'h8068;
17'h75e2:	data_out=16'h8a00;
17'h75e3:	data_out=16'h89fe;
17'h75e4:	data_out=16'h4ec;
17'h75e5:	data_out=16'h89e7;
17'h75e6:	data_out=16'h9f0;
17'h75e7:	data_out=16'ha00;
17'h75e8:	data_out=16'h9fd;
17'h75e9:	data_out=16'h875;
17'h75ea:	data_out=16'h9fd;
17'h75eb:	data_out=16'h89a8;
17'h75ec:	data_out=16'h9e1;
17'h75ed:	data_out=16'h89fd;
17'h75ee:	data_out=16'h9fd;
17'h75ef:	data_out=16'h89e0;
17'h75f0:	data_out=16'h9fd;
17'h75f1:	data_out=16'h89ff;
17'h75f2:	data_out=16'h89ab;
17'h75f3:	data_out=16'h89e8;
17'h75f4:	data_out=16'h82b;
17'h75f5:	data_out=16'h8a00;
17'h75f6:	data_out=16'h9e7;
17'h75f7:	data_out=16'h8512;
17'h75f8:	data_out=16'h9f3;
17'h75f9:	data_out=16'h9fc;
17'h75fa:	data_out=16'h8a00;
17'h75fb:	data_out=16'h9fd;
17'h75fc:	data_out=16'h86a6;
17'h75fd:	data_out=16'h89ef;
17'h75fe:	data_out=16'h8a00;
17'h75ff:	data_out=16'h85eb;
17'h7600:	data_out=16'h9d6;
17'h7601:	data_out=16'h962;
17'h7602:	data_out=16'h8045;
17'h7603:	data_out=16'h850;
17'h7604:	data_out=16'h7d0;
17'h7605:	data_out=16'h8430;
17'h7606:	data_out=16'h8a00;
17'h7607:	data_out=16'h8a00;
17'h7608:	data_out=16'h7d4;
17'h7609:	data_out=16'h89f6;
17'h760a:	data_out=16'h8a00;
17'h760b:	data_out=16'h848d;
17'h760c:	data_out=16'h8a00;
17'h760d:	data_out=16'h89cf;
17'h760e:	data_out=16'h9fe;
17'h760f:	data_out=16'h869e;
17'h7610:	data_out=16'h8ff;
17'h7611:	data_out=16'h948;
17'h7612:	data_out=16'h8a00;
17'h7613:	data_out=16'h89df;
17'h7614:	data_out=16'h8a00;
17'h7615:	data_out=16'h96c;
17'h7616:	data_out=16'h32b;
17'h7617:	data_out=16'h8a00;
17'h7618:	data_out=16'h8a00;
17'h7619:	data_out=16'h9d6;
17'h761a:	data_out=16'h843a;
17'h761b:	data_out=16'h89e8;
17'h761c:	data_out=16'h9d7;
17'h761d:	data_out=16'h85c;
17'h761e:	data_out=16'h89c4;
17'h761f:	data_out=16'h89fb;
17'h7620:	data_out=16'h75a;
17'h7621:	data_out=16'h9fe;
17'h7622:	data_out=16'h8149;
17'h7623:	data_out=16'h89e8;
17'h7624:	data_out=16'h89e7;
17'h7625:	data_out=16'h899d;
17'h7626:	data_out=16'h82a9;
17'h7627:	data_out=16'h863;
17'h7628:	data_out=16'h9fe;
17'h7629:	data_out=16'ha00;
17'h762a:	data_out=16'h8fb;
17'h762b:	data_out=16'h89fe;
17'h762c:	data_out=16'h126;
17'h762d:	data_out=16'h256;
17'h762e:	data_out=16'h8a00;
17'h762f:	data_out=16'h8f2;
17'h7630:	data_out=16'h828;
17'h7631:	data_out=16'h9ad;
17'h7632:	data_out=16'h86aa;
17'h7633:	data_out=16'h89f9;
17'h7634:	data_out=16'h899;
17'h7635:	data_out=16'h729;
17'h7636:	data_out=16'h886;
17'h7637:	data_out=16'h88a3;
17'h7638:	data_out=16'h8a00;
17'h7639:	data_out=16'h89d6;
17'h763a:	data_out=16'h89eb;
17'h763b:	data_out=16'h8a00;
17'h763c:	data_out=16'h9bd;
17'h763d:	data_out=16'h982;
17'h763e:	data_out=16'h9fe;
17'h763f:	data_out=16'h845f;
17'h7640:	data_out=16'h586;
17'h7641:	data_out=16'h9ce;
17'h7642:	data_out=16'h983;
17'h7643:	data_out=16'h9ff;
17'h7644:	data_out=16'h890;
17'h7645:	data_out=16'h956;
17'h7646:	data_out=16'h9fd;
17'h7647:	data_out=16'h8a00;
17'h7648:	data_out=16'h8a00;
17'h7649:	data_out=16'h8945;
17'h764a:	data_out=16'h8765;
17'h764b:	data_out=16'h95a;
17'h764c:	data_out=16'h89ce;
17'h764d:	data_out=16'h82e0;
17'h764e:	data_out=16'h4ee;
17'h764f:	data_out=16'h89db;
17'h7650:	data_out=16'h896f;
17'h7651:	data_out=16'h89f4;
17'h7652:	data_out=16'h89fd;
17'h7653:	data_out=16'h9d;
17'h7654:	data_out=16'h614;
17'h7655:	data_out=16'h89cc;
17'h7656:	data_out=16'h9e3;
17'h7657:	data_out=16'h898a;
17'h7658:	data_out=16'h89f4;
17'h7659:	data_out=16'h82d;
17'h765a:	data_out=16'h8a00;
17'h765b:	data_out=16'h940;
17'h765c:	data_out=16'h9bb;
17'h765d:	data_out=16'h9f9;
17'h765e:	data_out=16'ha00;
17'h765f:	data_out=16'h862d;
17'h7660:	data_out=16'h8a00;
17'h7661:	data_out=16'h8e1;
17'h7662:	data_out=16'h8a00;
17'h7663:	data_out=16'h8a00;
17'h7664:	data_out=16'h45c;
17'h7665:	data_out=16'h8584;
17'h7666:	data_out=16'h8442;
17'h7667:	data_out=16'ha00;
17'h7668:	data_out=16'h9ff;
17'h7669:	data_out=16'h6c4;
17'h766a:	data_out=16'h9fe;
17'h766b:	data_out=16'h894b;
17'h766c:	data_out=16'h9bc;
17'h766d:	data_out=16'h8a00;
17'h766e:	data_out=16'h9fe;
17'h766f:	data_out=16'h89d5;
17'h7670:	data_out=16'h9fe;
17'h7671:	data_out=16'h8a00;
17'h7672:	data_out=16'h8029;
17'h7673:	data_out=16'h85a1;
17'h7674:	data_out=16'h4cb;
17'h7675:	data_out=16'h899c;
17'h7676:	data_out=16'h8773;
17'h7677:	data_out=16'h81a4;
17'h7678:	data_out=16'h9c3;
17'h7679:	data_out=16'h9f6;
17'h767a:	data_out=16'h8a00;
17'h767b:	data_out=16'h9fe;
17'h767c:	data_out=16'h8a00;
17'h767d:	data_out=16'h89ea;
17'h767e:	data_out=16'h8a00;
17'h767f:	data_out=16'h89a4;
17'h7680:	data_out=16'h958;
17'h7681:	data_out=16'h831f;
17'h7682:	data_out=16'hf0;
17'h7683:	data_out=16'h90a;
17'h7684:	data_out=16'h87a;
17'h7685:	data_out=16'h899f;
17'h7686:	data_out=16'h8a00;
17'h7687:	data_out=16'h8a00;
17'h7688:	data_out=16'h83d;
17'h7689:	data_out=16'h89f9;
17'h768a:	data_out=16'h8735;
17'h768b:	data_out=16'h9de;
17'h768c:	data_out=16'h89ff;
17'h768d:	data_out=16'h89f5;
17'h768e:	data_out=16'h9fb;
17'h768f:	data_out=16'h8a00;
17'h7690:	data_out=16'h975;
17'h7691:	data_out=16'h9df;
17'h7692:	data_out=16'h8a00;
17'h7693:	data_out=16'h898b;
17'h7694:	data_out=16'h89bc;
17'h7695:	data_out=16'h86a9;
17'h7696:	data_out=16'h89b7;
17'h7697:	data_out=16'h89b7;
17'h7698:	data_out=16'h8a00;
17'h7699:	data_out=16'h80ce;
17'h769a:	data_out=16'h891a;
17'h769b:	data_out=16'h9e9;
17'h769c:	data_out=16'h9df;
17'h769d:	data_out=16'h950;
17'h769e:	data_out=16'h89c7;
17'h769f:	data_out=16'h89fa;
17'h76a0:	data_out=16'h866e;
17'h76a1:	data_out=16'h9fb;
17'h76a2:	data_out=16'h9c3;
17'h76a3:	data_out=16'h89ea;
17'h76a4:	data_out=16'h89ea;
17'h76a5:	data_out=16'h8992;
17'h76a6:	data_out=16'h45f;
17'h76a7:	data_out=16'h951;
17'h76a8:	data_out=16'h9fa;
17'h76a9:	data_out=16'ha00;
17'h76aa:	data_out=16'h89ff;
17'h76ab:	data_out=16'h8a00;
17'h76ac:	data_out=16'h89a2;
17'h76ad:	data_out=16'h643;
17'h76ae:	data_out=16'h8a00;
17'h76af:	data_out=16'h90c;
17'h76b0:	data_out=16'h1bf;
17'h76b1:	data_out=16'h9e6;
17'h76b2:	data_out=16'h8831;
17'h76b3:	data_out=16'h89e4;
17'h76b4:	data_out=16'h692;
17'h76b5:	data_out=16'h901;
17'h76b6:	data_out=16'h85c;
17'h76b7:	data_out=16'h68;
17'h76b8:	data_out=16'h8a00;
17'h76b9:	data_out=16'h89da;
17'h76ba:	data_out=16'h89f7;
17'h76bb:	data_out=16'h8a00;
17'h76bc:	data_out=16'h9f6;
17'h76bd:	data_out=16'h818;
17'h76be:	data_out=16'h9fa;
17'h76bf:	data_out=16'h899e;
17'h76c0:	data_out=16'h808e;
17'h76c1:	data_out=16'h9ed;
17'h76c2:	data_out=16'h9f7;
17'h76c3:	data_out=16'ha00;
17'h76c4:	data_out=16'h338;
17'h76c5:	data_out=16'h85db;
17'h76c6:	data_out=16'h9ed;
17'h76c7:	data_out=16'h8a00;
17'h76c8:	data_out=16'h8a00;
17'h76c9:	data_out=16'h88e1;
17'h76ca:	data_out=16'h89ff;
17'h76cb:	data_out=16'h9f5;
17'h76cc:	data_out=16'h89f3;
17'h76cd:	data_out=16'h984;
17'h76ce:	data_out=16'h8674;
17'h76cf:	data_out=16'h89f1;
17'h76d0:	data_out=16'h896f;
17'h76d1:	data_out=16'h89e9;
17'h76d2:	data_out=16'h89ee;
17'h76d3:	data_out=16'h3e7;
17'h76d4:	data_out=16'hab;
17'h76d5:	data_out=16'h89aa;
17'h76d6:	data_out=16'h9dd;
17'h76d7:	data_out=16'h899f;
17'h76d8:	data_out=16'h722;
17'h76d9:	data_out=16'h52;
17'h76da:	data_out=16'h811a;
17'h76db:	data_out=16'h644;
17'h76dc:	data_out=16'h9f0;
17'h76dd:	data_out=16'h9df;
17'h76de:	data_out=16'h9ff;
17'h76df:	data_out=16'h8a00;
17'h76e0:	data_out=16'h84b7;
17'h76e1:	data_out=16'h94d;
17'h76e2:	data_out=16'h8913;
17'h76e3:	data_out=16'h89f6;
17'h76e4:	data_out=16'h809;
17'h76e5:	data_out=16'h98e;
17'h76e6:	data_out=16'h89c0;
17'h76e7:	data_out=16'h9e8;
17'h76e8:	data_out=16'h9fa;
17'h76e9:	data_out=16'h74d;
17'h76ea:	data_out=16'h9fb;
17'h76eb:	data_out=16'h88d2;
17'h76ec:	data_out=16'h884;
17'h76ed:	data_out=16'h89f2;
17'h76ee:	data_out=16'h9fb;
17'h76ef:	data_out=16'h89e6;
17'h76f0:	data_out=16'h9fb;
17'h76f1:	data_out=16'h8a00;
17'h76f2:	data_out=16'h87d5;
17'h76f3:	data_out=16'h871b;
17'h76f4:	data_out=16'h80b2;
17'h76f5:	data_out=16'h9bf;
17'h76f6:	data_out=16'h89f1;
17'h76f7:	data_out=16'h7b1;
17'h76f8:	data_out=16'h9b5;
17'h76f9:	data_out=16'h9e5;
17'h76fa:	data_out=16'h89e1;
17'h76fb:	data_out=16'h9fa;
17'h76fc:	data_out=16'h8a00;
17'h76fd:	data_out=16'h89f6;
17'h76fe:	data_out=16'h86b3;
17'h76ff:	data_out=16'h89c1;
17'h7700:	data_out=16'h9ce;
17'h7701:	data_out=16'h9b0;
17'h7702:	data_out=16'h89ff;
17'h7703:	data_out=16'h9e9;
17'h7704:	data_out=16'h95d;
17'h7705:	data_out=16'h3e6;
17'h7706:	data_out=16'h89fc;
17'h7707:	data_out=16'h8a00;
17'h7708:	data_out=16'h9d5;
17'h7709:	data_out=16'h8a00;
17'h770a:	data_out=16'h100;
17'h770b:	data_out=16'ha00;
17'h770c:	data_out=16'h89e4;
17'h770d:	data_out=16'h89fb;
17'h770e:	data_out=16'h8566;
17'h770f:	data_out=16'h89ff;
17'h7710:	data_out=16'h9ad;
17'h7711:	data_out=16'h9fc;
17'h7712:	data_out=16'h8a00;
17'h7713:	data_out=16'h433;
17'h7714:	data_out=16'h9c5;
17'h7715:	data_out=16'h242;
17'h7716:	data_out=16'h5b7;
17'h7717:	data_out=16'h99b;
17'h7718:	data_out=16'h8a00;
17'h7719:	data_out=16'h85ca;
17'h771a:	data_out=16'h89d1;
17'h771b:	data_out=16'ha00;
17'h771c:	data_out=16'h9ff;
17'h771d:	data_out=16'h9d3;
17'h771e:	data_out=16'h81cc;
17'h771f:	data_out=16'h8a00;
17'h7720:	data_out=16'h8d4;
17'h7721:	data_out=16'h8574;
17'h7722:	data_out=16'h987;
17'h7723:	data_out=16'h8a00;
17'h7724:	data_out=16'h8a00;
17'h7725:	data_out=16'h89fe;
17'h7726:	data_out=16'h236;
17'h7727:	data_out=16'h9aa;
17'h7728:	data_out=16'h82c6;
17'h7729:	data_out=16'ha00;
17'h772a:	data_out=16'h8a00;
17'h772b:	data_out=16'h898f;
17'h772c:	data_out=16'h5c8;
17'h772d:	data_out=16'h7c0;
17'h772e:	data_out=16'h89f7;
17'h772f:	data_out=16'h9c2;
17'h7730:	data_out=16'h8202;
17'h7731:	data_out=16'h9fb;
17'h7732:	data_out=16'h8a00;
17'h7733:	data_out=16'h126;
17'h7734:	data_out=16'h57a;
17'h7735:	data_out=16'h9a1;
17'h7736:	data_out=16'h997;
17'h7737:	data_out=16'h89fe;
17'h7738:	data_out=16'h9ce;
17'h7739:	data_out=16'h830c;
17'h773a:	data_out=16'h8a00;
17'h773b:	data_out=16'h89fe;
17'h773c:	data_out=16'h9fb;
17'h773d:	data_out=16'h832;
17'h773e:	data_out=16'h8299;
17'h773f:	data_out=16'h37d;
17'h7740:	data_out=16'h8a00;
17'h7741:	data_out=16'ha00;
17'h7742:	data_out=16'h9ff;
17'h7743:	data_out=16'ha00;
17'h7744:	data_out=16'h99d;
17'h7745:	data_out=16'h3f2;
17'h7746:	data_out=16'h9fe;
17'h7747:	data_out=16'h8a00;
17'h7748:	data_out=16'h89fb;
17'h7749:	data_out=16'h852c;
17'h774a:	data_out=16'h87e1;
17'h774b:	data_out=16'ha00;
17'h774c:	data_out=16'h8a00;
17'h774d:	data_out=16'h7ca;
17'h774e:	data_out=16'h83a2;
17'h774f:	data_out=16'h8a00;
17'h7750:	data_out=16'h81b6;
17'h7751:	data_out=16'h89fc;
17'h7752:	data_out=16'h8a00;
17'h7753:	data_out=16'h9e4;
17'h7754:	data_out=16'h81d;
17'h7755:	data_out=16'h89c7;
17'h7756:	data_out=16'h8129;
17'h7757:	data_out=16'h8a00;
17'h7758:	data_out=16'h9f4;
17'h7759:	data_out=16'h8a00;
17'h775a:	data_out=16'ha00;
17'h775b:	data_out=16'h73d;
17'h775c:	data_out=16'ha00;
17'h775d:	data_out=16'h9c7;
17'h775e:	data_out=16'ha00;
17'h775f:	data_out=16'h8a00;
17'h7760:	data_out=16'h8223;
17'h7761:	data_out=16'h863;
17'h7762:	data_out=16'h9f1;
17'h7763:	data_out=16'h32e;
17'h7764:	data_out=16'h9e5;
17'h7765:	data_out=16'h967;
17'h7766:	data_out=16'h89c8;
17'h7767:	data_out=16'h46b;
17'h7768:	data_out=16'h84d9;
17'h7769:	data_out=16'h99f;
17'h776a:	data_out=16'h8599;
17'h776b:	data_out=16'h877d;
17'h776c:	data_out=16'h984;
17'h776d:	data_out=16'h378;
17'h776e:	data_out=16'h8599;
17'h776f:	data_out=16'h8a00;
17'h7770:	data_out=16'h8570;
17'h7771:	data_out=16'h8a00;
17'h7772:	data_out=16'h89dd;
17'h7773:	data_out=16'h89f0;
17'h7774:	data_out=16'h832b;
17'h7775:	data_out=16'h9f4;
17'h7776:	data_out=16'h89ee;
17'h7777:	data_out=16'h904;
17'h7778:	data_out=16'h9d7;
17'h7779:	data_out=16'h91b;
17'h777a:	data_out=16'h9ba;
17'h777b:	data_out=16'h828f;
17'h777c:	data_out=16'h8a00;
17'h777d:	data_out=16'h89fe;
17'h777e:	data_out=16'h9cf;
17'h777f:	data_out=16'h89f4;
17'h7780:	data_out=16'h9f4;
17'h7781:	data_out=16'h9d3;
17'h7782:	data_out=16'h89fc;
17'h7783:	data_out=16'h9e4;
17'h7784:	data_out=16'h85a8;
17'h7785:	data_out=16'h8a00;
17'h7786:	data_out=16'h89ff;
17'h7787:	data_out=16'h8a00;
17'h7788:	data_out=16'h9f2;
17'h7789:	data_out=16'h89c8;
17'h778a:	data_out=16'h9bc;
17'h778b:	data_out=16'ha00;
17'h778c:	data_out=16'h8123;
17'h778d:	data_out=16'h89fc;
17'h778e:	data_out=16'h89f8;
17'h778f:	data_out=16'h89fb;
17'h7790:	data_out=16'h9d8;
17'h7791:	data_out=16'h9fe;
17'h7792:	data_out=16'h89ff;
17'h7793:	data_out=16'h5c3;
17'h7794:	data_out=16'h9f6;
17'h7795:	data_out=16'h5e3;
17'h7796:	data_out=16'h86c;
17'h7797:	data_out=16'h9d2;
17'h7798:	data_out=16'h8a00;
17'h7799:	data_out=16'h8977;
17'h779a:	data_out=16'h8a00;
17'h779b:	data_out=16'ha00;
17'h779c:	data_out=16'ha00;
17'h779d:	data_out=16'h9fd;
17'h779e:	data_out=16'h943;
17'h779f:	data_out=16'h89f9;
17'h77a0:	data_out=16'h9a6;
17'h77a1:	data_out=16'h89f9;
17'h77a2:	data_out=16'h89b5;
17'h77a3:	data_out=16'h8a00;
17'h77a4:	data_out=16'h8a00;
17'h77a5:	data_out=16'h89f5;
17'h77a6:	data_out=16'h8297;
17'h77a7:	data_out=16'h9f1;
17'h77a8:	data_out=16'h89f9;
17'h77a9:	data_out=16'h9eb;
17'h77aa:	data_out=16'h89ff;
17'h77ab:	data_out=16'h97d;
17'h77ac:	data_out=16'h870;
17'h77ad:	data_out=16'h9c8;
17'h77ae:	data_out=16'h8967;
17'h77af:	data_out=16'h9cc;
17'h77b0:	data_out=16'h86ef;
17'h77b1:	data_out=16'h9fa;
17'h77b2:	data_out=16'h8a00;
17'h77b3:	data_out=16'h9ff;
17'h77b4:	data_out=16'h9b2;
17'h77b5:	data_out=16'h8af;
17'h77b6:	data_out=16'h9ca;
17'h77b7:	data_out=16'h89ee;
17'h77b8:	data_out=16'ha00;
17'h77b9:	data_out=16'h9ff;
17'h77ba:	data_out=16'h89f0;
17'h77bb:	data_out=16'h89fe;
17'h77bc:	data_out=16'h9c9;
17'h77bd:	data_out=16'h6b1;
17'h77be:	data_out=16'h89f9;
17'h77bf:	data_out=16'h8a00;
17'h77c0:	data_out=16'h8a00;
17'h77c1:	data_out=16'ha00;
17'h77c2:	data_out=16'h9d6;
17'h77c3:	data_out=16'ha00;
17'h77c4:	data_out=16'h9b9;
17'h77c5:	data_out=16'h808;
17'h77c6:	data_out=16'h9e9;
17'h77c7:	data_out=16'h8a00;
17'h77c8:	data_out=16'h89ee;
17'h77c9:	data_out=16'h89d9;
17'h77ca:	data_out=16'h882a;
17'h77cb:	data_out=16'h9fd;
17'h77cc:	data_out=16'h8a00;
17'h77cd:	data_out=16'h89e4;
17'h77ce:	data_out=16'h89de;
17'h77cf:	data_out=16'h8a00;
17'h77d0:	data_out=16'h300;
17'h77d1:	data_out=16'h89da;
17'h77d2:	data_out=16'h8a00;
17'h77d3:	data_out=16'h9ff;
17'h77d4:	data_out=16'h876;
17'h77d5:	data_out=16'h83bc;
17'h77d6:	data_out=16'h89bf;
17'h77d7:	data_out=16'h89fe;
17'h77d8:	data_out=16'h9ff;
17'h77d9:	data_out=16'h8a00;
17'h77da:	data_out=16'ha00;
17'h77db:	data_out=16'h5b6;
17'h77dc:	data_out=16'ha00;
17'h77dd:	data_out=16'h9bb;
17'h77de:	data_out=16'h9ff;
17'h77df:	data_out=16'h89fd;
17'h77e0:	data_out=16'h59d;
17'h77e1:	data_out=16'h830b;
17'h77e2:	data_out=16'ha00;
17'h77e3:	data_out=16'h9f9;
17'h77e4:	data_out=16'h9fe;
17'h77e5:	data_out=16'h38;
17'h77e6:	data_out=16'h88c0;
17'h77e7:	data_out=16'h89d1;
17'h77e8:	data_out=16'h89f9;
17'h77e9:	data_out=16'h9d7;
17'h77ea:	data_out=16'h89f7;
17'h77eb:	data_out=16'h8914;
17'h77ec:	data_out=16'h9b6;
17'h77ed:	data_out=16'h9fa;
17'h77ee:	data_out=16'h89f7;
17'h77ef:	data_out=16'h8a00;
17'h77f0:	data_out=16'h89f7;
17'h77f1:	data_out=16'h8a00;
17'h77f2:	data_out=16'h8a00;
17'h77f3:	data_out=16'h8a00;
17'h77f4:	data_out=16'h8834;
17'h77f5:	data_out=16'h9c5;
17'h77f6:	data_out=16'h89d1;
17'h77f7:	data_out=16'h89a8;
17'h77f8:	data_out=16'h755;
17'h77f9:	data_out=16'h8227;
17'h77fa:	data_out=16'h9f7;
17'h77fb:	data_out=16'h89f9;
17'h77fc:	data_out=16'h8a00;
17'h77fd:	data_out=16'h8a00;
17'h77fe:	data_out=16'ha00;
17'h77ff:	data_out=16'h8a00;
17'h7800:	data_out=16'h9fa;
17'h7801:	data_out=16'h9e5;
17'h7802:	data_out=16'h89ea;
17'h7803:	data_out=16'h8ef;
17'h7804:	data_out=16'h89d0;
17'h7805:	data_out=16'h8a00;
17'h7806:	data_out=16'h8a00;
17'h7807:	data_out=16'h89ff;
17'h7808:	data_out=16'h9ee;
17'h7809:	data_out=16'h89c5;
17'h780a:	data_out=16'h9c3;
17'h780b:	data_out=16'ha00;
17'h780c:	data_out=16'h4db;
17'h780d:	data_out=16'h8a00;
17'h780e:	data_out=16'h89f5;
17'h780f:	data_out=16'h89ca;
17'h7810:	data_out=16'h51f;
17'h7811:	data_out=16'ha00;
17'h7812:	data_out=16'h884e;
17'h7813:	data_out=16'hc0;
17'h7814:	data_out=16'h9af;
17'h7815:	data_out=16'h83b1;
17'h7816:	data_out=16'h65c;
17'h7817:	data_out=16'h97d;
17'h7818:	data_out=16'h89fd;
17'h7819:	data_out=16'h89ba;
17'h781a:	data_out=16'h8a00;
17'h781b:	data_out=16'h9ff;
17'h781c:	data_out=16'h9f0;
17'h781d:	data_out=16'ha00;
17'h781e:	data_out=16'h435;
17'h781f:	data_out=16'h899f;
17'h7820:	data_out=16'h6f0;
17'h7821:	data_out=16'h89f7;
17'h7822:	data_out=16'h89dc;
17'h7823:	data_out=16'h8a00;
17'h7824:	data_out=16'h8a00;
17'h7825:	data_out=16'h8a00;
17'h7826:	data_out=16'h8e4;
17'h7827:	data_out=16'h9fe;
17'h7828:	data_out=16'h89f5;
17'h7829:	data_out=16'h8555;
17'h782a:	data_out=16'h8a00;
17'h782b:	data_out=16'h9fd;
17'h782c:	data_out=16'h621;
17'h782d:	data_out=16'h9f0;
17'h782e:	data_out=16'h8843;
17'h782f:	data_out=16'h982;
17'h7830:	data_out=16'h8a00;
17'h7831:	data_out=16'h9d6;
17'h7832:	data_out=16'h8a00;
17'h7833:	data_out=16'h9fe;
17'h7834:	data_out=16'h9f4;
17'h7835:	data_out=16'h888;
17'h7836:	data_out=16'h9cb;
17'h7837:	data_out=16'h89d6;
17'h7838:	data_out=16'ha00;
17'h7839:	data_out=16'h9ff;
17'h783a:	data_out=16'h89d8;
17'h783b:	data_out=16'h26d;
17'h783c:	data_out=16'h826;
17'h783d:	data_out=16'h20e;
17'h783e:	data_out=16'h89f5;
17'h783f:	data_out=16'h8a00;
17'h7840:	data_out=16'h8a00;
17'h7841:	data_out=16'ha00;
17'h7842:	data_out=16'h941;
17'h7843:	data_out=16'h87fc;
17'h7844:	data_out=16'h99e;
17'h7845:	data_out=16'h828c;
17'h7846:	data_out=16'ha0;
17'h7847:	data_out=16'h89ae;
17'h7848:	data_out=16'h89f3;
17'h7849:	data_out=16'h8a00;
17'h784a:	data_out=16'h8798;
17'h784b:	data_out=16'h9b4;
17'h784c:	data_out=16'h8a00;
17'h784d:	data_out=16'h8a00;
17'h784e:	data_out=16'h89d6;
17'h784f:	data_out=16'h8a00;
17'h7850:	data_out=16'h8a00;
17'h7851:	data_out=16'h89ff;
17'h7852:	data_out=16'h8a00;
17'h7853:	data_out=16'h9f4;
17'h7854:	data_out=16'h348;
17'h7855:	data_out=16'h898e;
17'h7856:	data_out=16'h89fd;
17'h7857:	data_out=16'h8a00;
17'h7858:	data_out=16'h83a5;
17'h7859:	data_out=16'h8a00;
17'h785a:	data_out=16'ha00;
17'h785b:	data_out=16'h9f4;
17'h785c:	data_out=16'h99e;
17'h785d:	data_out=16'h82bc;
17'h785e:	data_out=16'ha00;
17'h785f:	data_out=16'h89ed;
17'h7860:	data_out=16'h965;
17'h7861:	data_out=16'h8a00;
17'h7862:	data_out=16'h9e2;
17'h7863:	data_out=16'h9fd;
17'h7864:	data_out=16'ha00;
17'h7865:	data_out=16'h8a00;
17'h7866:	data_out=16'h88af;
17'h7867:	data_out=16'h89fe;
17'h7868:	data_out=16'h89f8;
17'h7869:	data_out=16'h9d8;
17'h786a:	data_out=16'h89f1;
17'h786b:	data_out=16'h8a00;
17'h786c:	data_out=16'h9e1;
17'h786d:	data_out=16'h9fe;
17'h786e:	data_out=16'h89f2;
17'h786f:	data_out=16'h8a00;
17'h7870:	data_out=16'h89f4;
17'h7871:	data_out=16'h89cb;
17'h7872:	data_out=16'h8a00;
17'h7873:	data_out=16'h8a00;
17'h7874:	data_out=16'h8a00;
17'h7875:	data_out=16'h88b1;
17'h7876:	data_out=16'h852b;
17'h7877:	data_out=16'h89f5;
17'h7878:	data_out=16'h85ba;
17'h7879:	data_out=16'h8994;
17'h787a:	data_out=16'h9d7;
17'h787b:	data_out=16'h89f5;
17'h787c:	data_out=16'h89fc;
17'h787d:	data_out=16'h89d1;
17'h787e:	data_out=16'ha00;
17'h787f:	data_out=16'h8a00;
17'h7880:	data_out=16'h97e;
17'h7881:	data_out=16'h9e0;
17'h7882:	data_out=16'h89db;
17'h7883:	data_out=16'h48c;
17'h7884:	data_out=16'h89d8;
17'h7885:	data_out=16'h89fe;
17'h7886:	data_out=16'h89be;
17'h7887:	data_out=16'h89f9;
17'h7888:	data_out=16'h5f;
17'h7889:	data_out=16'h8999;
17'h788a:	data_out=16'h9b5;
17'h788b:	data_out=16'ha00;
17'h788c:	data_out=16'h86b5;
17'h788d:	data_out=16'h8a00;
17'h788e:	data_out=16'h80bf;
17'h788f:	data_out=16'h89ba;
17'h7890:	data_out=16'h89e7;
17'h7891:	data_out=16'ha00;
17'h7892:	data_out=16'h28f;
17'h7893:	data_out=16'h864a;
17'h7894:	data_out=16'h9f2;
17'h7895:	data_out=16'h89fd;
17'h7896:	data_out=16'h1cf;
17'h7897:	data_out=16'h9db;
17'h7898:	data_out=16'h89fd;
17'h7899:	data_out=16'h89fa;
17'h789a:	data_out=16'h89ff;
17'h789b:	data_out=16'h9f0;
17'h789c:	data_out=16'h68e;
17'h789d:	data_out=16'ha00;
17'h789e:	data_out=16'h982;
17'h789f:	data_out=16'h8927;
17'h78a0:	data_out=16'h8f4;
17'h78a1:	data_out=16'h8216;
17'h78a2:	data_out=16'h89d4;
17'h78a3:	data_out=16'h89fe;
17'h78a4:	data_out=16'h89fe;
17'h78a5:	data_out=16'h8a00;
17'h78a6:	data_out=16'h9c7;
17'h78a7:	data_out=16'h9fe;
17'h78a8:	data_out=16'h8111;
17'h78a9:	data_out=16'h89aa;
17'h78aa:	data_out=16'h8239;
17'h78ab:	data_out=16'h9fd;
17'h78ac:	data_out=16'h8005;
17'h78ad:	data_out=16'h9f7;
17'h78ae:	data_out=16'h83a9;
17'h78af:	data_out=16'h979;
17'h78b0:	data_out=16'h8a00;
17'h78b1:	data_out=16'h9d9;
17'h78b2:	data_out=16'h8a00;
17'h78b3:	data_out=16'h9fe;
17'h78b4:	data_out=16'h9f6;
17'h78b5:	data_out=16'h9c2;
17'h78b6:	data_out=16'h9bd;
17'h78b7:	data_out=16'h896a;
17'h78b8:	data_out=16'ha00;
17'h78b9:	data_out=16'h9fe;
17'h78ba:	data_out=16'h89db;
17'h78bb:	data_out=16'h92b;
17'h78bc:	data_out=16'h85a;
17'h78bd:	data_out=16'h718;
17'h78be:	data_out=16'h80ea;
17'h78bf:	data_out=16'h89fe;
17'h78c0:	data_out=16'h8a00;
17'h78c1:	data_out=16'h9d5;
17'h78c2:	data_out=16'h869;
17'h78c3:	data_out=16'h8860;
17'h78c4:	data_out=16'h9e2;
17'h78c5:	data_out=16'h89b9;
17'h78c6:	data_out=16'h89a0;
17'h78c7:	data_out=16'h264;
17'h78c8:	data_out=16'h89da;
17'h78c9:	data_out=16'h89f8;
17'h78ca:	data_out=16'h86ef;
17'h78cb:	data_out=16'h996;
17'h78cc:	data_out=16'h8a00;
17'h78cd:	data_out=16'h89e8;
17'h78ce:	data_out=16'h256;
17'h78cf:	data_out=16'h8a00;
17'h78d0:	data_out=16'h8a00;
17'h78d1:	data_out=16'h8a00;
17'h78d2:	data_out=16'h89fe;
17'h78d3:	data_out=16'h9d0;
17'h78d4:	data_out=16'h7b8;
17'h78d5:	data_out=16'h8133;
17'h78d6:	data_out=16'h89fb;
17'h78d7:	data_out=16'h89f9;
17'h78d8:	data_out=16'h880b;
17'h78d9:	data_out=16'h8a00;
17'h78da:	data_out=16'h9fc;
17'h78db:	data_out=16'h9ea;
17'h78dc:	data_out=16'h8ce;
17'h78dd:	data_out=16'h865b;
17'h78de:	data_out=16'ha00;
17'h78df:	data_out=16'h89e7;
17'h78e0:	data_out=16'h9ca;
17'h78e1:	data_out=16'h8523;
17'h78e2:	data_out=16'h9f5;
17'h78e3:	data_out=16'h9fa;
17'h78e4:	data_out=16'h9e9;
17'h78e5:	data_out=16'h89fc;
17'h78e6:	data_out=16'h89c8;
17'h78e7:	data_out=16'h8a00;
17'h78e8:	data_out=16'h8228;
17'h78e9:	data_out=16'h46f;
17'h78ea:	data_out=16'h8012;
17'h78eb:	data_out=16'h89f8;
17'h78ec:	data_out=16'h92b;
17'h78ed:	data_out=16'h9fc;
17'h78ee:	data_out=16'h8018;
17'h78ef:	data_out=16'h89ff;
17'h78f0:	data_out=16'h806c;
17'h78f1:	data_out=16'h89b6;
17'h78f2:	data_out=16'h8a00;
17'h78f3:	data_out=16'h8a00;
17'h78f4:	data_out=16'h8a00;
17'h78f5:	data_out=16'h89ea;
17'h78f6:	data_out=16'h9d0;
17'h78f7:	data_out=16'h89f5;
17'h78f8:	data_out=16'h89fb;
17'h78f9:	data_out=16'h89f1;
17'h78fa:	data_out=16'h9f2;
17'h78fb:	data_out=16'h80e4;
17'h78fc:	data_out=16'h89fb;
17'h78fd:	data_out=16'h89af;
17'h78fe:	data_out=16'ha00;
17'h78ff:	data_out=16'h8a00;
17'h7900:	data_out=16'h5e9;
17'h7901:	data_out=16'ha00;
17'h7902:	data_out=16'h82d1;
17'h7903:	data_out=16'h8526;
17'h7904:	data_out=16'h898f;
17'h7905:	data_out=16'h89f8;
17'h7906:	data_out=16'h5c5;
17'h7907:	data_out=16'h8a00;
17'h7908:	data_out=16'h8954;
17'h7909:	data_out=16'h89e5;
17'h790a:	data_out=16'ha00;
17'h790b:	data_out=16'h9fd;
17'h790c:	data_out=16'h89fa;
17'h790d:	data_out=16'h8a00;
17'h790e:	data_out=16'h9f7;
17'h790f:	data_out=16'h89ee;
17'h7910:	data_out=16'h89fd;
17'h7911:	data_out=16'ha00;
17'h7912:	data_out=16'h19;
17'h7913:	data_out=16'h8284;
17'h7914:	data_out=16'h9b7;
17'h7915:	data_out=16'h89fb;
17'h7916:	data_out=16'h89f7;
17'h7917:	data_out=16'h973;
17'h7918:	data_out=16'h8a00;
17'h7919:	data_out=16'h89e6;
17'h791a:	data_out=16'h89f9;
17'h791b:	data_out=16'h9d5;
17'h791c:	data_out=16'h451;
17'h791d:	data_out=16'ha00;
17'h791e:	data_out=16'h97f;
17'h791f:	data_out=16'h89cf;
17'h7920:	data_out=16'h4e9;
17'h7921:	data_out=16'h948;
17'h7922:	data_out=16'h8957;
17'h7923:	data_out=16'h4fb;
17'h7924:	data_out=16'h4ad;
17'h7925:	data_out=16'h89de;
17'h7926:	data_out=16'h9d5;
17'h7927:	data_out=16'h9f8;
17'h7928:	data_out=16'h9aa;
17'h7929:	data_out=16'h833d;
17'h792a:	data_out=16'h1f5;
17'h792b:	data_out=16'h9dd;
17'h792c:	data_out=16'h89f7;
17'h792d:	data_out=16'ha00;
17'h792e:	data_out=16'h9ed;
17'h792f:	data_out=16'h9b;
17'h7930:	data_out=16'h8a00;
17'h7931:	data_out=16'ha00;
17'h7932:	data_out=16'h89f8;
17'h7933:	data_out=16'h9c2;
17'h7934:	data_out=16'ha00;
17'h7935:	data_out=16'h9f0;
17'h7936:	data_out=16'h8305;
17'h7937:	data_out=16'h9cb;
17'h7938:	data_out=16'ha00;
17'h7939:	data_out=16'h999;
17'h793a:	data_out=16'h89e3;
17'h793b:	data_out=16'h9b6;
17'h793c:	data_out=16'h9f9;
17'h793d:	data_out=16'h36e;
17'h793e:	data_out=16'h9b6;
17'h793f:	data_out=16'h89f8;
17'h7940:	data_out=16'h89f8;
17'h7941:	data_out=16'h86f2;
17'h7942:	data_out=16'h8a00;
17'h7943:	data_out=16'h8919;
17'h7944:	data_out=16'h9f7;
17'h7945:	data_out=16'h89fb;
17'h7946:	data_out=16'h9d9;
17'h7947:	data_out=16'h8125;
17'h7948:	data_out=16'h8582;
17'h7949:	data_out=16'h89e0;
17'h794a:	data_out=16'h89d4;
17'h794b:	data_out=16'h84e9;
17'h794c:	data_out=16'h89fe;
17'h794d:	data_out=16'h89d2;
17'h794e:	data_out=16'h343;
17'h794f:	data_out=16'h89ec;
17'h7950:	data_out=16'h89fc;
17'h7951:	data_out=16'h89fb;
17'h7952:	data_out=16'h85db;
17'h7953:	data_out=16'h9c2;
17'h7954:	data_out=16'h97a;
17'h7955:	data_out=16'h93e;
17'h7956:	data_out=16'h8960;
17'h7957:	data_out=16'h84b9;
17'h7958:	data_out=16'h88e7;
17'h7959:	data_out=16'h89f0;
17'h795a:	data_out=16'h9e2;
17'h795b:	data_out=16'ha00;
17'h795c:	data_out=16'h9d1;
17'h795d:	data_out=16'h8548;
17'h795e:	data_out=16'h3ec;
17'h795f:	data_out=16'h88e7;
17'h7960:	data_out=16'h9df;
17'h7961:	data_out=16'h9a0;
17'h7962:	data_out=16'h9ea;
17'h7963:	data_out=16'h9c6;
17'h7964:	data_out=16'h9fb;
17'h7965:	data_out=16'h818a;
17'h7966:	data_out=16'h89cc;
17'h7967:	data_out=16'h89de;
17'h7968:	data_out=16'h943;
17'h7969:	data_out=16'h89d1;
17'h796a:	data_out=16'h9f8;
17'h796b:	data_out=16'h89ed;
17'h796c:	data_out=16'h247;
17'h796d:	data_out=16'h9c5;
17'h796e:	data_out=16'h9f8;
17'h796f:	data_out=16'h89ff;
17'h7970:	data_out=16'h9f8;
17'h7971:	data_out=16'hb4;
17'h7972:	data_out=16'h8906;
17'h7973:	data_out=16'h8470;
17'h7974:	data_out=16'h8a00;
17'h7975:	data_out=16'h977;
17'h7976:	data_out=16'h9e6;
17'h7977:	data_out=16'h89fd;
17'h7978:	data_out=16'h8a00;
17'h7979:	data_out=16'h8a00;
17'h797a:	data_out=16'h9b7;
17'h797b:	data_out=16'h9b7;
17'h797c:	data_out=16'h8a00;
17'h797d:	data_out=16'h89d6;
17'h797e:	data_out=16'ha00;
17'h797f:	data_out=16'h8a00;
17'h7980:	data_out=16'h88dc;
17'h7981:	data_out=16'h9ff;
17'h7982:	data_out=16'h8e1;
17'h7983:	data_out=16'h88fb;
17'h7984:	data_out=16'h85dd;
17'h7985:	data_out=16'h89f0;
17'h7986:	data_out=16'h98e;
17'h7987:	data_out=16'h8a00;
17'h7988:	data_out=16'h897c;
17'h7989:	data_out=16'h89e5;
17'h798a:	data_out=16'ha00;
17'h798b:	data_out=16'h9ef;
17'h798c:	data_out=16'h89d3;
17'h798d:	data_out=16'h8a00;
17'h798e:	data_out=16'h9f9;
17'h798f:	data_out=16'h8972;
17'h7990:	data_out=16'h89f4;
17'h7991:	data_out=16'ha00;
17'h7992:	data_out=16'h1f7;
17'h7993:	data_out=16'h6dc;
17'h7994:	data_out=16'h9bd;
17'h7995:	data_out=16'h89fb;
17'h7996:	data_out=16'h89fe;
17'h7997:	data_out=16'h6a5;
17'h7998:	data_out=16'h8a00;
17'h7999:	data_out=16'h89ad;
17'h799a:	data_out=16'h89ef;
17'h799b:	data_out=16'h9df;
17'h799c:	data_out=16'h18b;
17'h799d:	data_out=16'ha00;
17'h799e:	data_out=16'h999;
17'h799f:	data_out=16'h8222;
17'h79a0:	data_out=16'h80d1;
17'h79a1:	data_out=16'h9f7;
17'h79a2:	data_out=16'h88dc;
17'h79a3:	data_out=16'ha00;
17'h79a4:	data_out=16'ha00;
17'h79a5:	data_out=16'h8950;
17'h79a6:	data_out=16'h8597;
17'h79a7:	data_out=16'h9dd;
17'h79a8:	data_out=16'h9f6;
17'h79a9:	data_out=16'h8170;
17'h79aa:	data_out=16'hd;
17'h79ab:	data_out=16'h62;
17'h79ac:	data_out=16'h89fd;
17'h79ad:	data_out=16'ha00;
17'h79ae:	data_out=16'h9fc;
17'h79af:	data_out=16'h835c;
17'h79b0:	data_out=16'h8a00;
17'h79b1:	data_out=16'ha00;
17'h79b2:	data_out=16'h8783;
17'h79b3:	data_out=16'h993;
17'h79b4:	data_out=16'h9fd;
17'h79b5:	data_out=16'h96b;
17'h79b6:	data_out=16'h83b6;
17'h79b7:	data_out=16'h9e1;
17'h79b8:	data_out=16'h9ff;
17'h79b9:	data_out=16'h7d0;
17'h79ba:	data_out=16'h89e5;
17'h79bb:	data_out=16'h501;
17'h79bc:	data_out=16'ha00;
17'h79bd:	data_out=16'h81bc;
17'h79be:	data_out=16'h9f6;
17'h79bf:	data_out=16'h89f0;
17'h79c0:	data_out=16'h87ff;
17'h79c1:	data_out=16'h8a00;
17'h79c2:	data_out=16'h89ca;
17'h79c3:	data_out=16'h89fb;
17'h79c4:	data_out=16'h9fc;
17'h79c5:	data_out=16'h89fb;
17'h79c6:	data_out=16'h9f7;
17'h79c7:	data_out=16'h87bb;
17'h79c8:	data_out=16'h96b;
17'h79c9:	data_out=16'h88c9;
17'h79ca:	data_out=16'h89ef;
17'h79cb:	data_out=16'h89bf;
17'h79cc:	data_out=16'h89f0;
17'h79cd:	data_out=16'h88e5;
17'h79ce:	data_out=16'h391;
17'h79cf:	data_out=16'h899b;
17'h79d0:	data_out=16'h89fe;
17'h79d1:	data_out=16'h89ff;
17'h79d2:	data_out=16'h8425;
17'h79d3:	data_out=16'h9c9;
17'h79d4:	data_out=16'h82f7;
17'h79d5:	data_out=16'h98d;
17'h79d6:	data_out=16'h81f1;
17'h79d7:	data_out=16'h98c;
17'h79d8:	data_out=16'h89d6;
17'h79d9:	data_out=16'h88cf;
17'h79da:	data_out=16'h96c;
17'h79db:	data_out=16'ha00;
17'h79dc:	data_out=16'h9d5;
17'h79dd:	data_out=16'h882a;
17'h79de:	data_out=16'h80cd;
17'h79df:	data_out=16'h88d9;
17'h79e0:	data_out=16'h9e3;
17'h79e1:	data_out=16'h9b6;
17'h79e2:	data_out=16'h9f1;
17'h79e3:	data_out=16'h98e;
17'h79e4:	data_out=16'h9f3;
17'h79e5:	data_out=16'h8093;
17'h79e6:	data_out=16'h89c5;
17'h79e7:	data_out=16'h89d1;
17'h79e8:	data_out=16'h9f7;
17'h79e9:	data_out=16'h89c4;
17'h79ea:	data_out=16'h9f9;
17'h79eb:	data_out=16'h89e2;
17'h79ec:	data_out=16'h89e4;
17'h79ed:	data_out=16'h992;
17'h79ee:	data_out=16'h9f9;
17'h79ef:	data_out=16'h89fe;
17'h79f0:	data_out=16'h9f9;
17'h79f1:	data_out=16'h573;
17'h79f2:	data_out=16'h8645;
17'h79f3:	data_out=16'h9a5;
17'h79f4:	data_out=16'h8a00;
17'h79f5:	data_out=16'h97e;
17'h79f6:	data_out=16'h9a6;
17'h79f7:	data_out=16'h89ff;
17'h79f8:	data_out=16'h8a00;
17'h79f9:	data_out=16'h8a00;
17'h79fa:	data_out=16'h9af;
17'h79fb:	data_out=16'h9f6;
17'h79fc:	data_out=16'h8a00;
17'h79fd:	data_out=16'h871f;
17'h79fe:	data_out=16'ha00;
17'h79ff:	data_out=16'h8a00;
17'h7a00:	data_out=16'h87b1;
17'h7a01:	data_out=16'h9fe;
17'h7a02:	data_out=16'h9de;
17'h7a03:	data_out=16'h89e0;
17'h7a04:	data_out=16'h83ee;
17'h7a05:	data_out=16'h89f1;
17'h7a06:	data_out=16'h817;
17'h7a07:	data_out=16'h8a00;
17'h7a08:	data_out=16'h8617;
17'h7a09:	data_out=16'h89ff;
17'h7a0a:	data_out=16'ha00;
17'h7a0b:	data_out=16'h328;
17'h7a0c:	data_out=16'h89c5;
17'h7a0d:	data_out=16'h8a00;
17'h7a0e:	data_out=16'h9f7;
17'h7a0f:	data_out=16'h8405;
17'h7a10:	data_out=16'h89fb;
17'h7a11:	data_out=16'ha00;
17'h7a12:	data_out=16'h409;
17'h7a13:	data_out=16'h614;
17'h7a14:	data_out=16'h84a0;
17'h7a15:	data_out=16'h89f7;
17'h7a16:	data_out=16'h89ff;
17'h7a17:	data_out=16'h865a;
17'h7a18:	data_out=16'h8a00;
17'h7a19:	data_out=16'h89d0;
17'h7a1a:	data_out=16'h89f7;
17'h7a1b:	data_out=16'h9ee;
17'h7a1c:	data_out=16'h895d;
17'h7a1d:	data_out=16'ha00;
17'h7a1e:	data_out=16'h810e;
17'h7a1f:	data_out=16'h8465;
17'h7a20:	data_out=16'h85c4;
17'h7a21:	data_out=16'h9f6;
17'h7a22:	data_out=16'h89f4;
17'h7a23:	data_out=16'ha00;
17'h7a24:	data_out=16'ha00;
17'h7a25:	data_out=16'h89fb;
17'h7a26:	data_out=16'h8715;
17'h7a27:	data_out=16'h9fb;
17'h7a28:	data_out=16'h9f5;
17'h7a29:	data_out=16'h89dd;
17'h7a2a:	data_out=16'h491;
17'h7a2b:	data_out=16'h8476;
17'h7a2c:	data_out=16'h89ff;
17'h7a2d:	data_out=16'ha00;
17'h7a2e:	data_out=16'h9fa;
17'h7a2f:	data_out=16'h8774;
17'h7a30:	data_out=16'h8a00;
17'h7a31:	data_out=16'ha00;
17'h7a32:	data_out=16'h885a;
17'h7a33:	data_out=16'h2fc;
17'h7a34:	data_out=16'h9ff;
17'h7a35:	data_out=16'h6c1;
17'h7a36:	data_out=16'h82c7;
17'h7a37:	data_out=16'h9ea;
17'h7a38:	data_out=16'h9fe;
17'h7a39:	data_out=16'h80ed;
17'h7a3a:	data_out=16'h89fd;
17'h7a3b:	data_out=16'h8270;
17'h7a3c:	data_out=16'h9fe;
17'h7a3d:	data_out=16'h86be;
17'h7a3e:	data_out=16'h9f5;
17'h7a3f:	data_out=16'h89f2;
17'h7a40:	data_out=16'h875f;
17'h7a41:	data_out=16'h89ab;
17'h7a42:	data_out=16'h89c9;
17'h7a43:	data_out=16'h89ff;
17'h7a44:	data_out=16'h9ff;
17'h7a45:	data_out=16'h89f8;
17'h7a46:	data_out=16'h9fd;
17'h7a47:	data_out=16'h89e3;
17'h7a48:	data_out=16'h923;
17'h7a49:	data_out=16'h89d0;
17'h7a4a:	data_out=16'h892a;
17'h7a4b:	data_out=16'h89be;
17'h7a4c:	data_out=16'h89fa;
17'h7a4d:	data_out=16'h89ed;
17'h7a4e:	data_out=16'h5f1;
17'h7a4f:	data_out=16'h89c1;
17'h7a50:	data_out=16'h8a00;
17'h7a51:	data_out=16'h89fe;
17'h7a52:	data_out=16'h62;
17'h7a53:	data_out=16'h9f9;
17'h7a54:	data_out=16'h857f;
17'h7a55:	data_out=16'h1c9;
17'h7a56:	data_out=16'h82bb;
17'h7a57:	data_out=16'h837b;
17'h7a58:	data_out=16'h89c4;
17'h7a59:	data_out=16'h895f;
17'h7a5a:	data_out=16'h9ab;
17'h7a5b:	data_out=16'ha00;
17'h7a5c:	data_out=16'h9fc;
17'h7a5d:	data_out=16'h893d;
17'h7a5e:	data_out=16'h866d;
17'h7a5f:	data_out=16'h893d;
17'h7a60:	data_out=16'h967;
17'h7a61:	data_out=16'h9c4;
17'h7a62:	data_out=16'h80ff;
17'h7a63:	data_out=16'h524;
17'h7a64:	data_out=16'h952;
17'h7a65:	data_out=16'h8974;
17'h7a66:	data_out=16'h89c3;
17'h7a67:	data_out=16'h8991;
17'h7a68:	data_out=16'h9f5;
17'h7a69:	data_out=16'h898b;
17'h7a6a:	data_out=16'h9f7;
17'h7a6b:	data_out=16'h89c5;
17'h7a6c:	data_out=16'h8975;
17'h7a6d:	data_out=16'h4f8;
17'h7a6e:	data_out=16'h9f7;
17'h7a6f:	data_out=16'h89fe;
17'h7a70:	data_out=16'h9f7;
17'h7a71:	data_out=16'h6c3;
17'h7a72:	data_out=16'h8981;
17'h7a73:	data_out=16'h88d2;
17'h7a74:	data_out=16'h8a00;
17'h7a75:	data_out=16'h997;
17'h7a76:	data_out=16'h8ba;
17'h7a77:	data_out=16'h89ff;
17'h7a78:	data_out=16'h8a00;
17'h7a79:	data_out=16'h89f2;
17'h7a7a:	data_out=16'h4aa;
17'h7a7b:	data_out=16'h9f5;
17'h7a7c:	data_out=16'h89ff;
17'h7a7d:	data_out=16'h89fe;
17'h7a7e:	data_out=16'ha00;
17'h7a7f:	data_out=16'h8a00;
17'h7a80:	data_out=16'h889a;
17'h7a81:	data_out=16'h201;
17'h7a82:	data_out=16'h117;
17'h7a83:	data_out=16'h89f3;
17'h7a84:	data_out=16'h8773;
17'h7a85:	data_out=16'h89f7;
17'h7a86:	data_out=16'h905;
17'h7a87:	data_out=16'h89ef;
17'h7a88:	data_out=16'h8615;
17'h7a89:	data_out=16'h8a00;
17'h7a8a:	data_out=16'h52d;
17'h7a8b:	data_out=16'h888d;
17'h7a8c:	data_out=16'h89ae;
17'h7a8d:	data_out=16'h8a00;
17'h7a8e:	data_out=16'h9f8;
17'h7a8f:	data_out=16'h8882;
17'h7a90:	data_out=16'h89f8;
17'h7a91:	data_out=16'ha00;
17'h7a92:	data_out=16'h6d9;
17'h7a93:	data_out=16'h678;
17'h7a94:	data_out=16'h89a6;
17'h7a95:	data_out=16'h89f8;
17'h7a96:	data_out=16'h89fd;
17'h7a97:	data_out=16'h89ae;
17'h7a98:	data_out=16'h89f0;
17'h7a99:	data_out=16'h89e5;
17'h7a9a:	data_out=16'h89f7;
17'h7a9b:	data_out=16'h8879;
17'h7a9c:	data_out=16'h89bd;
17'h7a9d:	data_out=16'h9fe;
17'h7a9e:	data_out=16'h89ba;
17'h7a9f:	data_out=16'h89bf;
17'h7aa0:	data_out=16'h895b;
17'h7aa1:	data_out=16'h9f7;
17'h7aa2:	data_out=16'h89ff;
17'h7aa3:	data_out=16'ha00;
17'h7aa4:	data_out=16'ha00;
17'h7aa5:	data_out=16'h89fd;
17'h7aa6:	data_out=16'h85f8;
17'h7aa7:	data_out=16'h816c;
17'h7aa8:	data_out=16'h9f6;
17'h7aa9:	data_out=16'h89f5;
17'h7aaa:	data_out=16'h8721;
17'h7aab:	data_out=16'h8999;
17'h7aac:	data_out=16'h89fd;
17'h7aad:	data_out=16'ha00;
17'h7aae:	data_out=16'h83ed;
17'h7aaf:	data_out=16'h895d;
17'h7ab0:	data_out=16'h8a00;
17'h7ab1:	data_out=16'h9fd;
17'h7ab2:	data_out=16'h89e0;
17'h7ab3:	data_out=16'h89c6;
17'h7ab4:	data_out=16'h1ad;
17'h7ab5:	data_out=16'h81cd;
17'h7ab6:	data_out=16'h864e;
17'h7ab7:	data_out=16'h8a5;
17'h7ab8:	data_out=16'h8f6;
17'h7ab9:	data_out=16'h89d7;
17'h7aba:	data_out=16'h8a00;
17'h7abb:	data_out=16'h8994;
17'h7abc:	data_out=16'h59e;
17'h7abd:	data_out=16'h8994;
17'h7abe:	data_out=16'h9f6;
17'h7abf:	data_out=16'h89f7;
17'h7ac0:	data_out=16'h89c1;
17'h7ac1:	data_out=16'h89a1;
17'h7ac2:	data_out=16'h899c;
17'h7ac3:	data_out=16'h89fe;
17'h7ac4:	data_out=16'h86f4;
17'h7ac5:	data_out=16'h89f9;
17'h7ac6:	data_out=16'h9fc;
17'h7ac7:	data_out=16'h89e3;
17'h7ac8:	data_out=16'h86f3;
17'h7ac9:	data_out=16'h89fa;
17'h7aca:	data_out=16'h88f0;
17'h7acb:	data_out=16'h8958;
17'h7acc:	data_out=16'h89fe;
17'h7acd:	data_out=16'h89fa;
17'h7ace:	data_out=16'h88a0;
17'h7acf:	data_out=16'h89f2;
17'h7ad0:	data_out=16'h89fe;
17'h7ad1:	data_out=16'h89fd;
17'h7ad2:	data_out=16'h52b;
17'h7ad3:	data_out=16'h9fb;
17'h7ad4:	data_out=16'h8841;
17'h7ad5:	data_out=16'h8990;
17'h7ad6:	data_out=16'h832e;
17'h7ad7:	data_out=16'h899b;
17'h7ad8:	data_out=16'h89a2;
17'h7ad9:	data_out=16'h89de;
17'h7ada:	data_out=16'h9f7;
17'h7adb:	data_out=16'ha00;
17'h7adc:	data_out=16'h9fb;
17'h7add:	data_out=16'h89d7;
17'h7ade:	data_out=16'h88e5;
17'h7adf:	data_out=16'h8994;
17'h7ae0:	data_out=16'h57c;
17'h7ae1:	data_out=16'h8db;
17'h7ae2:	data_out=16'h8969;
17'h7ae3:	data_out=16'h88df;
17'h7ae4:	data_out=16'h73d;
17'h7ae5:	data_out=16'h89fe;
17'h7ae6:	data_out=16'h89e0;
17'h7ae7:	data_out=16'h89e9;
17'h7ae8:	data_out=16'h9f7;
17'h7ae9:	data_out=16'h881b;
17'h7aea:	data_out=16'h9f8;
17'h7aeb:	data_out=16'h89f7;
17'h7aec:	data_out=16'h89b4;
17'h7aed:	data_out=16'h89b4;
17'h7aee:	data_out=16'h9f8;
17'h7aef:	data_out=16'h89f9;
17'h7af0:	data_out=16'h9f8;
17'h7af1:	data_out=16'h434;
17'h7af2:	data_out=16'h89f5;
17'h7af3:	data_out=16'h89f5;
17'h7af4:	data_out=16'h89fb;
17'h7af5:	data_out=16'h83f3;
17'h7af6:	data_out=16'h89a0;
17'h7af7:	data_out=16'h8a00;
17'h7af8:	data_out=16'h8a00;
17'h7af9:	data_out=16'h89ce;
17'h7afa:	data_out=16'h899a;
17'h7afb:	data_out=16'h9f6;
17'h7afc:	data_out=16'h83e9;
17'h7afd:	data_out=16'h89f9;
17'h7afe:	data_out=16'ha00;
17'h7aff:	data_out=16'h89ff;
17'h7b00:	data_out=16'h87d8;
17'h7b01:	data_out=16'h9fe;
17'h7b02:	data_out=16'h92b;
17'h7b03:	data_out=16'h89f6;
17'h7b04:	data_out=16'h8075;
17'h7b05:	data_out=16'h89f9;
17'h7b06:	data_out=16'h9f7;
17'h7b07:	data_out=16'h89db;
17'h7b08:	data_out=16'h988;
17'h7b09:	data_out=16'h8a00;
17'h7b0a:	data_out=16'h96f;
17'h7b0b:	data_out=16'h894c;
17'h7b0c:	data_out=16'h89cc;
17'h7b0d:	data_out=16'h89ff;
17'h7b0e:	data_out=16'h9fb;
17'h7b0f:	data_out=16'h3d1;
17'h7b10:	data_out=16'h89ff;
17'h7b11:	data_out=16'ha00;
17'h7b12:	data_out=16'h9e0;
17'h7b13:	data_out=16'h8364;
17'h7b14:	data_out=16'h89b5;
17'h7b15:	data_out=16'h89f8;
17'h7b16:	data_out=16'h89f9;
17'h7b17:	data_out=16'h89b2;
17'h7b18:	data_out=16'h9f9;
17'h7b19:	data_out=16'h89f9;
17'h7b1a:	data_out=16'h89fa;
17'h7b1b:	data_out=16'h88df;
17'h7b1c:	data_out=16'h89c0;
17'h7b1d:	data_out=16'ha00;
17'h7b1e:	data_out=16'h8990;
17'h7b1f:	data_out=16'h8912;
17'h7b20:	data_out=16'h894a;
17'h7b21:	data_out=16'h9fa;
17'h7b22:	data_out=16'h89ff;
17'h7b23:	data_out=16'ha00;
17'h7b24:	data_out=16'ha00;
17'h7b25:	data_out=16'h89ff;
17'h7b26:	data_out=16'h8e8;
17'h7b27:	data_out=16'ha00;
17'h7b28:	data_out=16'h9f9;
17'h7b29:	data_out=16'h89ef;
17'h7b2a:	data_out=16'h7ef;
17'h7b2b:	data_out=16'h89c3;
17'h7b2c:	data_out=16'h89fc;
17'h7b2d:	data_out=16'ha00;
17'h7b2e:	data_out=16'h798;
17'h7b2f:	data_out=16'h893f;
17'h7b30:	data_out=16'h89f9;
17'h7b31:	data_out=16'h736;
17'h7b32:	data_out=16'h89ea;
17'h7b33:	data_out=16'h89ab;
17'h7b34:	data_out=16'h9ff;
17'h7b35:	data_out=16'h8a5;
17'h7b36:	data_out=16'h8678;
17'h7b37:	data_out=16'h83b;
17'h7b38:	data_out=16'h9fa;
17'h7b39:	data_out=16'h89b6;
17'h7b3a:	data_out=16'h8a00;
17'h7b3b:	data_out=16'h15;
17'h7b3c:	data_out=16'h89b2;
17'h7b3d:	data_out=16'h8968;
17'h7b3e:	data_out=16'h9f9;
17'h7b3f:	data_out=16'h89f9;
17'h7b40:	data_out=16'h89ef;
17'h7b41:	data_out=16'h8985;
17'h7b42:	data_out=16'h897d;
17'h7b43:	data_out=16'h89ff;
17'h7b44:	data_out=16'h8648;
17'h7b45:	data_out=16'h89fa;
17'h7b46:	data_out=16'h9ff;
17'h7b47:	data_out=16'h89e7;
17'h7b48:	data_out=16'h86c8;
17'h7b49:	data_out=16'h89fd;
17'h7b4a:	data_out=16'h8908;
17'h7b4b:	data_out=16'h88c6;
17'h7b4c:	data_out=16'h89ff;
17'h7b4d:	data_out=16'h89ff;
17'h7b4e:	data_out=16'h73b;
17'h7b4f:	data_out=16'h89fe;
17'h7b50:	data_out=16'h89fe;
17'h7b51:	data_out=16'h89dc;
17'h7b52:	data_out=16'h9d9;
17'h7b53:	data_out=16'h66a;
17'h7b54:	data_out=16'h88c3;
17'h7b55:	data_out=16'h8977;
17'h7b56:	data_out=16'ha00;
17'h7b57:	data_out=16'h848f;
17'h7b58:	data_out=16'h8974;
17'h7b59:	data_out=16'h89f8;
17'h7b5a:	data_out=16'ha00;
17'h7b5b:	data_out=16'ha00;
17'h7b5c:	data_out=16'h78b;
17'h7b5d:	data_out=16'h89e7;
17'h7b5e:	data_out=16'h893b;
17'h7b5f:	data_out=16'h770;
17'h7b60:	data_out=16'h9f9;
17'h7b61:	data_out=16'h911;
17'h7b62:	data_out=16'h8990;
17'h7b63:	data_out=16'h8990;
17'h7b64:	data_out=16'h736;
17'h7b65:	data_out=16'h8a00;
17'h7b66:	data_out=16'h89ee;
17'h7b67:	data_out=16'h89fd;
17'h7b68:	data_out=16'h9f9;
17'h7b69:	data_out=16'h46a;
17'h7b6a:	data_out=16'h9fc;
17'h7b6b:	data_out=16'h89f9;
17'h7b6c:	data_out=16'h8001;
17'h7b6d:	data_out=16'h8993;
17'h7b6e:	data_out=16'h9fc;
17'h7b6f:	data_out=16'h89fb;
17'h7b70:	data_out=16'h9fb;
17'h7b71:	data_out=16'h9fc;
17'h7b72:	data_out=16'h89fd;
17'h7b73:	data_out=16'h89fa;
17'h7b74:	data_out=16'h89f3;
17'h7b75:	data_out=16'h81b4;
17'h7b76:	data_out=16'h89c7;
17'h7b77:	data_out=16'h8a00;
17'h7b78:	data_out=16'h8a00;
17'h7b79:	data_out=16'h8903;
17'h7b7a:	data_out=16'h898c;
17'h7b7b:	data_out=16'h9f9;
17'h7b7c:	data_out=16'h9fd;
17'h7b7d:	data_out=16'h89f9;
17'h7b7e:	data_out=16'h5dd;
17'h7b7f:	data_out=16'h8a00;
17'h7b80:	data_out=16'ha00;
17'h7b81:	data_out=16'ha00;
17'h7b82:	data_out=16'ha00;
17'h7b83:	data_out=16'h89fc;
17'h7b84:	data_out=16'ha00;
17'h7b85:	data_out=16'h89af;
17'h7b86:	data_out=16'h4e4;
17'h7b87:	data_out=16'h89f2;
17'h7b88:	data_out=16'ha00;
17'h7b89:	data_out=16'h8a00;
17'h7b8a:	data_out=16'ha00;
17'h7b8b:	data_out=16'h89d8;
17'h7b8c:	data_out=16'h89ff;
17'h7b8d:	data_out=16'h897b;
17'h7b8e:	data_out=16'ha00;
17'h7b8f:	data_out=16'ha00;
17'h7b90:	data_out=16'h8a00;
17'h7b91:	data_out=16'ha00;
17'h7b92:	data_out=16'ha00;
17'h7b93:	data_out=16'h873b;
17'h7b94:	data_out=16'h89fe;
17'h7b95:	data_out=16'ha00;
17'h7b96:	data_out=16'h4d9;
17'h7b97:	data_out=16'h8a00;
17'h7b98:	data_out=16'ha00;
17'h7b99:	data_out=16'h8a00;
17'h7b9a:	data_out=16'h89ea;
17'h7b9b:	data_out=16'h89b4;
17'h7b9c:	data_out=16'h88ba;
17'h7b9d:	data_out=16'ha00;
17'h7b9e:	data_out=16'h8946;
17'h7b9f:	data_out=16'h89e3;
17'h7ba0:	data_out=16'h88b0;
17'h7ba1:	data_out=16'ha00;
17'h7ba2:	data_out=16'h89ff;
17'h7ba3:	data_out=16'ha00;
17'h7ba4:	data_out=16'ha00;
17'h7ba5:	data_out=16'h8525;
17'h7ba6:	data_out=16'ha00;
17'h7ba7:	data_out=16'h954;
17'h7ba8:	data_out=16'h9fe;
17'h7ba9:	data_out=16'h8a00;
17'h7baa:	data_out=16'ha00;
17'h7bab:	data_out=16'h8a00;
17'h7bac:	data_out=16'h507;
17'h7bad:	data_out=16'ha00;
17'h7bae:	data_out=16'h476;
17'h7baf:	data_out=16'h89a5;
17'h7bb0:	data_out=16'h966;
17'h7bb1:	data_out=16'h84d;
17'h7bb2:	data_out=16'h9bf;
17'h7bb3:	data_out=16'h89fe;
17'h7bb4:	data_out=16'ha00;
17'h7bb5:	data_out=16'ha00;
17'h7bb6:	data_out=16'ha00;
17'h7bb7:	data_out=16'ha00;
17'h7bb8:	data_out=16'h9ce;
17'h7bb9:	data_out=16'h89fc;
17'h7bba:	data_out=16'h89ff;
17'h7bbb:	data_out=16'h9f7;
17'h7bbc:	data_out=16'h89ec;
17'h7bbd:	data_out=16'ha00;
17'h7bbe:	data_out=16'h9fe;
17'h7bbf:	data_out=16'h89a2;
17'h7bc0:	data_out=16'h87ea;
17'h7bc1:	data_out=16'h86f7;
17'h7bc2:	data_out=16'h642;
17'h7bc3:	data_out=16'h8a00;
17'h7bc4:	data_out=16'h841;
17'h7bc5:	data_out=16'ha00;
17'h7bc6:	data_out=16'ha00;
17'h7bc7:	data_out=16'h80e6;
17'h7bc8:	data_out=16'h887e;
17'h7bc9:	data_out=16'h2c9;
17'h7bca:	data_out=16'h89df;
17'h7bcb:	data_out=16'h892c;
17'h7bcc:	data_out=16'h953;
17'h7bcd:	data_out=16'h8a00;
17'h7bce:	data_out=16'h9fe;
17'h7bcf:	data_out=16'h9fe;
17'h7bd0:	data_out=16'h8a00;
17'h7bd1:	data_out=16'h8746;
17'h7bd2:	data_out=16'ha00;
17'h7bd3:	data_out=16'h893b;
17'h7bd4:	data_out=16'h8801;
17'h7bd5:	data_out=16'h8946;
17'h7bd6:	data_out=16'ha00;
17'h7bd7:	data_out=16'ha00;
17'h7bd8:	data_out=16'h9d5;
17'h7bd9:	data_out=16'h9fc;
17'h7bda:	data_out=16'h89e8;
17'h7bdb:	data_out=16'ha00;
17'h7bdc:	data_out=16'h89da;
17'h7bdd:	data_out=16'h995;
17'h7bde:	data_out=16'h89b6;
17'h7bdf:	data_out=16'ha00;
17'h7be0:	data_out=16'ha00;
17'h7be1:	data_out=16'ha00;
17'h7be2:	data_out=16'h89f6;
17'h7be3:	data_out=16'h89ff;
17'h7be4:	data_out=16'h889b;
17'h7be5:	data_out=16'h8a00;
17'h7be6:	data_out=16'h8a00;
17'h7be7:	data_out=16'h8a00;
17'h7be8:	data_out=16'h9ff;
17'h7be9:	data_out=16'ha00;
17'h7bea:	data_out=16'ha00;
17'h7beb:	data_out=16'h89fb;
17'h7bec:	data_out=16'ha00;
17'h7bed:	data_out=16'h89ff;
17'h7bee:	data_out=16'ha00;
17'h7bef:	data_out=16'h8a00;
17'h7bf0:	data_out=16'ha00;
17'h7bf1:	data_out=16'ha00;
17'h7bf2:	data_out=16'h813;
17'h7bf3:	data_out=16'h9c9;
17'h7bf4:	data_out=16'h9fa;
17'h7bf5:	data_out=16'h421;
17'h7bf6:	data_out=16'h89f6;
17'h7bf7:	data_out=16'h89fb;
17'h7bf8:	data_out=16'h8a00;
17'h7bf9:	data_out=16'ha00;
17'h7bfa:	data_out=16'h89fe;
17'h7bfb:	data_out=16'h9fe;
17'h7bfc:	data_out=16'ha00;
17'h7bfd:	data_out=16'h89fb;
17'h7bfe:	data_out=16'h84e4;
17'h7bff:	data_out=16'h3fb;
17'h7c00:	data_out=16'ha00;
17'h7c01:	data_out=16'ha00;
17'h7c02:	data_out=16'ha00;
17'h7c03:	data_out=16'h89c5;
17'h7c04:	data_out=16'ha00;
17'h7c05:	data_out=16'ha00;
17'h7c06:	data_out=16'h8a00;
17'h7c07:	data_out=16'h89d8;
17'h7c08:	data_out=16'ha00;
17'h7c09:	data_out=16'h8a00;
17'h7c0a:	data_out=16'ha00;
17'h7c0b:	data_out=16'h8a00;
17'h7c0c:	data_out=16'h848a;
17'h7c0d:	data_out=16'ha00;
17'h7c0e:	data_out=16'ha00;
17'h7c0f:	data_out=16'ha00;
17'h7c10:	data_out=16'h8a00;
17'h7c11:	data_out=16'h8e8;
17'h7c12:	data_out=16'ha00;
17'h7c13:	data_out=16'h8358;
17'h7c14:	data_out=16'h89ff;
17'h7c15:	data_out=16'ha00;
17'h7c16:	data_out=16'ha00;
17'h7c17:	data_out=16'h8a00;
17'h7c18:	data_out=16'ha00;
17'h7c19:	data_out=16'h8a00;
17'h7c1a:	data_out=16'ha00;
17'h7c1b:	data_out=16'h8136;
17'h7c1c:	data_out=16'ha00;
17'h7c1d:	data_out=16'h8e5;
17'h7c1e:	data_out=16'h9ff;
17'h7c1f:	data_out=16'h8366;
17'h7c20:	data_out=16'ha00;
17'h7c21:	data_out=16'ha00;
17'h7c22:	data_out=16'h89ff;
17'h7c23:	data_out=16'ha00;
17'h7c24:	data_out=16'ha00;
17'h7c25:	data_out=16'ha00;
17'h7c26:	data_out=16'ha00;
17'h7c27:	data_out=16'h942;
17'h7c28:	data_out=16'ha00;
17'h7c29:	data_out=16'h8a00;
17'h7c2a:	data_out=16'ha00;
17'h7c2b:	data_out=16'h8a00;
17'h7c2c:	data_out=16'ha00;
17'h7c2d:	data_out=16'h89eb;
17'h7c2e:	data_out=16'h9f4;
17'h7c2f:	data_out=16'h86ed;
17'h7c30:	data_out=16'ha00;
17'h7c31:	data_out=16'h84e1;
17'h7c32:	data_out=16'ha00;
17'h7c33:	data_out=16'h89ff;
17'h7c34:	data_out=16'h8146;
17'h7c35:	data_out=16'ha00;
17'h7c36:	data_out=16'ha00;
17'h7c37:	data_out=16'ha00;
17'h7c38:	data_out=16'h63c;
17'h7c39:	data_out=16'h890c;
17'h7c3a:	data_out=16'h89ff;
17'h7c3b:	data_out=16'ha00;
17'h7c3c:	data_out=16'h9ff;
17'h7c3d:	data_out=16'ha00;
17'h7c3e:	data_out=16'ha00;
17'h7c3f:	data_out=16'ha00;
17'h7c40:	data_out=16'ha00;
17'h7c41:	data_out=16'ha00;
17'h7c42:	data_out=16'h69a;
17'h7c43:	data_out=16'h8a00;
17'h7c44:	data_out=16'ha00;
17'h7c45:	data_out=16'ha00;
17'h7c46:	data_out=16'ha00;
17'h7c47:	data_out=16'h2f1;
17'h7c48:	data_out=16'h8946;
17'h7c49:	data_out=16'ha00;
17'h7c4a:	data_out=16'h85c0;
17'h7c4b:	data_out=16'h895c;
17'h7c4c:	data_out=16'ha00;
17'h7c4d:	data_out=16'h8a00;
17'h7c4e:	data_out=16'ha00;
17'h7c4f:	data_out=16'ha00;
17'h7c50:	data_out=16'h89ff;
17'h7c51:	data_out=16'ha00;
17'h7c52:	data_out=16'ha00;
17'h7c53:	data_out=16'h8914;
17'h7c54:	data_out=16'ha00;
17'h7c55:	data_out=16'ha00;
17'h7c56:	data_out=16'ha00;
17'h7c57:	data_out=16'ha00;
17'h7c58:	data_out=16'ha00;
17'h7c59:	data_out=16'ha00;
17'h7c5a:	data_out=16'h89c1;
17'h7c5b:	data_out=16'ha00;
17'h7c5c:	data_out=16'h88c6;
17'h7c5d:	data_out=16'ha00;
17'h7c5e:	data_out=16'h8923;
17'h7c5f:	data_out=16'ha00;
17'h7c60:	data_out=16'ha00;
17'h7c61:	data_out=16'ha00;
17'h7c62:	data_out=16'h89fe;
17'h7c63:	data_out=16'h8a00;
17'h7c64:	data_out=16'h89e9;
17'h7c65:	data_out=16'h8a00;
17'h7c66:	data_out=16'h8a00;
17'h7c67:	data_out=16'h8a00;
17'h7c68:	data_out=16'ha00;
17'h7c69:	data_out=16'ha00;
17'h7c6a:	data_out=16'ha00;
17'h7c6b:	data_out=16'h7cf;
17'h7c6c:	data_out=16'ha00;
17'h7c6d:	data_out=16'h89ff;
17'h7c6e:	data_out=16'ha00;
17'h7c6f:	data_out=16'h89fb;
17'h7c70:	data_out=16'ha00;
17'h7c71:	data_out=16'ha00;
17'h7c72:	data_out=16'ha00;
17'h7c73:	data_out=16'ha00;
17'h7c74:	data_out=16'ha00;
17'h7c75:	data_out=16'ha00;
17'h7c76:	data_out=16'h8a00;
17'h7c77:	data_out=16'h9f3;
17'h7c78:	data_out=16'h8a00;
17'h7c79:	data_out=16'ha00;
17'h7c7a:	data_out=16'h89ff;
17'h7c7b:	data_out=16'ha00;
17'h7c7c:	data_out=16'ha00;
17'h7c7d:	data_out=16'h89fd;
17'h7c7e:	data_out=16'h88a9;
17'h7c7f:	data_out=16'h9fe;
17'h7c80:	data_out=16'ha00;
17'h7c81:	data_out=16'ha00;
17'h7c82:	data_out=16'ha00;
17'h7c83:	data_out=16'h9e6;
17'h7c84:	data_out=16'ha00;
17'h7c85:	data_out=16'ha00;
17'h7c86:	data_out=16'hf8;
17'h7c87:	data_out=16'h51b;
17'h7c88:	data_out=16'ha00;
17'h7c89:	data_out=16'h884d;
17'h7c8a:	data_out=16'ha00;
17'h7c8b:	data_out=16'h8a00;
17'h7c8c:	data_out=16'h4a6;
17'h7c8d:	data_out=16'ha00;
17'h7c8e:	data_out=16'ha00;
17'h7c8f:	data_out=16'ha00;
17'h7c90:	data_out=16'h84df;
17'h7c91:	data_out=16'ha00;
17'h7c92:	data_out=16'h3bc;
17'h7c93:	data_out=16'h9cc;
17'h7c94:	data_out=16'h68e;
17'h7c95:	data_out=16'ha00;
17'h7c96:	data_out=16'ha00;
17'h7c97:	data_out=16'h88d8;
17'h7c98:	data_out=16'ha00;
17'h7c99:	data_out=16'h8a00;
17'h7c9a:	data_out=16'ha00;
17'h7c9b:	data_out=16'h6a2;
17'h7c9c:	data_out=16'ha00;
17'h7c9d:	data_out=16'h8fc;
17'h7c9e:	data_out=16'ha00;
17'h7c9f:	data_out=16'h9df;
17'h7ca0:	data_out=16'ha00;
17'h7ca1:	data_out=16'ha00;
17'h7ca2:	data_out=16'h89ff;
17'h7ca3:	data_out=16'ha00;
17'h7ca4:	data_out=16'ha00;
17'h7ca5:	data_out=16'ha00;
17'h7ca6:	data_out=16'ha00;
17'h7ca7:	data_out=16'ha00;
17'h7ca8:	data_out=16'ha00;
17'h7ca9:	data_out=16'h8a00;
17'h7caa:	data_out=16'ha00;
17'h7cab:	data_out=16'h8a00;
17'h7cac:	data_out=16'ha00;
17'h7cad:	data_out=16'h8a00;
17'h7cae:	data_out=16'h9df;
17'h7caf:	data_out=16'ha00;
17'h7cb0:	data_out=16'ha00;
17'h7cb1:	data_out=16'h8379;
17'h7cb2:	data_out=16'ha00;
17'h7cb3:	data_out=16'h75d;
17'h7cb4:	data_out=16'h8173;
17'h7cb5:	data_out=16'ha00;
17'h7cb6:	data_out=16'ha00;
17'h7cb7:	data_out=16'ha00;
17'h7cb8:	data_out=16'h611;
17'h7cb9:	data_out=16'h9e7;
17'h7cba:	data_out=16'h8764;
17'h7cbb:	data_out=16'ha00;
17'h7cbc:	data_out=16'h9ff;
17'h7cbd:	data_out=16'ha00;
17'h7cbe:	data_out=16'ha00;
17'h7cbf:	data_out=16'ha00;
17'h7cc0:	data_out=16'ha00;
17'h7cc1:	data_out=16'ha00;
17'h7cc2:	data_out=16'h83ed;
17'h7cc3:	data_out=16'h8a00;
17'h7cc4:	data_out=16'ha00;
17'h7cc5:	data_out=16'ha00;
17'h7cc6:	data_out=16'ha00;
17'h7cc7:	data_out=16'h9a2;
17'h7cc8:	data_out=16'h8684;
17'h7cc9:	data_out=16'ha00;
17'h7cca:	data_out=16'h7eb;
17'h7ccb:	data_out=16'h89dc;
17'h7ccc:	data_out=16'ha00;
17'h7ccd:	data_out=16'h89ff;
17'h7cce:	data_out=16'ha00;
17'h7ccf:	data_out=16'ha00;
17'h7cd0:	data_out=16'h6e1;
17'h7cd1:	data_out=16'ha00;
17'h7cd2:	data_out=16'ha00;
17'h7cd3:	data_out=16'ha00;
17'h7cd4:	data_out=16'ha00;
17'h7cd5:	data_out=16'ha00;
17'h7cd6:	data_out=16'ha00;
17'h7cd7:	data_out=16'ha00;
17'h7cd8:	data_out=16'ha00;
17'h7cd9:	data_out=16'ha00;
17'h7cda:	data_out=16'h89cd;
17'h7cdb:	data_out=16'ha00;
17'h7cdc:	data_out=16'h961;
17'h7cdd:	data_out=16'ha00;
17'h7cde:	data_out=16'h9fe;
17'h7cdf:	data_out=16'ha00;
17'h7ce0:	data_out=16'ha00;
17'h7ce1:	data_out=16'ha00;
17'h7ce2:	data_out=16'h89ff;
17'h7ce3:	data_out=16'h674;
17'h7ce4:	data_out=16'h89f9;
17'h7ce5:	data_out=16'h8a00;
17'h7ce6:	data_out=16'h8a00;
17'h7ce7:	data_out=16'h8a00;
17'h7ce8:	data_out=16'ha00;
17'h7ce9:	data_out=16'ha00;
17'h7cea:	data_out=16'ha00;
17'h7ceb:	data_out=16'ha00;
17'h7cec:	data_out=16'ha00;
17'h7ced:	data_out=16'h6fe;
17'h7cee:	data_out=16'ha00;
17'h7cef:	data_out=16'h98e;
17'h7cf0:	data_out=16'ha00;
17'h7cf1:	data_out=16'ha00;
17'h7cf2:	data_out=16'ha00;
17'h7cf3:	data_out=16'ha00;
17'h7cf4:	data_out=16'ha00;
17'h7cf5:	data_out=16'ha00;
17'h7cf6:	data_out=16'h8a00;
17'h7cf7:	data_out=16'h9fc;
17'h7cf8:	data_out=16'h8a00;
17'h7cf9:	data_out=16'ha00;
17'h7cfa:	data_out=16'h96a;
17'h7cfb:	data_out=16'ha00;
17'h7cfc:	data_out=16'ha00;
17'h7cfd:	data_out=16'h7a9;
17'h7cfe:	data_out=16'h8420;
17'h7cff:	data_out=16'ha00;
17'h7d00:	data_out=16'h9b7;
17'h7d01:	data_out=16'ha00;
17'h7d02:	data_out=16'ha00;
17'h7d03:	data_out=16'h48d;
17'h7d04:	data_out=16'ha00;
17'h7d05:	data_out=16'ha00;
17'h7d06:	data_out=16'h501;
17'h7d07:	data_out=16'h8a;
17'h7d08:	data_out=16'h9ff;
17'h7d09:	data_out=16'h8a00;
17'h7d0a:	data_out=16'ha00;
17'h7d0b:	data_out=16'h8a00;
17'h7d0c:	data_out=16'h822;
17'h7d0d:	data_out=16'h50f;
17'h7d0e:	data_out=16'h7e9;
17'h7d0f:	data_out=16'h9ff;
17'h7d10:	data_out=16'h8336;
17'h7d11:	data_out=16'ha00;
17'h7d12:	data_out=16'h84d2;
17'h7d13:	data_out=16'h3f4;
17'h7d14:	data_out=16'h2ac;
17'h7d15:	data_out=16'ha00;
17'h7d16:	data_out=16'h9ff;
17'h7d17:	data_out=16'h8311;
17'h7d18:	data_out=16'ha00;
17'h7d19:	data_out=16'h8a00;
17'h7d1a:	data_out=16'ha00;
17'h7d1b:	data_out=16'h8758;
17'h7d1c:	data_out=16'ha00;
17'h7d1d:	data_out=16'ha00;
17'h7d1e:	data_out=16'h6a2;
17'h7d1f:	data_out=16'h9de;
17'h7d20:	data_out=16'h9ff;
17'h7d21:	data_out=16'h7be;
17'h7d22:	data_out=16'h89e4;
17'h7d23:	data_out=16'h922;
17'h7d24:	data_out=16'h92b;
17'h7d25:	data_out=16'h8104;
17'h7d26:	data_out=16'he5;
17'h7d27:	data_out=16'h98c;
17'h7d28:	data_out=16'h78b;
17'h7d29:	data_out=16'h8525;
17'h7d2a:	data_out=16'h69a;
17'h7d2b:	data_out=16'h8a00;
17'h7d2c:	data_out=16'h9ff;
17'h7d2d:	data_out=16'h8a00;
17'h7d2e:	data_out=16'h9d0;
17'h7d2f:	data_out=16'h27d;
17'h7d30:	data_out=16'ha00;
17'h7d31:	data_out=16'h806c;
17'h7d32:	data_out=16'ha00;
17'h7d33:	data_out=16'h438;
17'h7d34:	data_out=16'h282;
17'h7d35:	data_out=16'h9ff;
17'h7d36:	data_out=16'h9ff;
17'h7d37:	data_out=16'ha00;
17'h7d38:	data_out=16'h9fb;
17'h7d39:	data_out=16'h58f;
17'h7d3a:	data_out=16'h8993;
17'h7d3b:	data_out=16'h9fd;
17'h7d3c:	data_out=16'ha00;
17'h7d3d:	data_out=16'ha00;
17'h7d3e:	data_out=16'h78b;
17'h7d3f:	data_out=16'ha00;
17'h7d40:	data_out=16'ha00;
17'h7d41:	data_out=16'h9ff;
17'h7d42:	data_out=16'h8058;
17'h7d43:	data_out=16'h9a;
17'h7d44:	data_out=16'h9fe;
17'h7d45:	data_out=16'ha00;
17'h7d46:	data_out=16'h8464;
17'h7d47:	data_out=16'h844a;
17'h7d48:	data_out=16'h86fd;
17'h7d49:	data_out=16'h8036;
17'h7d4a:	data_out=16'h8f1;
17'h7d4b:	data_out=16'h8899;
17'h7d4c:	data_out=16'h2b2;
17'h7d4d:	data_out=16'h89ea;
17'h7d4e:	data_out=16'ha00;
17'h7d4f:	data_out=16'h2da;
17'h7d50:	data_out=16'h9f5;
17'h7d51:	data_out=16'ha00;
17'h7d52:	data_out=16'ha00;
17'h7d53:	data_out=16'h809c;
17'h7d54:	data_out=16'h9ff;
17'h7d55:	data_out=16'h9fc;
17'h7d56:	data_out=16'ha00;
17'h7d57:	data_out=16'ha00;
17'h7d58:	data_out=16'ha00;
17'h7d59:	data_out=16'ha00;
17'h7d5a:	data_out=16'h86d3;
17'h7d5b:	data_out=16'ha00;
17'h7d5c:	data_out=16'h805;
17'h7d5d:	data_out=16'ha00;
17'h7d5e:	data_out=16'h1b0;
17'h7d5f:	data_out=16'h564;
17'h7d60:	data_out=16'h31a;
17'h7d61:	data_out=16'ha00;
17'h7d62:	data_out=16'h8643;
17'h7d63:	data_out=16'h3ab;
17'h7d64:	data_out=16'h85d2;
17'h7d65:	data_out=16'h8a00;
17'h7d66:	data_out=16'h8a00;
17'h7d67:	data_out=16'h8a00;
17'h7d68:	data_out=16'h7a1;
17'h7d69:	data_out=16'h9fd;
17'h7d6a:	data_out=16'h80a;
17'h7d6b:	data_out=16'h9fe;
17'h7d6c:	data_out=16'ha00;
17'h7d6d:	data_out=16'h3f2;
17'h7d6e:	data_out=16'h80a;
17'h7d6f:	data_out=16'h97c;
17'h7d70:	data_out=16'h7fa;
17'h7d71:	data_out=16'h9fe;
17'h7d72:	data_out=16'ha00;
17'h7d73:	data_out=16'ha00;
17'h7d74:	data_out=16'ha00;
17'h7d75:	data_out=16'ha00;
17'h7d76:	data_out=16'h8a00;
17'h7d77:	data_out=16'h9ff;
17'h7d78:	data_out=16'h12;
17'h7d79:	data_out=16'ha00;
17'h7d7a:	data_out=16'h344;
17'h7d7b:	data_out=16'h78b;
17'h7d7c:	data_out=16'h85c;
17'h7d7d:	data_out=16'h604;
17'h7d7e:	data_out=16'h880b;
17'h7d7f:	data_out=16'ha00;
17'h7d80:	data_out=16'h80f8;
17'h7d81:	data_out=16'h12c;
17'h7d82:	data_out=16'h7d;
17'h7d83:	data_out=16'h8192;
17'h7d84:	data_out=16'h12b;
17'h7d85:	data_out=16'h8;
17'h7d86:	data_out=16'h1a;
17'h7d87:	data_out=16'h83d3;
17'h7d88:	data_out=16'h80bc;
17'h7d89:	data_out=16'h8562;
17'h7d8a:	data_out=16'h171;
17'h7d8b:	data_out=16'h85ba;
17'h7d8c:	data_out=16'h8205;
17'h7d8d:	data_out=16'h8236;
17'h7d8e:	data_out=16'h134;
17'h7d8f:	data_out=16'h47;
17'h7d90:	data_out=16'h83d9;
17'h7d91:	data_out=16'h8040;
17'h7d92:	data_out=16'h8381;
17'h7d93:	data_out=16'h825f;
17'h7d94:	data_out=16'h821e;
17'h7d95:	data_out=16'hb5;
17'h7d96:	data_out=16'h80ba;
17'h7d97:	data_out=16'h82d0;
17'h7d98:	data_out=16'h8010;
17'h7d99:	data_out=16'h8291;
17'h7d9a:	data_out=16'h103;
17'h7d9b:	data_out=16'h8495;
17'h7d9c:	data_out=16'h132;
17'h7d9d:	data_out=16'h81fd;
17'h7d9e:	data_out=16'h825f;
17'h7d9f:	data_out=16'h13;
17'h7da0:	data_out=16'h82f2;
17'h7da1:	data_out=16'h118;
17'h7da2:	data_out=16'h8355;
17'h7da3:	data_out=16'h1d1;
17'h7da4:	data_out=16'h1d1;
17'h7da5:	data_out=16'h8383;
17'h7da6:	data_out=16'h8398;
17'h7da7:	data_out=16'h82f9;
17'h7da8:	data_out=16'hf8;
17'h7da9:	data_out=16'h81dc;
17'h7daa:	data_out=16'h8317;
17'h7dab:	data_out=16'h8592;
17'h7dac:	data_out=16'h80da;
17'h7dad:	data_out=16'h22;
17'h7dae:	data_out=16'h826e;
17'h7daf:	data_out=16'h82ad;
17'h7db0:	data_out=16'h139;
17'h7db1:	data_out=16'h8153;
17'h7db2:	data_out=16'h136;
17'h7db3:	data_out=16'h8252;
17'h7db4:	data_out=16'h80af;
17'h7db5:	data_out=16'h8109;
17'h7db6:	data_out=16'h810b;
17'h7db7:	data_out=16'h3a;
17'h7db8:	data_out=16'h47e;
17'h7db9:	data_out=16'h8227;
17'h7dba:	data_out=16'h83ee;
17'h7dbb:	data_out=16'h80d7;
17'h7dbc:	data_out=16'h8048;
17'h7dbd:	data_out=16'h81e3;
17'h7dbe:	data_out=16'hf3;
17'h7dbf:	data_out=16'h76;
17'h7dc0:	data_out=16'h80;
17'h7dc1:	data_out=16'h8176;
17'h7dc2:	data_out=16'h81e4;
17'h7dc3:	data_out=16'h80b5;
17'h7dc4:	data_out=16'h81de;
17'h7dc5:	data_out=16'h30;
17'h7dc6:	data_out=16'h80e0;
17'h7dc7:	data_out=16'h837e;
17'h7dc8:	data_out=16'h83bd;
17'h7dc9:	data_out=16'h831c;
17'h7dca:	data_out=16'h8249;
17'h7dcb:	data_out=16'h837a;
17'h7dcc:	data_out=16'h8250;
17'h7dcd:	data_out=16'h835a;
17'h7dce:	data_out=16'h8274;
17'h7dcf:	data_out=16'h82cd;
17'h7dd0:	data_out=16'he3;
17'h7dd1:	data_out=16'h184;
17'h7dd2:	data_out=16'h225;
17'h7dd3:	data_out=16'h8439;
17'h7dd4:	data_out=16'h8169;
17'h7dd5:	data_out=16'h6e;
17'h7dd6:	data_out=16'h60;
17'h7dd7:	data_out=16'h110;
17'h7dd8:	data_out=16'h150;
17'h7dd9:	data_out=16'hfb;
17'h7dda:	data_out=16'h8241;
17'h7ddb:	data_out=16'h5f7;
17'h7ddc:	data_out=16'h814f;
17'h7ddd:	data_out=16'h80ef;
17'h7dde:	data_out=16'h831f;
17'h7ddf:	data_out=16'h80c5;
17'h7de0:	data_out=16'h811a;
17'h7de1:	data_out=16'h1c1;
17'h7de2:	data_out=16'h823e;
17'h7de3:	data_out=16'h8268;
17'h7de4:	data_out=16'h82f1;
17'h7de5:	data_out=16'h846a;
17'h7de6:	data_out=16'h8490;
17'h7de7:	data_out=16'h838f;
17'h7de8:	data_out=16'h112;
17'h7de9:	data_out=16'h801d;
17'h7dea:	data_out=16'h14d;
17'h7deb:	data_out=16'h8064;
17'h7dec:	data_out=16'h76;
17'h7ded:	data_out=16'h8262;
17'h7dee:	data_out=16'h146;
17'h7def:	data_out=16'h8111;
17'h7df0:	data_out=16'h131;
17'h7df1:	data_out=16'h81d0;
17'h7df2:	data_out=16'h241;
17'h7df3:	data_out=16'hf3;
17'h7df4:	data_out=16'h145;
17'h7df5:	data_out=16'h39d;
17'h7df6:	data_out=16'h8612;
17'h7df7:	data_out=16'h80de;
17'h7df8:	data_out=16'h8197;
17'h7df9:	data_out=16'h8263;
17'h7dfa:	data_out=16'h825c;
17'h7dfb:	data_out=16'hf4;
17'h7dfc:	data_out=16'ha2;
17'h7dfd:	data_out=16'h809e;
17'h7dfe:	data_out=16'h84e4;
17'h7dff:	data_out=16'h36;
17'h7e00:	data_out=16'h3a;
17'h7e01:	data_out=16'h6c;
17'h7e02:	data_out=16'h61;
17'h7e03:	data_out=16'h52;
17'h7e04:	data_out=16'h5d;
17'h7e05:	data_out=16'h66;
17'h7e06:	data_out=16'h8010;
17'h7e07:	data_out=16'h4d;
17'h7e08:	data_out=16'h34;
17'h7e09:	data_out=16'h8013;
17'h7e0a:	data_out=16'h8a;
17'h7e0b:	data_out=16'h8009;
17'h7e0c:	data_out=16'h71;
17'h7e0d:	data_out=16'h33;
17'h7e0e:	data_out=16'h6;
17'h7e0f:	data_out=16'h48;
17'h7e10:	data_out=16'h3;
17'h7e11:	data_out=16'h63;
17'h7e12:	data_out=16'h4a;
17'h7e13:	data_out=16'h22;
17'h7e14:	data_out=16'h63;
17'h7e15:	data_out=16'h2a;
17'h7e16:	data_out=16'h40;
17'h7e17:	data_out=16'h65;
17'h7e18:	data_out=16'h6;
17'h7e19:	data_out=16'h11;
17'h7e1a:	data_out=16'h53;
17'h7e1b:	data_out=16'h2c;
17'h7e1c:	data_out=16'h8c;
17'h7e1d:	data_out=16'hbe;
17'h7e1e:	data_out=16'h69;
17'h7e1f:	data_out=16'h2e;
17'h7e20:	data_out=16'ha0;
17'h7e21:	data_out=16'h10;
17'h7e22:	data_out=16'h45;
17'h7e23:	data_out=16'hd;
17'h7e24:	data_out=16'hc;
17'h7e25:	data_out=16'h3d;
17'h7e26:	data_out=16'h8010;
17'h7e27:	data_out=16'hae;
17'h7e28:	data_out=16'h8001;
17'h7e29:	data_out=16'h2d;
17'h7e2a:	data_out=16'h1d;
17'h7e2b:	data_out=16'h39;
17'h7e2c:	data_out=16'h58;
17'h7e2d:	data_out=16'h2e;
17'h7e2e:	data_out=16'h2c;
17'h7e2f:	data_out=16'h6b;
17'h7e30:	data_out=16'h6f;
17'h7e31:	data_out=16'h69;
17'h7e32:	data_out=16'h69;
17'h7e33:	data_out=16'h67;
17'h7e34:	data_out=16'h38;
17'h7e35:	data_out=16'h66;
17'h7e36:	data_out=16'h33;
17'h7e37:	data_out=16'h7e;
17'h7e38:	data_out=16'h41;
17'h7e39:	data_out=16'h23;
17'h7e3a:	data_out=16'h66;
17'h7e3b:	data_out=16'h3b;
17'h7e3c:	data_out=16'h71;
17'h7e3d:	data_out=16'h3a;
17'h7e3e:	data_out=16'h11;
17'h7e3f:	data_out=16'h4a;
17'h7e40:	data_out=16'h61;
17'h7e41:	data_out=16'h4f;
17'h7e42:	data_out=16'h38;
17'h7e43:	data_out=16'h800b;
17'h7e44:	data_out=16'h42;
17'h7e45:	data_out=16'hf;
17'h7e46:	data_out=16'h66;
17'h7e47:	data_out=16'h4c;
17'h7e48:	data_out=16'h17;
17'h7e49:	data_out=16'h4e;
17'h7e4a:	data_out=16'h43;
17'h7e4b:	data_out=16'h7a;
17'h7e4c:	data_out=16'h49;
17'h7e4d:	data_out=16'h58;
17'h7e4e:	data_out=16'h56;
17'h7e4f:	data_out=16'h47;
17'h7e50:	data_out=16'h5d;
17'h7e51:	data_out=16'h2d;
17'h7e52:	data_out=16'hd;
17'h7e53:	data_out=16'hca;
17'h7e54:	data_out=16'h6f;
17'h7e55:	data_out=16'h21;
17'h7e56:	data_out=16'h57;
17'h7e57:	data_out=16'h3b;
17'h7e58:	data_out=16'h5e;
17'h7e59:	data_out=16'h41;
17'h7e5a:	data_out=16'h34;
17'h7e5b:	data_out=16'h49;
17'h7e5c:	data_out=16'h6d;
17'h7e5d:	data_out=16'h51;
17'h7e5e:	data_out=16'h67;
17'h7e5f:	data_out=16'h1d;
17'h7e60:	data_out=16'h1d;
17'h7e61:	data_out=16'h64;
17'h7e62:	data_out=16'h29;
17'h7e63:	data_out=16'h68;
17'h7e64:	data_out=16'h36;
17'h7e65:	data_out=16'h59;
17'h7e66:	data_out=16'h1e;
17'h7e67:	data_out=16'h29;
17'h7e68:	data_out=16'hf;
17'h7e69:	data_out=16'h47;
17'h7e6a:	data_out=16'h3;
17'h7e6b:	data_out=16'h5e;
17'h7e6c:	data_out=16'hd2;
17'h7e6d:	data_out=16'h68;
17'h7e6e:	data_out=16'h6;
17'h7e6f:	data_out=16'h7e;
17'h7e70:	data_out=16'h6;
17'h7e71:	data_out=16'h1b;
17'h7e72:	data_out=16'h4f;
17'h7e73:	data_out=16'h55;
17'h7e74:	data_out=16'h69;
17'h7e75:	data_out=16'h36;
17'h7e76:	data_out=16'h22;
17'h7e77:	data_out=16'h14;
17'h7e78:	data_out=16'h800f;
17'h7e79:	data_out=16'h3e;
17'h7e7a:	data_out=16'h63;
17'h7e7b:	data_out=16'h8000;
17'h7e7c:	data_out=16'h17;
17'h7e7d:	data_out=16'h8016;
17'h7e7e:	data_out=16'h801d;
17'h7e7f:	data_out=16'h3b;
17'h7e80:	data_out=16'h4e8;
17'h7e81:	data_out=16'h623;
17'h7e82:	data_out=16'h23a;
17'h7e83:	data_out=16'h32a;
17'h7e84:	data_out=16'h806a;
17'h7e85:	data_out=16'h7;
17'h7e86:	data_out=16'h82c8;
17'h7e87:	data_out=16'h1a4;
17'h7e88:	data_out=16'h30b;
17'h7e89:	data_out=16'h1a;
17'h7e8a:	data_out=16'h2c6;
17'h7e8b:	data_out=16'h44;
17'h7e8c:	data_out=16'h8006;
17'h7e8d:	data_out=16'h326;
17'h7e8e:	data_out=16'h11;
17'h7e8f:	data_out=16'h389;
17'h7e90:	data_out=16'h2a1;
17'h7e91:	data_out=16'h80a7;
17'h7e92:	data_out=16'h38b;
17'h7e93:	data_out=16'h2a6;
17'h7e94:	data_out=16'h232;
17'h7e95:	data_out=16'hef;
17'h7e96:	data_out=16'h1e7;
17'h7e97:	data_out=16'h2fd;
17'h7e98:	data_out=16'h80;
17'h7e99:	data_out=16'h8141;
17'h7e9a:	data_out=16'h80b4;
17'h7e9b:	data_out=16'h412;
17'h7e9c:	data_out=16'h800c;
17'h7e9d:	data_out=16'h515;
17'h7e9e:	data_out=16'h3d6;
17'h7e9f:	data_out=16'h8221;
17'h7ea0:	data_out=16'h775;
17'h7ea1:	data_out=16'hd;
17'h7ea2:	data_out=16'h400;
17'h7ea3:	data_out=16'h8094;
17'h7ea4:	data_out=16'h8086;
17'h7ea5:	data_out=16'h224;
17'h7ea6:	data_out=16'h80d2;
17'h7ea7:	data_out=16'h52f;
17'h7ea8:	data_out=16'h1a;
17'h7ea9:	data_out=16'h406;
17'h7eaa:	data_out=16'h5c2;
17'h7eab:	data_out=16'h131;
17'h7eac:	data_out=16'h166;
17'h7ead:	data_out=16'h590;
17'h7eae:	data_out=16'h4d2;
17'h7eaf:	data_out=16'h820;
17'h7eb0:	data_out=16'h8036;
17'h7eb1:	data_out=16'h266;
17'h7eb2:	data_out=16'h8017;
17'h7eb3:	data_out=16'h285;
17'h7eb4:	data_out=16'h25c;
17'h7eb5:	data_out=16'h80aa;
17'h7eb6:	data_out=16'h596;
17'h7eb7:	data_out=16'h231;
17'h7eb8:	data_out=16'h80a1;
17'h7eb9:	data_out=16'h2f2;
17'h7eba:	data_out=16'h5f7;
17'h7ebb:	data_out=16'h80a8;
17'h7ebc:	data_out=16'h3e1;
17'h7ebd:	data_out=16'h154;
17'h7ebe:	data_out=16'h14;
17'h7ebf:	data_out=16'h808d;
17'h7ec0:	data_out=16'h800a;
17'h7ec1:	data_out=16'h1ef;
17'h7ec2:	data_out=16'h6ba;
17'h7ec3:	data_out=16'h83cb;
17'h7ec4:	data_out=16'h803c;
17'h7ec5:	data_out=16'h804a;
17'h7ec6:	data_out=16'h2f7;
17'h7ec7:	data_out=16'h2d3;
17'h7ec8:	data_out=16'h3af;
17'h7ec9:	data_out=16'h1af;
17'h7eca:	data_out=16'h2c6;
17'h7ecb:	data_out=16'h692;
17'h7ecc:	data_out=16'h4e5;
17'h7ecd:	data_out=16'h458;
17'h7ece:	data_out=16'h54a;
17'h7ecf:	data_out=16'h40c;
17'h7ed0:	data_out=16'h810a;
17'h7ed1:	data_out=16'h8088;
17'h7ed2:	data_out=16'h80aa;
17'h7ed3:	data_out=16'h6ce;
17'h7ed4:	data_out=16'h86a;
17'h7ed5:	data_out=16'ha;
17'h7ed6:	data_out=16'h5d;
17'h7ed7:	data_out=16'h70;
17'h7ed8:	data_out=16'hf3;
17'h7ed9:	data_out=16'hd9;
17'h7eda:	data_out=16'h347;
17'h7edb:	data_out=16'h8215;
17'h7edc:	data_out=16'h30a;
17'h7edd:	data_out=16'h6a0;
17'h7ede:	data_out=16'h802;
17'h7edf:	data_out=16'h3a8;
17'h7ee0:	data_out=16'h14d;
17'h7ee1:	data_out=16'h80b7;
17'h7ee2:	data_out=16'h138;
17'h7ee3:	data_out=16'h281;
17'h7ee4:	data_out=16'h9e;
17'h7ee5:	data_out=16'h139;
17'h7ee6:	data_out=16'h8153;
17'h7ee7:	data_out=16'h2b4;
17'h7ee8:	data_out=16'ha;
17'h7ee9:	data_out=16'h36b;
17'h7eea:	data_out=16'h8007;
17'h7eeb:	data_out=16'h806c;
17'h7eec:	data_out=16'ha00;
17'h7eed:	data_out=16'h297;
17'h7eee:	data_out=16'h8007;
17'h7eef:	data_out=16'h1fa;
17'h7ef0:	data_out=16'h3;
17'h7ef1:	data_out=16'h1b6;
17'h7ef2:	data_out=16'h8046;
17'h7ef3:	data_out=16'h55;
17'h7ef4:	data_out=16'h8036;
17'h7ef5:	data_out=16'h82bf;
17'h7ef6:	data_out=16'h58;
17'h7ef7:	data_out=16'h810d;
17'h7ef8:	data_out=16'h83a9;
17'h7ef9:	data_out=16'h564;
17'h7efa:	data_out=16'h26a;
17'h7efb:	data_out=16'h12;
17'h7efc:	data_out=16'h140;
17'h7efd:	data_out=16'h8372;
17'h7efe:	data_out=16'h816a;
17'h7eff:	data_out=16'h805c;
17'h7f00:	data_out=16'ha00;
17'h7f01:	data_out=16'ha00;
17'h7f02:	data_out=16'h6d2;
17'h7f03:	data_out=16'ha00;
17'h7f04:	data_out=16'h528;
17'h7f05:	data_out=16'h783;
17'h7f06:	data_out=16'h8236;
17'h7f07:	data_out=16'ha00;
17'h7f08:	data_out=16'h823;
17'h7f09:	data_out=16'h54e;
17'h7f0a:	data_out=16'h9fa;
17'h7f0b:	data_out=16'h3a1;
17'h7f0c:	data_out=16'h2c5;
17'h7f0d:	data_out=16'h882;
17'h7f0e:	data_out=16'h53;
17'h7f0f:	data_out=16'ha00;
17'h7f10:	data_out=16'h91d;
17'h7f11:	data_out=16'h5ac;
17'h7f12:	data_out=16'ha00;
17'h7f13:	data_out=16'ha00;
17'h7f14:	data_out=16'h6e0;
17'h7f15:	data_out=16'h2a1;
17'h7f16:	data_out=16'h7ae;
17'h7f17:	data_out=16'h869;
17'h7f18:	data_out=16'he4;
17'h7f19:	data_out=16'h60;
17'h7f1a:	data_out=16'h55f;
17'h7f1b:	data_out=16'h9ff;
17'h7f1c:	data_out=16'h4e9;
17'h7f1d:	data_out=16'ha00;
17'h7f1e:	data_out=16'ha00;
17'h7f1f:	data_out=16'h94;
17'h7f20:	data_out=16'ha00;
17'h7f21:	data_out=16'h56;
17'h7f22:	data_out=16'ha00;
17'h7f23:	data_out=16'h84e1;
17'h7f24:	data_out=16'h84e2;
17'h7f25:	data_out=16'h8bd;
17'h7f26:	data_out=16'h224;
17'h7f27:	data_out=16'ha00;
17'h7f28:	data_out=16'h5f;
17'h7f29:	data_out=16'ha00;
17'h7f2a:	data_out=16'ha00;
17'h7f2b:	data_out=16'h611;
17'h7f2c:	data_out=16'h611;
17'h7f2d:	data_out=16'ha00;
17'h7f2e:	data_out=16'ha00;
17'h7f2f:	data_out=16'ha00;
17'h7f30:	data_out=16'h4bb;
17'h7f31:	data_out=16'h9fc;
17'h7f32:	data_out=16'h57e;
17'h7f33:	data_out=16'h89b;
17'h7f34:	data_out=16'h72e;
17'h7f35:	data_out=16'h64b;
17'h7f36:	data_out=16'ha00;
17'h7f37:	data_out=16'h6d5;
17'h7f38:	data_out=16'h45c;
17'h7f39:	data_out=16'h98b;
17'h7f3a:	data_out=16'ha00;
17'h7f3b:	data_out=16'h4b2;
17'h7f3c:	data_out=16'h930;
17'h7f3d:	data_out=16'ha00;
17'h7f3e:	data_out=16'h5f;
17'h7f3f:	data_out=16'h77e;
17'h7f40:	data_out=16'h6cf;
17'h7f41:	data_out=16'h216;
17'h7f42:	data_out=16'ha00;
17'h7f43:	data_out=16'h85ce;
17'h7f44:	data_out=16'h744;
17'h7f45:	data_out=16'h2ce;
17'h7f46:	data_out=16'h52c;
17'h7f47:	data_out=16'ha00;
17'h7f48:	data_out=16'ha00;
17'h7f49:	data_out=16'h835;
17'h7f4a:	data_out=16'ha00;
17'h7f4b:	data_out=16'ha00;
17'h7f4c:	data_out=16'h9fe;
17'h7f4d:	data_out=16'ha00;
17'h7f4e:	data_out=16'ha00;
17'h7f4f:	data_out=16'h9ff;
17'h7f50:	data_out=16'h13c;
17'h7f51:	data_out=16'h80f6;
17'h7f52:	data_out=16'h8539;
17'h7f53:	data_out=16'ha00;
17'h7f54:	data_out=16'ha00;
17'h7f55:	data_out=16'h8050;
17'h7f56:	data_out=16'h5c0;
17'h7f57:	data_out=16'h64d;
17'h7f58:	data_out=16'h29e;
17'h7f59:	data_out=16'h904;
17'h7f5a:	data_out=16'h9ff;
17'h7f5b:	data_out=16'he4;
17'h7f5c:	data_out=16'h9fd;
17'h7f5d:	data_out=16'ha00;
17'h7f5e:	data_out=16'ha00;
17'h7f5f:	data_out=16'h8ea;
17'h7f60:	data_out=16'h402;
17'h7f61:	data_out=16'h4a0;
17'h7f62:	data_out=16'h30c;
17'h7f63:	data_out=16'h870;
17'h7f64:	data_out=16'h508;
17'h7f65:	data_out=16'h9fe;
17'h7f66:	data_out=16'h802a;
17'h7f67:	data_out=16'h7cb;
17'h7f68:	data_out=16'h57;
17'h7f69:	data_out=16'h6d4;
17'h7f6a:	data_out=16'h4e;
17'h7f6b:	data_out=16'h6b3;
17'h7f6c:	data_out=16'ha00;
17'h7f6d:	data_out=16'h8be;
17'h7f6e:	data_out=16'h4f;
17'h7f6f:	data_out=16'h9ff;
17'h7f70:	data_out=16'h51;
17'h7f71:	data_out=16'h6c8;
17'h7f72:	data_out=16'h74f;
17'h7f73:	data_out=16'h936;
17'h7f74:	data_out=16'h4a2;
17'h7f75:	data_out=16'h8310;
17'h7f76:	data_out=16'h266;
17'h7f77:	data_out=16'hd6;
17'h7f78:	data_out=16'h8506;
17'h7f79:	data_out=16'h9ff;
17'h7f7a:	data_out=16'h7ab;
17'h7f7b:	data_out=16'h60;
17'h7f7c:	data_out=16'h2fc;
17'h7f7d:	data_out=16'h820d;
17'h7f7e:	data_out=16'h33d;
17'h7f7f:	data_out=16'h574;
17'h7f80:	data_out=16'h329;
17'h7f81:	data_out=16'ha00;
17'h7f82:	data_out=16'h9f4;
17'h7f83:	data_out=16'h99e;
17'h7f84:	data_out=16'h8677;
17'h7f85:	data_out=16'h9f8;
17'h7f86:	data_out=16'h85ab;
17'h7f87:	data_out=16'h2a9;
17'h7f88:	data_out=16'h975;
17'h7f89:	data_out=16'h8948;
17'h7f8a:	data_out=16'h5b9;
17'h7f8b:	data_out=16'ha00;
17'h7f8c:	data_out=16'h17d;
17'h7f8d:	data_out=16'h6fd;
17'h7f8e:	data_out=16'h82ba;
17'h7f8f:	data_out=16'h9ff;
17'h7f90:	data_out=16'h7e6;
17'h7f91:	data_out=16'h47e;
17'h7f92:	data_out=16'h9fd;
17'h7f93:	data_out=16'h973;
17'h7f94:	data_out=16'h9fd;
17'h7f95:	data_out=16'h88bc;
17'h7f96:	data_out=16'h83e9;
17'h7f97:	data_out=16'h9fc;
17'h7f98:	data_out=16'h81fc;
17'h7f99:	data_out=16'h4ad;
17'h7f9a:	data_out=16'h8168;
17'h7f9b:	data_out=16'h9f2;
17'h7f9c:	data_out=16'h73c;
17'h7f9d:	data_out=16'ha00;
17'h7f9e:	data_out=16'h9ff;
17'h7f9f:	data_out=16'h8811;
17'h7fa0:	data_out=16'ha00;
17'h7fa1:	data_out=16'h829e;
17'h7fa2:	data_out=16'h9fd;
17'h7fa3:	data_out=16'h8a00;
17'h7fa4:	data_out=16'h8a00;
17'h7fa5:	data_out=16'h81c0;
17'h7fa6:	data_out=16'h8a00;
17'h7fa7:	data_out=16'ha00;
17'h7fa8:	data_out=16'h8259;
17'h7fa9:	data_out=16'h9f2;
17'h7faa:	data_out=16'h9ff;
17'h7fab:	data_out=16'ha00;
17'h7fac:	data_out=16'h8679;
17'h7fad:	data_out=16'ha00;
17'h7fae:	data_out=16'ha00;
17'h7faf:	data_out=16'ha00;
17'h7fb0:	data_out=16'h8173;
17'h7fb1:	data_out=16'ha00;
17'h7fb2:	data_out=16'h81a3;
17'h7fb3:	data_out=16'ha00;
17'h7fb4:	data_out=16'ha00;
17'h7fb5:	data_out=16'h5ca;
17'h7fb6:	data_out=16'ha00;
17'h7fb7:	data_out=16'h9f8;
17'h7fb8:	data_out=16'ha00;
17'h7fb9:	data_out=16'ha00;
17'h7fba:	data_out=16'h9a0;
17'h7fbb:	data_out=16'h849a;
17'h7fbc:	data_out=16'h9f9;
17'h7fbd:	data_out=16'h69;
17'h7fbe:	data_out=16'h8255;
17'h7fbf:	data_out=16'h9d9;
17'h7fc0:	data_out=16'h861a;
17'h7fc1:	data_out=16'h9df;
17'h7fc2:	data_out=16'h99b;
17'h7fc3:	data_out=16'h89fc;
17'h7fc4:	data_out=16'h233;
17'h7fc5:	data_out=16'h88d1;
17'h7fc6:	data_out=16'h9f1;
17'h7fc7:	data_out=16'h8233;
17'h7fc8:	data_out=16'ha00;
17'h7fc9:	data_out=16'h8410;
17'h7fca:	data_out=16'ha00;
17'h7fcb:	data_out=16'h9fe;
17'h7fcc:	data_out=16'h8e3;
17'h7fcd:	data_out=16'h9ff;
17'h7fce:	data_out=16'ha00;
17'h7fcf:	data_out=16'h429;
17'h7fd0:	data_out=16'h889d;
17'h7fd1:	data_out=16'h89fa;
17'h7fd2:	data_out=16'h8a00;
17'h7fd3:	data_out=16'ha00;
17'h7fd4:	data_out=16'ha00;
17'h7fd5:	data_out=16'h8546;
17'h7fd6:	data_out=16'h8a00;
17'h7fd7:	data_out=16'h8a00;
17'h7fd8:	data_out=16'h20c;
17'h7fd9:	data_out=16'h89ef;
17'h7fda:	data_out=16'h9f7;
17'h7fdb:	data_out=16'h2af;
17'h7fdc:	data_out=16'h9fa;
17'h7fdd:	data_out=16'h9ff;
17'h7fde:	data_out=16'ha00;
17'h7fdf:	data_out=16'ha00;
17'h7fe0:	data_out=16'h89f8;
17'h7fe1:	data_out=16'h80b4;
17'h7fe2:	data_out=16'h9fd;
17'h7fe3:	data_out=16'ha00;
17'h7fe4:	data_out=16'h646;
17'h7fe5:	data_out=16'ha00;
17'h7fe6:	data_out=16'h425;
17'h7fe7:	data_out=16'ha00;
17'h7fe8:	data_out=16'h8293;
17'h7fe9:	data_out=16'h53b;
17'h7fea:	data_out=16'h82db;
17'h7feb:	data_out=16'h8098;
17'h7fec:	data_out=16'h9f9;
17'h7fed:	data_out=16'ha00;
17'h7fee:	data_out=16'h82da;
17'h7fef:	data_out=16'h9fc;
17'h7ff0:	data_out=16'h82c9;
17'h7ff1:	data_out=16'ha00;
17'h7ff2:	data_out=16'h8657;
17'h7ff3:	data_out=16'h5d;
17'h7ff4:	data_out=16'h819e;
17'h7ff5:	data_out=16'h924;
17'h7ff6:	data_out=16'h8ca;
17'h7ff7:	data_out=16'h87fa;
17'h7ff8:	data_out=16'h89fe;
17'h7ff9:	data_out=16'h9fc;
17'h7ffa:	data_out=16'ha00;
17'h7ffb:	data_out=16'h8254;
17'h7ffc:	data_out=16'h724;
17'h7ffd:	data_out=16'h831f;
17'h7ffe:	data_out=16'h89fa;
17'h7fff:	data_out=16'h89ff;
17'h8000:	data_out=16'h89ff;
17'h8001:	data_out=16'h9fb;
17'h8002:	data_out=16'h8b4;
17'h8003:	data_out=16'h895f;
17'h8004:	data_out=16'h8576;
17'h8005:	data_out=16'h9fe;
17'h8006:	data_out=16'h82bc;
17'h8007:	data_out=16'h2b8;
17'h8008:	data_out=16'h847a;
17'h8009:	data_out=16'h89ef;
17'h800a:	data_out=16'h89fb;
17'h800b:	data_out=16'h9f2;
17'h800c:	data_out=16'h8410;
17'h800d:	data_out=16'h8218;
17'h800e:	data_out=16'h851c;
17'h800f:	data_out=16'h9dd;
17'h8010:	data_out=16'h89fd;
17'h8011:	data_out=16'h449;
17'h8012:	data_out=16'h9f8;
17'h8013:	data_out=16'h845f;
17'h8014:	data_out=16'h923;
17'h8015:	data_out=16'h8a00;
17'h8016:	data_out=16'h8a00;
17'h8017:	data_out=16'h9ef;
17'h8018:	data_out=16'h8537;
17'h8019:	data_out=16'ha00;
17'h801a:	data_out=16'ha00;
17'h801b:	data_out=16'h94d;
17'h801c:	data_out=16'h67d;
17'h801d:	data_out=16'h9ff;
17'h801e:	data_out=16'h9cd;
17'h801f:	data_out=16'h875e;
17'h8020:	data_out=16'h9f9;
17'h8021:	data_out=16'h8488;
17'h8022:	data_out=16'h875;
17'h8023:	data_out=16'h8a00;
17'h8024:	data_out=16'h8a00;
17'h8025:	data_out=16'h89ff;
17'h8026:	data_out=16'h8a00;
17'h8027:	data_out=16'ha00;
17'h8028:	data_out=16'h838e;
17'h8029:	data_out=16'ha6;
17'h802a:	data_out=16'h954;
17'h802b:	data_out=16'ha00;
17'h802c:	data_out=16'h8a00;
17'h802d:	data_out=16'h818b;
17'h802e:	data_out=16'ha00;
17'h802f:	data_out=16'h9fd;
17'h8030:	data_out=16'h510;
17'h8031:	data_out=16'h9f7;
17'h8032:	data_out=16'h441;
17'h8033:	data_out=16'h9f5;
17'h8034:	data_out=16'h5ff;
17'h8035:	data_out=16'h77f;
17'h8036:	data_out=16'h78f;
17'h8037:	data_out=16'h949;
17'h8038:	data_out=16'ha00;
17'h8039:	data_out=16'h9ed;
17'h803a:	data_out=16'h319;
17'h803b:	data_out=16'h8952;
17'h803c:	data_out=16'h88b;
17'h803d:	data_out=16'h880f;
17'h803e:	data_out=16'h8387;
17'h803f:	data_out=16'h9fd;
17'h8040:	data_out=16'h854a;
17'h8041:	data_out=16'h71a;
17'h8042:	data_out=16'h8a00;
17'h8043:	data_out=16'h8851;
17'h8044:	data_out=16'h83cc;
17'h8045:	data_out=16'h8a00;
17'h8046:	data_out=16'h93b;
17'h8047:	data_out=16'h8879;
17'h8048:	data_out=16'ha00;
17'h8049:	data_out=16'h8a00;
17'h804a:	data_out=16'ha00;
17'h804b:	data_out=16'h877;
17'h804c:	data_out=16'h862c;
17'h804d:	data_out=16'h9ff;
17'h804e:	data_out=16'ha00;
17'h804f:	data_out=16'h89ff;
17'h8050:	data_out=16'h84b2;
17'h8051:	data_out=16'h8a00;
17'h8052:	data_out=16'h8a00;
17'h8053:	data_out=16'ha00;
17'h8054:	data_out=16'h9f4;
17'h8055:	data_out=16'h8a00;
17'h8056:	data_out=16'h8a00;
17'h8057:	data_out=16'h8a00;
17'h8058:	data_out=16'h89fe;
17'h8059:	data_out=16'h89e2;
17'h805a:	data_out=16'h9f9;
17'h805b:	data_out=16'h8de;
17'h805c:	data_out=16'h9fc;
17'h805d:	data_out=16'h9f0;
17'h805e:	data_out=16'h9f8;
17'h805f:	data_out=16'h9fe;
17'h8060:	data_out=16'h8a00;
17'h8061:	data_out=16'h8208;
17'h8062:	data_out=16'h9d8;
17'h8063:	data_out=16'ha00;
17'h8064:	data_out=16'h8393;
17'h8065:	data_out=16'ha00;
17'h8066:	data_out=16'ha00;
17'h8067:	data_out=16'ha00;
17'h8068:	data_out=16'h842f;
17'h8069:	data_out=16'h89fe;
17'h806a:	data_out=16'h85a5;
17'h806b:	data_out=16'h5c9;
17'h806c:	data_out=16'h230;
17'h806d:	data_out=16'h9fc;
17'h806e:	data_out=16'h85a3;
17'h806f:	data_out=16'ha00;
17'h8070:	data_out=16'h8553;
17'h8071:	data_out=16'h9f7;
17'h8072:	data_out=16'h89d9;
17'h8073:	data_out=16'h80a8;
17'h8074:	data_out=16'h4bb;
17'h8075:	data_out=16'h938;
17'h8076:	data_out=16'ha00;
17'h8077:	data_out=16'h89fa;
17'h8078:	data_out=16'hae;
17'h8079:	data_out=16'h964;
17'h807a:	data_out=16'h9f9;
17'h807b:	data_out=16'h8384;
17'h807c:	data_out=16'ha00;
17'h807d:	data_out=16'h9d1;
17'h807e:	data_out=16'h89f7;
17'h807f:	data_out=16'h85eb;
17'h8080:	data_out=16'h805b;
17'h8081:	data_out=16'h9ed;
17'h8082:	data_out=16'h420;
17'h8083:	data_out=16'h8a00;
17'h8084:	data_out=16'h8a7;
17'h8085:	data_out=16'h8144;
17'h8086:	data_out=16'h8977;
17'h8087:	data_out=16'h8148;
17'h8088:	data_out=16'h8165;
17'h8089:	data_out=16'h89e8;
17'h808a:	data_out=16'h89ff;
17'h808b:	data_out=16'h8538;
17'h808c:	data_out=16'h89f6;
17'h808d:	data_out=16'h8a00;
17'h808e:	data_out=16'h821f;
17'h808f:	data_out=16'h15c;
17'h8090:	data_out=16'h83b6;
17'h8091:	data_out=16'h9ff;
17'h8092:	data_out=16'h9e7;
17'h8093:	data_out=16'h8a00;
17'h8094:	data_out=16'h235;
17'h8095:	data_out=16'h89fd;
17'h8096:	data_out=16'h89ff;
17'h8097:	data_out=16'hd2;
17'h8098:	data_out=16'h2d9;
17'h8099:	data_out=16'ha00;
17'h809a:	data_out=16'h9ff;
17'h809b:	data_out=16'h497;
17'h809c:	data_out=16'h10d;
17'h809d:	data_out=16'h9f1;
17'h809e:	data_out=16'h80b;
17'h809f:	data_out=16'h8926;
17'h80a0:	data_out=16'h9f5;
17'h80a1:	data_out=16'h81ab;
17'h80a2:	data_out=16'h9fe;
17'h80a3:	data_out=16'h8a00;
17'h80a4:	data_out=16'h8a00;
17'h80a5:	data_out=16'h89ec;
17'h80a6:	data_out=16'h8a00;
17'h80a7:	data_out=16'h9f5;
17'h80a8:	data_out=16'h811a;
17'h80a9:	data_out=16'h83ed;
17'h80aa:	data_out=16'h9c2;
17'h80ab:	data_out=16'ha00;
17'h80ac:	data_out=16'h89ff;
17'h80ad:	data_out=16'h65a;
17'h80ae:	data_out=16'h9f3;
17'h80af:	data_out=16'h9e6;
17'h80b0:	data_out=16'hf7;
17'h80b1:	data_out=16'h24;
17'h80b2:	data_out=16'h136;
17'h80b3:	data_out=16'h9f7;
17'h80b4:	data_out=16'h8e0;
17'h80b5:	data_out=16'h6ea;
17'h80b6:	data_out=16'h9e1;
17'h80b7:	data_out=16'h420;
17'h80b8:	data_out=16'ha00;
17'h80b9:	data_out=16'h9f1;
17'h80ba:	data_out=16'h3d9;
17'h80bb:	data_out=16'h89ee;
17'h80bc:	data_out=16'h46b;
17'h80bd:	data_out=16'h645;
17'h80be:	data_out=16'h8118;
17'h80bf:	data_out=16'h8191;
17'h80c0:	data_out=16'h80bb;
17'h80c1:	data_out=16'h80a6;
17'h80c2:	data_out=16'h8a00;
17'h80c3:	data_out=16'h89ec;
17'h80c4:	data_out=16'h8705;
17'h80c5:	data_out=16'h89fd;
17'h80c6:	data_out=16'h929;
17'h80c7:	data_out=16'h842d;
17'h80c8:	data_out=16'h9ee;
17'h80c9:	data_out=16'h89f2;
17'h80ca:	data_out=16'ha00;
17'h80cb:	data_out=16'h8a00;
17'h80cc:	data_out=16'h898d;
17'h80cd:	data_out=16'ha00;
17'h80ce:	data_out=16'ha00;
17'h80cf:	data_out=16'h89ef;
17'h80d0:	data_out=16'h57;
17'h80d1:	data_out=16'h8a00;
17'h80d2:	data_out=16'h8a00;
17'h80d3:	data_out=16'ha00;
17'h80d4:	data_out=16'h9e7;
17'h80d5:	data_out=16'h8a00;
17'h80d6:	data_out=16'h89ff;
17'h80d7:	data_out=16'h89e6;
17'h80d8:	data_out=16'h89ff;
17'h80d9:	data_out=16'h80a2;
17'h80da:	data_out=16'h88e;
17'h80db:	data_out=16'ha00;
17'h80dc:	data_out=16'h9af;
17'h80dd:	data_out=16'h9c5;
17'h80de:	data_out=16'h9ce;
17'h80df:	data_out=16'h9ff;
17'h80e0:	data_out=16'h8a00;
17'h80e1:	data_out=16'h818d;
17'h80e2:	data_out=16'h138;
17'h80e3:	data_out=16'h9f8;
17'h80e4:	data_out=16'h991;
17'h80e5:	data_out=16'h6c;
17'h80e6:	data_out=16'h97c;
17'h80e7:	data_out=16'ha00;
17'h80e8:	data_out=16'h8169;
17'h80e9:	data_out=16'h89f0;
17'h80ea:	data_out=16'h8287;
17'h80eb:	data_out=16'h446;
17'h80ec:	data_out=16'h974;
17'h80ed:	data_out=16'h9f5;
17'h80ee:	data_out=16'h8284;
17'h80ef:	data_out=16'h8819;
17'h80f0:	data_out=16'h8248;
17'h80f1:	data_out=16'h9ee;
17'h80f2:	data_out=16'h84b6;
17'h80f3:	data_out=16'h18a;
17'h80f4:	data_out=16'h8030;
17'h80f5:	data_out=16'h8004;
17'h80f6:	data_out=16'ha00;
17'h80f7:	data_out=16'h89fc;
17'h80f8:	data_out=16'h820a;
17'h80f9:	data_out=16'h9fd;
17'h80fa:	data_out=16'h84e;
17'h80fb:	data_out=16'h8118;
17'h80fc:	data_out=16'ha00;
17'h80fd:	data_out=16'h8497;
17'h80fe:	data_out=16'h89e1;
17'h80ff:	data_out=16'h349;
17'h8100:	data_out=16'h8278;
17'h8101:	data_out=16'h992;
17'h8102:	data_out=16'h439;
17'h8103:	data_out=16'h89ff;
17'h8104:	data_out=16'h9c2;
17'h8105:	data_out=16'h89f6;
17'h8106:	data_out=16'h89e7;
17'h8107:	data_out=16'h85b5;
17'h8108:	data_out=16'h95f;
17'h8109:	data_out=16'h89fa;
17'h810a:	data_out=16'h85b7;
17'h810b:	data_out=16'h887e;
17'h810c:	data_out=16'h89c7;
17'h810d:	data_out=16'h89ff;
17'h810e:	data_out=16'h9c3;
17'h810f:	data_out=16'h87b4;
17'h8110:	data_out=16'h89fd;
17'h8111:	data_out=16'h9e4;
17'h8112:	data_out=16'hd6;
17'h8113:	data_out=16'h89ff;
17'h8114:	data_out=16'h89fe;
17'h8115:	data_out=16'h89ff;
17'h8116:	data_out=16'h89ff;
17'h8117:	data_out=16'h89fd;
17'h8118:	data_out=16'h8159;
17'h8119:	data_out=16'ha00;
17'h811a:	data_out=16'h2b8;
17'h811b:	data_out=16'h89fc;
17'h811c:	data_out=16'h8a00;
17'h811d:	data_out=16'h8048;
17'h811e:	data_out=16'h89fc;
17'h811f:	data_out=16'h89ea;
17'h8120:	data_out=16'h858;
17'h8121:	data_out=16'h9cd;
17'h8122:	data_out=16'h9ff;
17'h8123:	data_out=16'h89fd;
17'h8124:	data_out=16'h89fd;
17'h8125:	data_out=16'h89ec;
17'h8126:	data_out=16'h89fe;
17'h8127:	data_out=16'h82d1;
17'h8128:	data_out=16'h9de;
17'h8129:	data_out=16'h8606;
17'h812a:	data_out=16'h232;
17'h812b:	data_out=16'ha00;
17'h812c:	data_out=16'h89ff;
17'h812d:	data_out=16'h9e7;
17'h812e:	data_out=16'h660;
17'h812f:	data_out=16'h812b;
17'h8130:	data_out=16'h36d;
17'h8131:	data_out=16'h8a00;
17'h8132:	data_out=16'h341;
17'h8133:	data_out=16'h89fb;
17'h8134:	data_out=16'h1fa;
17'h8135:	data_out=16'h174;
17'h8136:	data_out=16'h595;
17'h8137:	data_out=16'h29d;
17'h8138:	data_out=16'h9a9;
17'h8139:	data_out=16'h887a;
17'h813a:	data_out=16'h89ee;
17'h813b:	data_out=16'h89fa;
17'h813c:	data_out=16'hb7;
17'h813d:	data_out=16'h8582;
17'h813e:	data_out=16'h9de;
17'h813f:	data_out=16'h89f6;
17'h8140:	data_out=16'h82b4;
17'h8141:	data_out=16'h89fc;
17'h8142:	data_out=16'h89ff;
17'h8143:	data_out=16'h89f0;
17'h8144:	data_out=16'h8959;
17'h8145:	data_out=16'h89ff;
17'h8146:	data_out=16'h9ef;
17'h8147:	data_out=16'h8634;
17'h8148:	data_out=16'h8230;
17'h8149:	data_out=16'h89f4;
17'h814a:	data_out=16'h6d1;
17'h814b:	data_out=16'h86d4;
17'h814c:	data_out=16'h87b3;
17'h814d:	data_out=16'h9ff;
17'h814e:	data_out=16'ha00;
17'h814f:	data_out=16'h89e3;
17'h8150:	data_out=16'h8771;
17'h8151:	data_out=16'h8a00;
17'h8152:	data_out=16'h8a00;
17'h8153:	data_out=16'h9bf;
17'h8154:	data_out=16'h98b;
17'h8155:	data_out=16'h8a00;
17'h8156:	data_out=16'h89fe;
17'h8157:	data_out=16'h89d7;
17'h8158:	data_out=16'h89fe;
17'h8159:	data_out=16'h8041;
17'h815a:	data_out=16'h82f4;
17'h815b:	data_out=16'h950;
17'h815c:	data_out=16'h4ca;
17'h815d:	data_out=16'h7e8;
17'h815e:	data_out=16'h8443;
17'h815f:	data_out=16'h9f5;
17'h8160:	data_out=16'h89f6;
17'h8161:	data_out=16'h8225;
17'h8162:	data_out=16'h89fe;
17'h8163:	data_out=16'h89f7;
17'h8164:	data_out=16'h5ce;
17'h8165:	data_out=16'h8733;
17'h8166:	data_out=16'h6e7;
17'h8167:	data_out=16'ha00;
17'h8168:	data_out=16'h9d8;
17'h8169:	data_out=16'h2ac;
17'h816a:	data_out=16'h9ba;
17'h816b:	data_out=16'h89f9;
17'h816c:	data_out=16'h8df;
17'h816d:	data_out=16'h89fa;
17'h816e:	data_out=16'h9ba;
17'h816f:	data_out=16'h89f7;
17'h8170:	data_out=16'h9bf;
17'h8171:	data_out=16'h93c;
17'h8172:	data_out=16'h86c2;
17'h8173:	data_out=16'h1bb;
17'h8174:	data_out=16'h20f;
17'h8175:	data_out=16'h89ec;
17'h8176:	data_out=16'ha00;
17'h8177:	data_out=16'h89fc;
17'h8178:	data_out=16'h16f;
17'h8179:	data_out=16'ha00;
17'h817a:	data_out=16'h89fc;
17'h817b:	data_out=16'h9dd;
17'h817c:	data_out=16'h9fb;
17'h817d:	data_out=16'h8952;
17'h817e:	data_out=16'h89e6;
17'h817f:	data_out=16'h8118;
17'h8180:	data_out=16'h4a0;
17'h8181:	data_out=16'h8044;
17'h8182:	data_out=16'h5d2;
17'h8183:	data_out=16'h89fa;
17'h8184:	data_out=16'h25c;
17'h8185:	data_out=16'h89f9;
17'h8186:	data_out=16'h8a00;
17'h8187:	data_out=16'h89ff;
17'h8188:	data_out=16'h84c;
17'h8189:	data_out=16'h89ee;
17'h818a:	data_out=16'h8908;
17'h818b:	data_out=16'h8882;
17'h818c:	data_out=16'h890e;
17'h818d:	data_out=16'h8a00;
17'h818e:	data_out=16'h9eb;
17'h818f:	data_out=16'h13e;
17'h8190:	data_out=16'h89f6;
17'h8191:	data_out=16'h881a;
17'h8192:	data_out=16'h8540;
17'h8193:	data_out=16'h89fe;
17'h8194:	data_out=16'h89fd;
17'h8195:	data_out=16'h89fd;
17'h8196:	data_out=16'h89fd;
17'h8197:	data_out=16'h89fc;
17'h8198:	data_out=16'h836c;
17'h8199:	data_out=16'ha00;
17'h819a:	data_out=16'h871a;
17'h819b:	data_out=16'h89fc;
17'h819c:	data_out=16'h89fe;
17'h819d:	data_out=16'h86e5;
17'h819e:	data_out=16'h89fb;
17'h819f:	data_out=16'h89ed;
17'h81a0:	data_out=16'h89da;
17'h81a1:	data_out=16'h9ea;
17'h81a2:	data_out=16'h9f7;
17'h81a3:	data_out=16'h89fc;
17'h81a4:	data_out=16'h89fc;
17'h81a5:	data_out=16'h89e1;
17'h81a6:	data_out=16'h410;
17'h81a7:	data_out=16'h89ab;
17'h81a8:	data_out=16'h9e1;
17'h81a9:	data_out=16'h84a9;
17'h81aa:	data_out=16'h823;
17'h81ab:	data_out=16'ha00;
17'h81ac:	data_out=16'h89fe;
17'h81ad:	data_out=16'h9f4;
17'h81ae:	data_out=16'h2d8;
17'h81af:	data_out=16'h89f6;
17'h81b0:	data_out=16'h77e;
17'h81b1:	data_out=16'h89ff;
17'h81b2:	data_out=16'h8004;
17'h81b3:	data_out=16'h89fa;
17'h81b4:	data_out=16'h13f;
17'h81b5:	data_out=16'h89f5;
17'h81b6:	data_out=16'h21;
17'h81b7:	data_out=16'hac;
17'h81b8:	data_out=16'h87b9;
17'h81b9:	data_out=16'h89f9;
17'h81ba:	data_out=16'h89e1;
17'h81bb:	data_out=16'h89f9;
17'h81bc:	data_out=16'h89fe;
17'h81bd:	data_out=16'h89d8;
17'h81be:	data_out=16'h9e1;
17'h81bf:	data_out=16'h89f9;
17'h81c0:	data_out=16'h88b5;
17'h81c1:	data_out=16'h89f8;
17'h81c2:	data_out=16'h89a5;
17'h81c3:	data_out=16'h89b0;
17'h81c4:	data_out=16'h89ea;
17'h81c5:	data_out=16'h89fd;
17'h81c6:	data_out=16'h9fb;
17'h81c7:	data_out=16'h15f;
17'h81c8:	data_out=16'h89fb;
17'h81c9:	data_out=16'h89e4;
17'h81ca:	data_out=16'h9c2;
17'h81cb:	data_out=16'h89fb;
17'h81cc:	data_out=16'h732;
17'h81cd:	data_out=16'h9dc;
17'h81ce:	data_out=16'ha00;
17'h81cf:	data_out=16'h8713;
17'h81d0:	data_out=16'h89f9;
17'h81d1:	data_out=16'h8a00;
17'h81d2:	data_out=16'h89fc;
17'h81d3:	data_out=16'h8919;
17'h81d4:	data_out=16'h8403;
17'h81d5:	data_out=16'h8a00;
17'h81d6:	data_out=16'h8934;
17'h81d7:	data_out=16'h89ce;
17'h81d8:	data_out=16'h8a00;
17'h81d9:	data_out=16'h89b7;
17'h81da:	data_out=16'h89fd;
17'h81db:	data_out=16'h89c2;
17'h81dc:	data_out=16'h89ff;
17'h81dd:	data_out=16'h6cc;
17'h81de:	data_out=16'h89fc;
17'h81df:	data_out=16'h9f2;
17'h81e0:	data_out=16'h87c;
17'h81e1:	data_out=16'h8661;
17'h81e2:	data_out=16'h89fc;
17'h81e3:	data_out=16'h89f9;
17'h81e4:	data_out=16'h85c1;
17'h81e5:	data_out=16'h89ed;
17'h81e6:	data_out=16'ha00;
17'h81e7:	data_out=16'ha00;
17'h81e8:	data_out=16'h9e8;
17'h81e9:	data_out=16'h4b2;
17'h81ea:	data_out=16'h9eb;
17'h81eb:	data_out=16'h89ea;
17'h81ec:	data_out=16'h984;
17'h81ed:	data_out=16'h89f9;
17'h81ee:	data_out=16'h9eb;
17'h81ef:	data_out=16'h89f5;
17'h81f0:	data_out=16'h9ea;
17'h81f1:	data_out=16'h98c;
17'h81f2:	data_out=16'h89e4;
17'h81f3:	data_out=16'h885a;
17'h81f4:	data_out=16'h627;
17'h81f5:	data_out=16'h8a00;
17'h81f6:	data_out=16'ha00;
17'h81f7:	data_out=16'h89f5;
17'h81f8:	data_out=16'h6b9;
17'h81f9:	data_out=16'h9ea;
17'h81fa:	data_out=16'h89fc;
17'h81fb:	data_out=16'h9e1;
17'h81fc:	data_out=16'h9fb;
17'h81fd:	data_out=16'h89cb;
17'h81fe:	data_out=16'h89df;
17'h81ff:	data_out=16'h8397;
17'h8200:	data_out=16'h9dc;
17'h8201:	data_out=16'h868c;
17'h8202:	data_out=16'h845;
17'h8203:	data_out=16'h8996;
17'h8204:	data_out=16'h8744;
17'h8205:	data_out=16'h89fa;
17'h8206:	data_out=16'h8a00;
17'h8207:	data_out=16'h89ff;
17'h8208:	data_out=16'h914;
17'h8209:	data_out=16'h89d2;
17'h820a:	data_out=16'h8a00;
17'h820b:	data_out=16'h87a1;
17'h820c:	data_out=16'h87b3;
17'h820d:	data_out=16'h89df;
17'h820e:	data_out=16'h9ff;
17'h820f:	data_out=16'h9e4;
17'h8210:	data_out=16'h89d0;
17'h8211:	data_out=16'h89ed;
17'h8212:	data_out=16'h89d0;
17'h8213:	data_out=16'h89b4;
17'h8214:	data_out=16'h89ed;
17'h8215:	data_out=16'h89f3;
17'h8216:	data_out=16'h89d9;
17'h8217:	data_out=16'h89e9;
17'h8218:	data_out=16'h275;
17'h8219:	data_out=16'h9fa;
17'h821a:	data_out=16'h89f1;
17'h821b:	data_out=16'h89f8;
17'h821c:	data_out=16'h89f0;
17'h821d:	data_out=16'h89c8;
17'h821e:	data_out=16'h89db;
17'h821f:	data_out=16'h89f3;
17'h8220:	data_out=16'h89e2;
17'h8221:	data_out=16'h9ff;
17'h8222:	data_out=16'ha00;
17'h8223:	data_out=16'h89ed;
17'h8224:	data_out=16'h89ed;
17'h8225:	data_out=16'h89b8;
17'h8226:	data_out=16'h9fe;
17'h8227:	data_out=16'h89e6;
17'h8228:	data_out=16'h9fe;
17'h8229:	data_out=16'h105;
17'h822a:	data_out=16'h9f6;
17'h822b:	data_out=16'ha00;
17'h822c:	data_out=16'h89e3;
17'h822d:	data_out=16'ha00;
17'h822e:	data_out=16'h81fe;
17'h822f:	data_out=16'h89ef;
17'h8230:	data_out=16'h7e1;
17'h8231:	data_out=16'h8a00;
17'h8232:	data_out=16'h889f;
17'h8233:	data_out=16'h89f6;
17'h8234:	data_out=16'h847a;
17'h8235:	data_out=16'h89ea;
17'h8236:	data_out=16'h9b5;
17'h8237:	data_out=16'h86d6;
17'h8238:	data_out=16'h89fd;
17'h8239:	data_out=16'h89f0;
17'h823a:	data_out=16'h8960;
17'h823b:	data_out=16'h89f5;
17'h823c:	data_out=16'h89ea;
17'h823d:	data_out=16'h8956;
17'h823e:	data_out=16'h9fe;
17'h823f:	data_out=16'h89fa;
17'h8240:	data_out=16'h8882;
17'h8241:	data_out=16'h89ed;
17'h8242:	data_out=16'h8417;
17'h8243:	data_out=16'h1a6;
17'h8244:	data_out=16'h89ec;
17'h8245:	data_out=16'h89f2;
17'h8246:	data_out=16'ha00;
17'h8247:	data_out=16'ha00;
17'h8248:	data_out=16'h89fc;
17'h8249:	data_out=16'h8996;
17'h824a:	data_out=16'h933;
17'h824b:	data_out=16'h8953;
17'h824c:	data_out=16'h9f9;
17'h824d:	data_out=16'ha00;
17'h824e:	data_out=16'ha00;
17'h824f:	data_out=16'h9fb;
17'h8250:	data_out=16'h89f3;
17'h8251:	data_out=16'h89f9;
17'h8252:	data_out=16'h8912;
17'h8253:	data_out=16'h89ea;
17'h8254:	data_out=16'h86b6;
17'h8255:	data_out=16'h89d8;
17'h8256:	data_out=16'h11e;
17'h8257:	data_out=16'h89a7;
17'h8258:	data_out=16'h89ff;
17'h8259:	data_out=16'h1;
17'h825a:	data_out=16'h8a00;
17'h825b:	data_out=16'h89e9;
17'h825c:	data_out=16'h8a00;
17'h825d:	data_out=16'h9d3;
17'h825e:	data_out=16'h89f5;
17'h825f:	data_out=16'h9ff;
17'h8260:	data_out=16'h9fe;
17'h8261:	data_out=16'h89f2;
17'h8262:	data_out=16'h89f0;
17'h8263:	data_out=16'h89fb;
17'h8264:	data_out=16'h85c4;
17'h8265:	data_out=16'h89f7;
17'h8266:	data_out=16'h9eb;
17'h8267:	data_out=16'ha00;
17'h8268:	data_out=16'h9ff;
17'h8269:	data_out=16'h958;
17'h826a:	data_out=16'h9ff;
17'h826b:	data_out=16'h89f0;
17'h826c:	data_out=16'ha00;
17'h826d:	data_out=16'h89fa;
17'h826e:	data_out=16'h9ff;
17'h826f:	data_out=16'h89f4;
17'h8270:	data_out=16'h9ff;
17'h8271:	data_out=16'h86c;
17'h8272:	data_out=16'h89ba;
17'h8273:	data_out=16'h89d3;
17'h8274:	data_out=16'h662;
17'h8275:	data_out=16'h8a00;
17'h8276:	data_out=16'ha00;
17'h8277:	data_out=16'h882c;
17'h8278:	data_out=16'h9a4;
17'h8279:	data_out=16'h9c7;
17'h827a:	data_out=16'h89fa;
17'h827b:	data_out=16'h9fe;
17'h827c:	data_out=16'h9e1;
17'h827d:	data_out=16'h89ee;
17'h827e:	data_out=16'h89c6;
17'h827f:	data_out=16'h89fd;
17'h8280:	data_out=16'h9fa;
17'h8281:	data_out=16'h511;
17'h8282:	data_out=16'h96a;
17'h8283:	data_out=16'h8918;
17'h8284:	data_out=16'hab;
17'h8285:	data_out=16'h8a00;
17'h8286:	data_out=16'h8a00;
17'h8287:	data_out=16'h8a00;
17'h8288:	data_out=16'h772;
17'h8289:	data_out=16'h89d2;
17'h828a:	data_out=16'h89ba;
17'h828b:	data_out=16'h88e0;
17'h828c:	data_out=16'h89d6;
17'h828d:	data_out=16'h89e1;
17'h828e:	data_out=16'ha00;
17'h828f:	data_out=16'h9e9;
17'h8290:	data_out=16'h88f7;
17'h8291:	data_out=16'h89b8;
17'h8292:	data_out=16'h89d7;
17'h8293:	data_out=16'h89a0;
17'h8294:	data_out=16'h89d9;
17'h8295:	data_out=16'h89f1;
17'h8296:	data_out=16'h89be;
17'h8297:	data_out=16'h89cb;
17'h8298:	data_out=16'h957;
17'h8299:	data_out=16'ha00;
17'h829a:	data_out=16'h89f9;
17'h829b:	data_out=16'h89eb;
17'h829c:	data_out=16'h89bc;
17'h829d:	data_out=16'h887c;
17'h829e:	data_out=16'h89b7;
17'h829f:	data_out=16'h89f3;
17'h82a0:	data_out=16'h8975;
17'h82a1:	data_out=16'ha00;
17'h82a2:	data_out=16'ha00;
17'h82a3:	data_out=16'h84ff;
17'h82a4:	data_out=16'h8508;
17'h82a5:	data_out=16'h8881;
17'h82a6:	data_out=16'ha00;
17'h82a7:	data_out=16'h89e8;
17'h82a8:	data_out=16'ha00;
17'h82a9:	data_out=16'h9fd;
17'h82aa:	data_out=16'h9ff;
17'h82ab:	data_out=16'h9f3;
17'h82ac:	data_out=16'h89cf;
17'h82ad:	data_out=16'ha00;
17'h82ae:	data_out=16'h8815;
17'h82af:	data_out=16'h89cf;
17'h82b0:	data_out=16'ha00;
17'h82b1:	data_out=16'h8a00;
17'h82b2:	data_out=16'h166;
17'h82b3:	data_out=16'h89e6;
17'h82b4:	data_out=16'h80fc;
17'h82b5:	data_out=16'h89ec;
17'h82b6:	data_out=16'h9b1;
17'h82b7:	data_out=16'h87d0;
17'h82b8:	data_out=16'h89fe;
17'h82b9:	data_out=16'h89e0;
17'h82ba:	data_out=16'h420;
17'h82bb:	data_out=16'h8a00;
17'h82bc:	data_out=16'h8961;
17'h82bd:	data_out=16'h9f4;
17'h82be:	data_out=16'ha00;
17'h82bf:	data_out=16'h8a00;
17'h82c0:	data_out=16'h51e;
17'h82c1:	data_out=16'h84e9;
17'h82c2:	data_out=16'ha00;
17'h82c3:	data_out=16'h59b;
17'h82c4:	data_out=16'h89f5;
17'h82c5:	data_out=16'h89f0;
17'h82c6:	data_out=16'ha00;
17'h82c7:	data_out=16'h9fa;
17'h82c8:	data_out=16'h89ff;
17'h82c9:	data_out=16'h863b;
17'h82ca:	data_out=16'h30a;
17'h82cb:	data_out=16'h844f;
17'h82cc:	data_out=16'ha00;
17'h82cd:	data_out=16'ha00;
17'h82ce:	data_out=16'h9df;
17'h82cf:	data_out=16'ha00;
17'h82d0:	data_out=16'h89c8;
17'h82d1:	data_out=16'h89fa;
17'h82d2:	data_out=16'hcc;
17'h82d3:	data_out=16'h89ef;
17'h82d4:	data_out=16'h745;
17'h82d5:	data_out=16'h89cb;
17'h82d6:	data_out=16'h9ad;
17'h82d7:	data_out=16'h11c;
17'h82d8:	data_out=16'h89fd;
17'h82d9:	data_out=16'h92c;
17'h82da:	data_out=16'h8a00;
17'h82db:	data_out=16'h89ae;
17'h82dc:	data_out=16'h8a00;
17'h82dd:	data_out=16'ha00;
17'h82de:	data_out=16'h89c1;
17'h82df:	data_out=16'ha00;
17'h82e0:	data_out=16'ha00;
17'h82e1:	data_out=16'h8980;
17'h82e2:	data_out=16'h89c4;
17'h82e3:	data_out=16'h89f8;
17'h82e4:	data_out=16'h83ab;
17'h82e5:	data_out=16'h89eb;
17'h82e6:	data_out=16'ha00;
17'h82e7:	data_out=16'ha00;
17'h82e8:	data_out=16'ha00;
17'h82e9:	data_out=16'h89c;
17'h82ea:	data_out=16'ha00;
17'h82eb:	data_out=16'h89f7;
17'h82ec:	data_out=16'ha00;
17'h82ed:	data_out=16'h89f3;
17'h82ee:	data_out=16'ha00;
17'h82ef:	data_out=16'h89dc;
17'h82f0:	data_out=16'ha00;
17'h82f1:	data_out=16'h698;
17'h82f2:	data_out=16'h88eb;
17'h82f3:	data_out=16'h88f5;
17'h82f4:	data_out=16'ha00;
17'h82f5:	data_out=16'h8a00;
17'h82f6:	data_out=16'ha00;
17'h82f7:	data_out=16'h9ff;
17'h82f8:	data_out=16'h9e1;
17'h82f9:	data_out=16'h9c5;
17'h82fa:	data_out=16'h89ec;
17'h82fb:	data_out=16'ha00;
17'h82fc:	data_out=16'h93d;
17'h82fd:	data_out=16'h8a00;
17'h82fe:	data_out=16'h89d7;
17'h82ff:	data_out=16'h8a00;
17'h8300:	data_out=16'h9f6;
17'h8301:	data_out=16'h6be;
17'h8302:	data_out=16'h619;
17'h8303:	data_out=16'h9e8;
17'h8304:	data_out=16'h436;
17'h8305:	data_out=16'h8a00;
17'h8306:	data_out=16'h8a00;
17'h8307:	data_out=16'h8a00;
17'h8308:	data_out=16'h442;
17'h8309:	data_out=16'h89e6;
17'h830a:	data_out=16'h8942;
17'h830b:	data_out=16'h89d8;
17'h830c:	data_out=16'h89ed;
17'h830d:	data_out=16'h8a00;
17'h830e:	data_out=16'ha00;
17'h830f:	data_out=16'h872;
17'h8310:	data_out=16'h9d3;
17'h8311:	data_out=16'h72;
17'h8312:	data_out=16'h89fb;
17'h8313:	data_out=16'h882f;
17'h8314:	data_out=16'h8a00;
17'h8315:	data_out=16'h9bc;
17'h8316:	data_out=16'h4c8;
17'h8317:	data_out=16'h8a00;
17'h8318:	data_out=16'h6ed;
17'h8319:	data_out=16'ha00;
17'h831a:	data_out=16'h8a00;
17'h831b:	data_out=16'h89f9;
17'h831c:	data_out=16'h87ee;
17'h831d:	data_out=16'h1bd;
17'h831e:	data_out=16'h89e2;
17'h831f:	data_out=16'h8a00;
17'h8320:	data_out=16'h40e;
17'h8321:	data_out=16'ha00;
17'h8322:	data_out=16'h9fd;
17'h8323:	data_out=16'h8442;
17'h8324:	data_out=16'h8407;
17'h8325:	data_out=16'h9fc;
17'h8326:	data_out=16'ha00;
17'h8327:	data_out=16'h80d9;
17'h8328:	data_out=16'h9fe;
17'h8329:	data_out=16'h9fb;
17'h832a:	data_out=16'h997;
17'h832b:	data_out=16'h8ff;
17'h832c:	data_out=16'h27c;
17'h832d:	data_out=16'h9fc;
17'h832e:	data_out=16'h8a00;
17'h832f:	data_out=16'h54f;
17'h8330:	data_out=16'ha00;
17'h8331:	data_out=16'h8a00;
17'h8332:	data_out=16'h2fc;
17'h8333:	data_out=16'h8a00;
17'h8334:	data_out=16'h7f8;
17'h8335:	data_out=16'h8378;
17'h8336:	data_out=16'h86f;
17'h8337:	data_out=16'h89ee;
17'h8338:	data_out=16'h8a00;
17'h8339:	data_out=16'h89fc;
17'h833a:	data_out=16'h235;
17'h833b:	data_out=16'h8a00;
17'h833c:	data_out=16'h895f;
17'h833d:	data_out=16'h9ee;
17'h833e:	data_out=16'h9fe;
17'h833f:	data_out=16'h8a00;
17'h8340:	data_out=16'h5d0;
17'h8341:	data_out=16'h95d;
17'h8342:	data_out=16'ha00;
17'h8343:	data_out=16'h8a;
17'h8344:	data_out=16'h8a00;
17'h8345:	data_out=16'h98c;
17'h8346:	data_out=16'ha00;
17'h8347:	data_out=16'h8b1;
17'h8348:	data_out=16'h8a00;
17'h8349:	data_out=16'ha00;
17'h834a:	data_out=16'h89fd;
17'h834b:	data_out=16'h9b3;
17'h834c:	data_out=16'ha00;
17'h834d:	data_out=16'h9fc;
17'h834e:	data_out=16'h74d;
17'h834f:	data_out=16'ha00;
17'h8350:	data_out=16'h89ea;
17'h8351:	data_out=16'h8a00;
17'h8352:	data_out=16'h5f1;
17'h8353:	data_out=16'h8a00;
17'h8354:	data_out=16'h7aa;
17'h8355:	data_out=16'h89eb;
17'h8356:	data_out=16'h9f5;
17'h8357:	data_out=16'h9d0;
17'h8358:	data_out=16'h89fe;
17'h8359:	data_out=16'h9ff;
17'h835a:	data_out=16'h8a00;
17'h835b:	data_out=16'h89fa;
17'h835c:	data_out=16'h8a00;
17'h835d:	data_out=16'ha00;
17'h835e:	data_out=16'h93a;
17'h835f:	data_out=16'h9f5;
17'h8360:	data_out=16'h9e3;
17'h8361:	data_out=16'h89de;
17'h8362:	data_out=16'h8a00;
17'h8363:	data_out=16'h8a00;
17'h8364:	data_out=16'h71b;
17'h8365:	data_out=16'h89f4;
17'h8366:	data_out=16'h9f5;
17'h8367:	data_out=16'ha00;
17'h8368:	data_out=16'ha00;
17'h8369:	data_out=16'h7b3;
17'h836a:	data_out=16'ha00;
17'h836b:	data_out=16'h89fc;
17'h836c:	data_out=16'h9fc;
17'h836d:	data_out=16'h8a00;
17'h836e:	data_out=16'ha00;
17'h836f:	data_out=16'h89f3;
17'h8370:	data_out=16'ha00;
17'h8371:	data_out=16'h89e9;
17'h8372:	data_out=16'h6e1;
17'h8373:	data_out=16'h8775;
17'h8374:	data_out=16'ha00;
17'h8375:	data_out=16'h8a00;
17'h8376:	data_out=16'ha00;
17'h8377:	data_out=16'h9ee;
17'h8378:	data_out=16'h9ba;
17'h8379:	data_out=16'h9ee;
17'h837a:	data_out=16'h8a00;
17'h837b:	data_out=16'h9fe;
17'h837c:	data_out=16'h89ae;
17'h837d:	data_out=16'h8a00;
17'h837e:	data_out=16'h8a00;
17'h837f:	data_out=16'h89e3;
17'h8380:	data_out=16'h9e9;
17'h8381:	data_out=16'h886;
17'h8382:	data_out=16'h91c;
17'h8383:	data_out=16'h9c0;
17'h8384:	data_out=16'h7d4;
17'h8385:	data_out=16'h8a00;
17'h8386:	data_out=16'h8a00;
17'h8387:	data_out=16'h89ff;
17'h8388:	data_out=16'h299;
17'h8389:	data_out=16'h89ef;
17'h838a:	data_out=16'h4f7;
17'h838b:	data_out=16'h89ea;
17'h838c:	data_out=16'h89ff;
17'h838d:	data_out=16'h3c8;
17'h838e:	data_out=16'ha00;
17'h838f:	data_out=16'h7e5;
17'h8390:	data_out=16'h94d;
17'h8391:	data_out=16'h6f9;
17'h8392:	data_out=16'h89fb;
17'h8393:	data_out=16'h597;
17'h8394:	data_out=16'h8a00;
17'h8395:	data_out=16'h9f0;
17'h8396:	data_out=16'h929;
17'h8397:	data_out=16'h8a00;
17'h8398:	data_out=16'h698;
17'h8399:	data_out=16'h8c4;
17'h839a:	data_out=16'h89ff;
17'h839b:	data_out=16'h89f6;
17'h839c:	data_out=16'h9c4;
17'h839d:	data_out=16'h498;
17'h839e:	data_out=16'h7d1;
17'h839f:	data_out=16'h8a00;
17'h83a0:	data_out=16'h548;
17'h83a1:	data_out=16'ha00;
17'h83a2:	data_out=16'h9ca;
17'h83a3:	data_out=16'h54a;
17'h83a4:	data_out=16'h554;
17'h83a5:	data_out=16'h9d9;
17'h83a6:	data_out=16'h9f2;
17'h83a7:	data_out=16'h1ac;
17'h83a8:	data_out=16'ha00;
17'h83a9:	data_out=16'h9fc;
17'h83aa:	data_out=16'h840;
17'h83ab:	data_out=16'h89fb;
17'h83ac:	data_out=16'h92e;
17'h83ad:	data_out=16'h804f;
17'h83ae:	data_out=16'h8a00;
17'h83af:	data_out=16'h816;
17'h83b0:	data_out=16'ha00;
17'h83b1:	data_out=16'h89f3;
17'h83b2:	data_out=16'h804f;
17'h83b3:	data_out=16'h8a00;
17'h83b4:	data_out=16'h86e;
17'h83b5:	data_out=16'h6a;
17'h83b6:	data_out=16'h691;
17'h83b7:	data_out=16'h85ea;
17'h83b8:	data_out=16'h8a00;
17'h83b9:	data_out=16'h8a00;
17'h83ba:	data_out=16'h89ca;
17'h83bb:	data_out=16'h8a00;
17'h83bc:	data_out=16'h988;
17'h83bd:	data_out=16'h9d8;
17'h83be:	data_out=16'ha00;
17'h83bf:	data_out=16'h8a00;
17'h83c0:	data_out=16'h741;
17'h83c1:	data_out=16'h965;
17'h83c2:	data_out=16'h9fc;
17'h83c3:	data_out=16'h837a;
17'h83c4:	data_out=16'h8a00;
17'h83c5:	data_out=16'h9ec;
17'h83c6:	data_out=16'h9c7;
17'h83c7:	data_out=16'h654;
17'h83c8:	data_out=16'h8a00;
17'h83c9:	data_out=16'ha00;
17'h83ca:	data_out=16'h89fe;
17'h83cb:	data_out=16'h965;
17'h83cc:	data_out=16'ha00;
17'h83cd:	data_out=16'h793;
17'h83ce:	data_out=16'h3f4;
17'h83cf:	data_out=16'ha00;
17'h83d0:	data_out=16'h89b4;
17'h83d1:	data_out=16'h89ff;
17'h83d2:	data_out=16'h9a7;
17'h83d3:	data_out=16'h8a00;
17'h83d4:	data_out=16'h549;
17'h83d5:	data_out=16'h89ed;
17'h83d6:	data_out=16'ha00;
17'h83d7:	data_out=16'h9f2;
17'h83d8:	data_out=16'h37a;
17'h83d9:	data_out=16'h9e9;
17'h83da:	data_out=16'h8a00;
17'h83db:	data_out=16'h185;
17'h83dc:	data_out=16'h8a00;
17'h83dd:	data_out=16'ha00;
17'h83de:	data_out=16'ha00;
17'h83df:	data_out=16'h999;
17'h83e0:	data_out=16'h89d;
17'h83e1:	data_out=16'h33c;
17'h83e2:	data_out=16'h8a00;
17'h83e3:	data_out=16'h8a00;
17'h83e4:	data_out=16'h818d;
17'h83e5:	data_out=16'h89fc;
17'h83e6:	data_out=16'h52f;
17'h83e7:	data_out=16'ha00;
17'h83e8:	data_out=16'ha00;
17'h83e9:	data_out=16'h7db;
17'h83ea:	data_out=16'ha00;
17'h83eb:	data_out=16'h898a;
17'h83ec:	data_out=16'h9db;
17'h83ed:	data_out=16'h8a00;
17'h83ee:	data_out=16'ha00;
17'h83ef:	data_out=16'h8826;
17'h83f0:	data_out=16'ha00;
17'h83f1:	data_out=16'h89fe;
17'h83f2:	data_out=16'h9c8;
17'h83f3:	data_out=16'h94b;
17'h83f4:	data_out=16'h412;
17'h83f5:	data_out=16'h8a00;
17'h83f6:	data_out=16'h8236;
17'h83f7:	data_out=16'h93e;
17'h83f8:	data_out=16'h164;
17'h83f9:	data_out=16'ha00;
17'h83fa:	data_out=16'h8a00;
17'h83fb:	data_out=16'ha00;
17'h83fc:	data_out=16'h8361;
17'h83fd:	data_out=16'h8a00;
17'h83fe:	data_out=16'h8a00;
17'h83ff:	data_out=16'h82dc;
17'h8400:	data_out=16'h9e0;
17'h8401:	data_out=16'h91a;
17'h8402:	data_out=16'hf3;
17'h8403:	data_out=16'h9c9;
17'h8404:	data_out=16'h8268;
17'h8405:	data_out=16'h89c6;
17'h8406:	data_out=16'h8a00;
17'h8407:	data_out=16'h89ff;
17'h8408:	data_out=16'h3e5;
17'h8409:	data_out=16'h89eb;
17'h840a:	data_out=16'h8469;
17'h840b:	data_out=16'h89df;
17'h840c:	data_out=16'h89ff;
17'h840d:	data_out=16'h89cb;
17'h840e:	data_out=16'h9f9;
17'h840f:	data_out=16'h81f;
17'h8410:	data_out=16'h71d;
17'h8411:	data_out=16'h9b2;
17'h8412:	data_out=16'h89fe;
17'h8413:	data_out=16'hcc;
17'h8414:	data_out=16'h89f0;
17'h8415:	data_out=16'h9bf;
17'h8416:	data_out=16'h8c1;
17'h8417:	data_out=16'h89df;
17'h8418:	data_out=16'h87f5;
17'h8419:	data_out=16'h8986;
17'h841a:	data_out=16'h89cc;
17'h841b:	data_out=16'h89d0;
17'h841c:	data_out=16'h983;
17'h841d:	data_out=16'h8f5;
17'h841e:	data_out=16'h882a;
17'h841f:	data_out=16'h8a00;
17'h8420:	data_out=16'h896c;
17'h8421:	data_out=16'h9f7;
17'h8422:	data_out=16'h325;
17'h8423:	data_out=16'h80df;
17'h8424:	data_out=16'h8079;
17'h8425:	data_out=16'h81af;
17'h8426:	data_out=16'h9b2;
17'h8427:	data_out=16'h7bd;
17'h8428:	data_out=16'h9f4;
17'h8429:	data_out=16'ha00;
17'h842a:	data_out=16'h7e6;
17'h842b:	data_out=16'h89ff;
17'h842c:	data_out=16'h8c9;
17'h842d:	data_out=16'h865f;
17'h842e:	data_out=16'h8a00;
17'h842f:	data_out=16'h91b;
17'h8430:	data_out=16'h82d9;
17'h8431:	data_out=16'h9cd;
17'h8432:	data_out=16'h89e9;
17'h8433:	data_out=16'h8a00;
17'h8434:	data_out=16'h93a;
17'h8435:	data_out=16'h8221;
17'h8436:	data_out=16'h6c8;
17'h8437:	data_out=16'h89f9;
17'h8438:	data_out=16'h8a00;
17'h8439:	data_out=16'h89f9;
17'h843a:	data_out=16'h89d7;
17'h843b:	data_out=16'h8a00;
17'h843c:	data_out=16'h9a3;
17'h843d:	data_out=16'h95a;
17'h843e:	data_out=16'h9f4;
17'h843f:	data_out=16'h89c5;
17'h8440:	data_out=16'h575;
17'h8441:	data_out=16'h9ea;
17'h8442:	data_out=16'ha00;
17'h8443:	data_out=16'h8653;
17'h8444:	data_out=16'h897d;
17'h8445:	data_out=16'h9b8;
17'h8446:	data_out=16'h99f;
17'h8447:	data_out=16'h64b;
17'h8448:	data_out=16'h89ff;
17'h8449:	data_out=16'h9a0;
17'h844a:	data_out=16'h89f2;
17'h844b:	data_out=16'h9ff;
17'h844c:	data_out=16'h9c7;
17'h844d:	data_out=16'h888b;
17'h844e:	data_out=16'h2fc;
17'h844f:	data_out=16'h9c8;
17'h8450:	data_out=16'h8987;
17'h8451:	data_out=16'h89fd;
17'h8452:	data_out=16'h9df;
17'h8453:	data_out=16'h89d0;
17'h8454:	data_out=16'h5ae;
17'h8455:	data_out=16'h89cd;
17'h8456:	data_out=16'h9fe;
17'h8457:	data_out=16'h6f;
17'h8458:	data_out=16'h51c;
17'h8459:	data_out=16'h92a;
17'h845a:	data_out=16'h8a00;
17'h845b:	data_out=16'h890c;
17'h845c:	data_out=16'h9ea;
17'h845d:	data_out=16'h9f1;
17'h845e:	data_out=16'ha00;
17'h845f:	data_out=16'h971;
17'h8460:	data_out=16'h630;
17'h8461:	data_out=16'h89ee;
17'h8462:	data_out=16'h89f2;
17'h8463:	data_out=16'h8a00;
17'h8464:	data_out=16'h892;
17'h8465:	data_out=16'h8664;
17'h8466:	data_out=16'h89c9;
17'h8467:	data_out=16'h9fd;
17'h8468:	data_out=16'h9f6;
17'h8469:	data_out=16'h8cc;
17'h846a:	data_out=16'h9fa;
17'h846b:	data_out=16'h8938;
17'h846c:	data_out=16'h9cb;
17'h846d:	data_out=16'h8a00;
17'h846e:	data_out=16'h9fa;
17'h846f:	data_out=16'h89d6;
17'h8470:	data_out=16'h9f9;
17'h8471:	data_out=16'h89ff;
17'h8472:	data_out=16'h6f4;
17'h8473:	data_out=16'h85e8;
17'h8474:	data_out=16'h8524;
17'h8475:	data_out=16'h89f0;
17'h8476:	data_out=16'h89fb;
17'h8477:	data_out=16'h897;
17'h8478:	data_out=16'h89ef;
17'h8479:	data_out=16'h9fc;
17'h847a:	data_out=16'h8a00;
17'h847b:	data_out=16'h9f4;
17'h847c:	data_out=16'h8a00;
17'h847d:	data_out=16'h8a00;
17'h847e:	data_out=16'h8a00;
17'h847f:	data_out=16'h89e0;
17'h8480:	data_out=16'h9ed;
17'h8481:	data_out=16'h9dd;
17'h8482:	data_out=16'h8a00;
17'h8483:	data_out=16'h8bf;
17'h8484:	data_out=16'h8248;
17'h8485:	data_out=16'h8991;
17'h8486:	data_out=16'h89fc;
17'h8487:	data_out=16'h8a00;
17'h8488:	data_out=16'h465;
17'h8489:	data_out=16'h89fe;
17'h848a:	data_out=16'h9b1;
17'h848b:	data_out=16'h89dd;
17'h848c:	data_out=16'h89e4;
17'h848d:	data_out=16'h89ea;
17'h848e:	data_out=16'h8050;
17'h848f:	data_out=16'h89fe;
17'h8490:	data_out=16'h8828;
17'h8491:	data_out=16'h9ff;
17'h8492:	data_out=16'h8a00;
17'h8493:	data_out=16'h16b;
17'h8494:	data_out=16'h89d6;
17'h8495:	data_out=16'h84da;
17'h8496:	data_out=16'h6b0;
17'h8497:	data_out=16'h89af;
17'h8498:	data_out=16'h8a00;
17'h8499:	data_out=16'h8a00;
17'h849a:	data_out=16'h89b7;
17'h849b:	data_out=16'h480;
17'h849c:	data_out=16'h84e;
17'h849d:	data_out=16'h9fb;
17'h849e:	data_out=16'h89ee;
17'h849f:	data_out=16'h8a00;
17'h84a0:	data_out=16'h897a;
17'h84a1:	data_out=16'h819e;
17'h84a2:	data_out=16'h89ff;
17'h84a3:	data_out=16'h89e0;
17'h84a4:	data_out=16'h89e0;
17'h84a5:	data_out=16'h8a00;
17'h84a6:	data_out=16'h661;
17'h84a7:	data_out=16'h8e8;
17'h84a8:	data_out=16'h82d4;
17'h84a9:	data_out=16'h9ec;
17'h84aa:	data_out=16'h8211;
17'h84ab:	data_out=16'h8a00;
17'h84ac:	data_out=16'hf3;
17'h84ad:	data_out=16'h8899;
17'h84ae:	data_out=16'h89ff;
17'h84af:	data_out=16'h974;
17'h84b0:	data_out=16'h87be;
17'h84b1:	data_out=16'h9fe;
17'h84b2:	data_out=16'h8a00;
17'h84b3:	data_out=16'h89fa;
17'h84b4:	data_out=16'h9e3;
17'h84b5:	data_out=16'h83f4;
17'h84b6:	data_out=16'h553;
17'h84b7:	data_out=16'h8a00;
17'h84b8:	data_out=16'h9d7;
17'h84b9:	data_out=16'h89fa;
17'h84ba:	data_out=16'h8a00;
17'h84bb:	data_out=16'h8a00;
17'h84bc:	data_out=16'h9cd;
17'h84bd:	data_out=16'h663;
17'h84be:	data_out=16'h82d0;
17'h84bf:	data_out=16'h8992;
17'h84c0:	data_out=16'h89fc;
17'h84c1:	data_out=16'h9f7;
17'h84c2:	data_out=16'ha00;
17'h84c3:	data_out=16'h89d3;
17'h84c4:	data_out=16'h82db;
17'h84c5:	data_out=16'h8368;
17'h84c6:	data_out=16'h9bd;
17'h84c7:	data_out=16'h8a00;
17'h84c8:	data_out=16'h88f6;
17'h84c9:	data_out=16'h8a00;
17'h84ca:	data_out=16'h89cf;
17'h84cb:	data_out=16'ha00;
17'h84cc:	data_out=16'h92c;
17'h84cd:	data_out=16'h89ff;
17'h84ce:	data_out=16'h891a;
17'h84cf:	data_out=16'h91f;
17'h84d0:	data_out=16'h899b;
17'h84d1:	data_out=16'h89fe;
17'h84d2:	data_out=16'h8202;
17'h84d3:	data_out=16'h87bf;
17'h84d4:	data_out=16'h4ba;
17'h84d5:	data_out=16'h89e5;
17'h84d6:	data_out=16'h9ed;
17'h84d7:	data_out=16'h8a00;
17'h84d8:	data_out=16'h633;
17'h84d9:	data_out=16'h8772;
17'h84da:	data_out=16'h996;
17'h84db:	data_out=16'h89b9;
17'h84dc:	data_out=16'ha00;
17'h84dd:	data_out=16'h9d3;
17'h84de:	data_out=16'ha00;
17'h84df:	data_out=16'h881f;
17'h84e0:	data_out=16'h8a00;
17'h84e1:	data_out=16'h895d;
17'h84e2:	data_out=16'h89b5;
17'h84e3:	data_out=16'h89f2;
17'h84e4:	data_out=16'h93a;
17'h84e5:	data_out=16'h9d6;
17'h84e6:	data_out=16'h8a00;
17'h84e7:	data_out=16'h214;
17'h84e8:	data_out=16'h825d;
17'h84e9:	data_out=16'h70c;
17'h84ea:	data_out=16'h5d;
17'h84eb:	data_out=16'h8947;
17'h84ec:	data_out=16'h9db;
17'h84ed:	data_out=16'h89f4;
17'h84ee:	data_out=16'h5b;
17'h84ef:	data_out=16'h89da;
17'h84f0:	data_out=16'h7;
17'h84f1:	data_out=16'h8a00;
17'h84f2:	data_out=16'h2b6;
17'h84f3:	data_out=16'h8725;
17'h84f4:	data_out=16'h88af;
17'h84f5:	data_out=16'h384;
17'h84f6:	data_out=16'h8a00;
17'h84f7:	data_out=16'hbb;
17'h84f8:	data_out=16'h89f7;
17'h84f9:	data_out=16'h7b8;
17'h84fa:	data_out=16'h89e6;
17'h84fb:	data_out=16'h82ce;
17'h84fc:	data_out=16'h8a00;
17'h84fd:	data_out=16'h8a00;
17'h84fe:	data_out=16'h8a00;
17'h84ff:	data_out=16'h89f1;
17'h8500:	data_out=16'ha00;
17'h8501:	data_out=16'h9ea;
17'h8502:	data_out=16'h8a00;
17'h8503:	data_out=16'h97f;
17'h8504:	data_out=16'h8a00;
17'h8505:	data_out=16'h8355;
17'h8506:	data_out=16'h67e;
17'h8507:	data_out=16'h8a00;
17'h8508:	data_out=16'h9da;
17'h8509:	data_out=16'h8a00;
17'h850a:	data_out=16'h8092;
17'h850b:	data_out=16'h99b;
17'h850c:	data_out=16'h81ba;
17'h850d:	data_out=16'h8538;
17'h850e:	data_out=16'h8a00;
17'h850f:	data_out=16'h8a00;
17'h8510:	data_out=16'h3c1;
17'h8511:	data_out=16'h9fe;
17'h8512:	data_out=16'h8a00;
17'h8513:	data_out=16'h4e1;
17'h8514:	data_out=16'h487;
17'h8515:	data_out=16'h86fa;
17'h8516:	data_out=16'h918;
17'h8517:	data_out=16'h99c;
17'h8518:	data_out=16'h8a00;
17'h8519:	data_out=16'h8a00;
17'h851a:	data_out=16'h89f2;
17'h851b:	data_out=16'h9c5;
17'h851c:	data_out=16'h9f9;
17'h851d:	data_out=16'ha00;
17'h851e:	data_out=16'h84aa;
17'h851f:	data_out=16'h8a00;
17'h8520:	data_out=16'h954;
17'h8521:	data_out=16'h8a00;
17'h8522:	data_out=16'h8a00;
17'h8523:	data_out=16'h8a00;
17'h8524:	data_out=16'h8a00;
17'h8525:	data_out=16'h8a00;
17'h8526:	data_out=16'h8a00;
17'h8527:	data_out=16'h9c4;
17'h8528:	data_out=16'h8a00;
17'h8529:	data_out=16'h8805;
17'h852a:	data_out=16'h8a00;
17'h852b:	data_out=16'h89c8;
17'h852c:	data_out=16'h910;
17'h852d:	data_out=16'h8244;
17'h852e:	data_out=16'h89fe;
17'h852f:	data_out=16'h9e2;
17'h8530:	data_out=16'h8960;
17'h8531:	data_out=16'h9fe;
17'h8532:	data_out=16'h8a00;
17'h8533:	data_out=16'h852b;
17'h8534:	data_out=16'h9ff;
17'h8535:	data_out=16'h8a00;
17'h8536:	data_out=16'h62a;
17'h8537:	data_out=16'h8a00;
17'h8538:	data_out=16'ha00;
17'h8539:	data_out=16'h804b;
17'h853a:	data_out=16'h8a00;
17'h853b:	data_out=16'h8a00;
17'h853c:	data_out=16'h9dc;
17'h853d:	data_out=16'h81af;
17'h853e:	data_out=16'h8a00;
17'h853f:	data_out=16'h83b1;
17'h8540:	data_out=16'h8a00;
17'h8541:	data_out=16'ha00;
17'h8542:	data_out=16'h9e8;
17'h8543:	data_out=16'h89fd;
17'h8544:	data_out=16'h9ca;
17'h8545:	data_out=16'h8523;
17'h8546:	data_out=16'h9e4;
17'h8547:	data_out=16'h8a00;
17'h8548:	data_out=16'h8350;
17'h8549:	data_out=16'h8a00;
17'h854a:	data_out=16'h88aa;
17'h854b:	data_out=16'ha00;
17'h854c:	data_out=16'h8a00;
17'h854d:	data_out=16'h8a00;
17'h854e:	data_out=16'h8a00;
17'h854f:	data_out=16'h8a00;
17'h8550:	data_out=16'h887;
17'h8551:	data_out=16'h89fd;
17'h8552:	data_out=16'h8a00;
17'h8553:	data_out=16'h9ff;
17'h8554:	data_out=16'h9cf;
17'h8555:	data_out=16'h89fe;
17'h8556:	data_out=16'h8a00;
17'h8557:	data_out=16'h8a00;
17'h8558:	data_out=16'h3d2;
17'h8559:	data_out=16'h8a00;
17'h855a:	data_out=16'ha00;
17'h855b:	data_out=16'h89db;
17'h855c:	data_out=16'ha00;
17'h855d:	data_out=16'h8e0;
17'h855e:	data_out=16'ha00;
17'h855f:	data_out=16'h89b7;
17'h8560:	data_out=16'h8a00;
17'h8561:	data_out=16'h8a00;
17'h8562:	data_out=16'h989;
17'h8563:	data_out=16'h1a5;
17'h8564:	data_out=16'ha00;
17'h8565:	data_out=16'h958;
17'h8566:	data_out=16'h8a00;
17'h8567:	data_out=16'h8a00;
17'h8568:	data_out=16'h8a00;
17'h8569:	data_out=16'h6c5;
17'h856a:	data_out=16'h8a00;
17'h856b:	data_out=16'h8853;
17'h856c:	data_out=16'h9e1;
17'h856d:	data_out=16'h147;
17'h856e:	data_out=16'h8a00;
17'h856f:	data_out=16'h8a00;
17'h8570:	data_out=16'h8a00;
17'h8571:	data_out=16'h8a00;
17'h8572:	data_out=16'h8a00;
17'h8573:	data_out=16'h89e5;
17'h8574:	data_out=16'h8982;
17'h8575:	data_out=16'ha00;
17'h8576:	data_out=16'h8a00;
17'h8577:	data_out=16'h8a00;
17'h8578:	data_out=16'h89ed;
17'h8579:	data_out=16'h85a1;
17'h857a:	data_out=16'h536;
17'h857b:	data_out=16'h8a00;
17'h857c:	data_out=16'h8a00;
17'h857d:	data_out=16'h8a00;
17'h857e:	data_out=16'h8a00;
17'h857f:	data_out=16'h89f5;
17'h8580:	data_out=16'ha00;
17'h8581:	data_out=16'h9ef;
17'h8582:	data_out=16'h8a00;
17'h8583:	data_out=16'h9dd;
17'h8584:	data_out=16'h8a00;
17'h8585:	data_out=16'h8602;
17'h8586:	data_out=16'h9c9;
17'h8587:	data_out=16'h8a00;
17'h8588:	data_out=16'h998;
17'h8589:	data_out=16'h8a00;
17'h858a:	data_out=16'h8a00;
17'h858b:	data_out=16'h9ff;
17'h858c:	data_out=16'h84aa;
17'h858d:	data_out=16'h7d7;
17'h858e:	data_out=16'h8a00;
17'h858f:	data_out=16'h8a00;
17'h8590:	data_out=16'h80f9;
17'h8591:	data_out=16'h9fc;
17'h8592:	data_out=16'h770;
17'h8593:	data_out=16'h876;
17'h8594:	data_out=16'h9fc;
17'h8595:	data_out=16'h643;
17'h8596:	data_out=16'h9bd;
17'h8597:	data_out=16'h9fe;
17'h8598:	data_out=16'h8a00;
17'h8599:	data_out=16'h8a00;
17'h859a:	data_out=16'h8a00;
17'h859b:	data_out=16'h9e5;
17'h859c:	data_out=16'h9f7;
17'h859d:	data_out=16'ha00;
17'h859e:	data_out=16'h91e;
17'h859f:	data_out=16'h89bd;
17'h85a0:	data_out=16'h9fd;
17'h85a1:	data_out=16'h8a00;
17'h85a2:	data_out=16'h8a00;
17'h85a3:	data_out=16'h8a00;
17'h85a4:	data_out=16'h8a00;
17'h85a5:	data_out=16'h8a00;
17'h85a6:	data_out=16'h8a00;
17'h85a7:	data_out=16'h9ec;
17'h85a8:	data_out=16'h8a00;
17'h85a9:	data_out=16'h89ee;
17'h85aa:	data_out=16'h8a00;
17'h85ab:	data_out=16'h9fa;
17'h85ac:	data_out=16'h9ce;
17'h85ad:	data_out=16'hbe;
17'h85ae:	data_out=16'h8986;
17'h85af:	data_out=16'h9fb;
17'h85b0:	data_out=16'h8a00;
17'h85b1:	data_out=16'h9f5;
17'h85b2:	data_out=16'h8a00;
17'h85b3:	data_out=16'ha00;
17'h85b4:	data_out=16'ha00;
17'h85b5:	data_out=16'h8a00;
17'h85b6:	data_out=16'h723;
17'h85b7:	data_out=16'h8a00;
17'h85b8:	data_out=16'ha00;
17'h85b9:	data_out=16'ha00;
17'h85ba:	data_out=16'h8a00;
17'h85bb:	data_out=16'h8a00;
17'h85bc:	data_out=16'h880;
17'h85bd:	data_out=16'h8273;
17'h85be:	data_out=16'h8a00;
17'h85bf:	data_out=16'h8674;
17'h85c0:	data_out=16'h8a00;
17'h85c1:	data_out=16'ha00;
17'h85c2:	data_out=16'h8e1;
17'h85c3:	data_out=16'h8a00;
17'h85c4:	data_out=16'h9ba;
17'h85c5:	data_out=16'h7b7;
17'h85c6:	data_out=16'h89e1;
17'h85c7:	data_out=16'h8a00;
17'h85c8:	data_out=16'h820;
17'h85c9:	data_out=16'h8a00;
17'h85ca:	data_out=16'h9ef;
17'h85cb:	data_out=16'h9f9;
17'h85cc:	data_out=16'h8a00;
17'h85cd:	data_out=16'h8a00;
17'h85ce:	data_out=16'h8852;
17'h85cf:	data_out=16'h8a00;
17'h85d0:	data_out=16'h98e;
17'h85d1:	data_out=16'h89fa;
17'h85d2:	data_out=16'h8a00;
17'h85d3:	data_out=16'ha00;
17'h85d4:	data_out=16'h9fd;
17'h85d5:	data_out=16'h89fc;
17'h85d6:	data_out=16'h8a00;
17'h85d7:	data_out=16'h8a00;
17'h85d8:	data_out=16'h9df;
17'h85d9:	data_out=16'h8a00;
17'h85da:	data_out=16'ha00;
17'h85db:	data_out=16'h89e7;
17'h85dc:	data_out=16'ha00;
17'h85dd:	data_out=16'h9d0;
17'h85de:	data_out=16'ha00;
17'h85df:	data_out=16'h83ea;
17'h85e0:	data_out=16'h8a00;
17'h85e1:	data_out=16'h8a00;
17'h85e2:	data_out=16'ha00;
17'h85e3:	data_out=16'ha00;
17'h85e4:	data_out=16'ha00;
17'h85e5:	data_out=16'h922;
17'h85e6:	data_out=16'h89e0;
17'h85e7:	data_out=16'h8a00;
17'h85e8:	data_out=16'h8a00;
17'h85e9:	data_out=16'h885f;
17'h85ea:	data_out=16'h8a00;
17'h85eb:	data_out=16'h8ec;
17'h85ec:	data_out=16'h9f2;
17'h85ed:	data_out=16'ha00;
17'h85ee:	data_out=16'h8a00;
17'h85ef:	data_out=16'h8a00;
17'h85f0:	data_out=16'h8a00;
17'h85f1:	data_out=16'h89ff;
17'h85f2:	data_out=16'h8a00;
17'h85f3:	data_out=16'h8a00;
17'h85f4:	data_out=16'h8a00;
17'h85f5:	data_out=16'h994;
17'h85f6:	data_out=16'h8a00;
17'h85f7:	data_out=16'h8a00;
17'h85f8:	data_out=16'h8a00;
17'h85f9:	data_out=16'h8932;
17'h85fa:	data_out=16'ha00;
17'h85fb:	data_out=16'h8a00;
17'h85fc:	data_out=16'h89fe;
17'h85fd:	data_out=16'h89fa;
17'h85fe:	data_out=16'h72e;
17'h85ff:	data_out=16'h89fd;
17'h8600:	data_out=16'h9ff;
17'h8601:	data_out=16'h9ee;
17'h8602:	data_out=16'h8a00;
17'h8603:	data_out=16'h892;
17'h8604:	data_out=16'h8a00;
17'h8605:	data_out=16'h8a00;
17'h8606:	data_out=16'h9ff;
17'h8607:	data_out=16'h8a00;
17'h8608:	data_out=16'h81f4;
17'h8609:	data_out=16'h89b2;
17'h860a:	data_out=16'h89c3;
17'h860b:	data_out=16'ha00;
17'h860c:	data_out=16'h89c3;
17'h860d:	data_out=16'h814c;
17'h860e:	data_out=16'h8a00;
17'h860f:	data_out=16'h89fc;
17'h8610:	data_out=16'h8a00;
17'h8611:	data_out=16'ha00;
17'h8612:	data_out=16'h9d0;
17'h8613:	data_out=16'h3a7;
17'h8614:	data_out=16'h9fb;
17'h8615:	data_out=16'h8a00;
17'h8616:	data_out=16'h7b9;
17'h8617:	data_out=16'h9fc;
17'h8618:	data_out=16'h89fe;
17'h8619:	data_out=16'h8a00;
17'h861a:	data_out=16'h8a00;
17'h861b:	data_out=16'h522;
17'h861c:	data_out=16'h996;
17'h861d:	data_out=16'ha00;
17'h861e:	data_out=16'h944;
17'h861f:	data_out=16'h87d4;
17'h8620:	data_out=16'h9ee;
17'h8621:	data_out=16'h8a00;
17'h8622:	data_out=16'h8a00;
17'h8623:	data_out=16'h8a00;
17'h8624:	data_out=16'h8a00;
17'h8625:	data_out=16'h8a00;
17'h8626:	data_out=16'h8a00;
17'h8627:	data_out=16'h9ff;
17'h8628:	data_out=16'h8a00;
17'h8629:	data_out=16'h8a00;
17'h862a:	data_out=16'h8a00;
17'h862b:	data_out=16'ha00;
17'h862c:	data_out=16'h7da;
17'h862d:	data_out=16'ha00;
17'h862e:	data_out=16'h86d9;
17'h862f:	data_out=16'h9f8;
17'h8630:	data_out=16'h8a00;
17'h8631:	data_out=16'h9c0;
17'h8632:	data_out=16'h8a00;
17'h8633:	data_out=16'ha00;
17'h8634:	data_out=16'ha00;
17'h8635:	data_out=16'h89ff;
17'h8636:	data_out=16'h62a;
17'h8637:	data_out=16'h8a00;
17'h8638:	data_out=16'ha00;
17'h8639:	data_out=16'ha00;
17'h863a:	data_out=16'h8a00;
17'h863b:	data_out=16'h8a00;
17'h863c:	data_out=16'h8a00;
17'h863d:	data_out=16'h89fb;
17'h863e:	data_out=16'h8a00;
17'h863f:	data_out=16'h8a00;
17'h8640:	data_out=16'h8a00;
17'h8641:	data_out=16'h9fe;
17'h8642:	data_out=16'h451;
17'h8643:	data_out=16'h8a00;
17'h8644:	data_out=16'h946;
17'h8645:	data_out=16'h8a00;
17'h8646:	data_out=16'h89fe;
17'h8647:	data_out=16'h8988;
17'h8648:	data_out=16'h9f7;
17'h8649:	data_out=16'h8a00;
17'h864a:	data_out=16'h9f7;
17'h864b:	data_out=16'h9e3;
17'h864c:	data_out=16'h8a00;
17'h864d:	data_out=16'h8a00;
17'h864e:	data_out=16'h238;
17'h864f:	data_out=16'h8a00;
17'h8650:	data_out=16'h89fc;
17'h8651:	data_out=16'h8a00;
17'h8652:	data_out=16'h8a00;
17'h8653:	data_out=16'ha00;
17'h8654:	data_out=16'h9f1;
17'h8655:	data_out=16'h89f9;
17'h8656:	data_out=16'h8a00;
17'h8657:	data_out=16'h8a00;
17'h8658:	data_out=16'h89f9;
17'h8659:	data_out=16'h8a00;
17'h865a:	data_out=16'ha00;
17'h865b:	data_out=16'h89b1;
17'h865c:	data_out=16'h990;
17'h865d:	data_out=16'h53a;
17'h865e:	data_out=16'ha00;
17'h865f:	data_out=16'h205;
17'h8660:	data_out=16'h8a00;
17'h8661:	data_out=16'h8a00;
17'h8662:	data_out=16'h9d7;
17'h8663:	data_out=16'ha00;
17'h8664:	data_out=16'ha00;
17'h8665:	data_out=16'h21d;
17'h8666:	data_out=16'h89be;
17'h8667:	data_out=16'h8a00;
17'h8668:	data_out=16'h8a00;
17'h8669:	data_out=16'h89de;
17'h866a:	data_out=16'h8a00;
17'h866b:	data_out=16'h89fd;
17'h866c:	data_out=16'h9f3;
17'h866d:	data_out=16'ha00;
17'h866e:	data_out=16'h8a00;
17'h866f:	data_out=16'h8a00;
17'h8670:	data_out=16'h8a00;
17'h8671:	data_out=16'h8119;
17'h8672:	data_out=16'h8a00;
17'h8673:	data_out=16'h8a00;
17'h8674:	data_out=16'h8a00;
17'h8675:	data_out=16'h8a00;
17'h8676:	data_out=16'h89a4;
17'h8677:	data_out=16'h8a00;
17'h8678:	data_out=16'h8a00;
17'h8679:	data_out=16'h89c8;
17'h867a:	data_out=16'ha00;
17'h867b:	data_out=16'h8a00;
17'h867c:	data_out=16'h89f6;
17'h867d:	data_out=16'h8980;
17'h867e:	data_out=16'ha00;
17'h867f:	data_out=16'h8a00;
17'h8680:	data_out=16'h9aa;
17'h8681:	data_out=16'h9fa;
17'h8682:	data_out=16'h8a00;
17'h8683:	data_out=16'h730;
17'h8684:	data_out=16'h89ff;
17'h8685:	data_out=16'h8a00;
17'h8686:	data_out=16'ha00;
17'h8687:	data_out=16'h89f7;
17'h8688:	data_out=16'h81b8;
17'h8689:	data_out=16'h8995;
17'h868a:	data_out=16'h9ce;
17'h868b:	data_out=16'ha00;
17'h868c:	data_out=16'h89cb;
17'h868d:	data_out=16'h8a00;
17'h868e:	data_out=16'h89f9;
17'h868f:	data_out=16'h89c7;
17'h8690:	data_out=16'h89da;
17'h8691:	data_out=16'ha00;
17'h8692:	data_out=16'h986;
17'h8693:	data_out=16'h82bb;
17'h8694:	data_out=16'h9fa;
17'h8695:	data_out=16'h89ff;
17'h8696:	data_out=16'h8931;
17'h8697:	data_out=16'h9f9;
17'h8698:	data_out=16'h89ff;
17'h8699:	data_out=16'h8a00;
17'h869a:	data_out=16'h89ff;
17'h869b:	data_out=16'h76f;
17'h869c:	data_out=16'h855c;
17'h869d:	data_out=16'ha00;
17'h869e:	data_out=16'h9e4;
17'h869f:	data_out=16'h29a;
17'h86a0:	data_out=16'h9f1;
17'h86a1:	data_out=16'h89fa;
17'h86a2:	data_out=16'h89e9;
17'h86a3:	data_out=16'h8a00;
17'h86a4:	data_out=16'h8a00;
17'h86a5:	data_out=16'h8a00;
17'h86a6:	data_out=16'h8078;
17'h86a7:	data_out=16'ha00;
17'h86a8:	data_out=16'h89f7;
17'h86a9:	data_out=16'h89fe;
17'h86aa:	data_out=16'h8015;
17'h86ab:	data_out=16'ha00;
17'h86ac:	data_out=16'h89fc;
17'h86ad:	data_out=16'ha00;
17'h86ae:	data_out=16'h9f1;
17'h86af:	data_out=16'h9f3;
17'h86b0:	data_out=16'h8a00;
17'h86b1:	data_out=16'h9ed;
17'h86b2:	data_out=16'h8a00;
17'h86b3:	data_out=16'ha00;
17'h86b4:	data_out=16'ha00;
17'h86b5:	data_out=16'h829c;
17'h86b6:	data_out=16'h693;
17'h86b7:	data_out=16'h89f5;
17'h86b8:	data_out=16'ha00;
17'h86b9:	data_out=16'ha00;
17'h86ba:	data_out=16'h89d2;
17'h86bb:	data_out=16'h89fa;
17'h86bc:	data_out=16'h88ea;
17'h86bd:	data_out=16'h89bf;
17'h86be:	data_out=16'h89f7;
17'h86bf:	data_out=16'h8a00;
17'h86c0:	data_out=16'h8a00;
17'h86c1:	data_out=16'h9af;
17'h86c2:	data_out=16'h352;
17'h86c3:	data_out=16'h8a00;
17'h86c4:	data_out=16'h9e4;
17'h86c5:	data_out=16'h89ff;
17'h86c6:	data_out=16'h1c6;
17'h86c7:	data_out=16'h829;
17'h86c8:	data_out=16'h9e6;
17'h86c9:	data_out=16'h8a00;
17'h86ca:	data_out=16'h9d4;
17'h86cb:	data_out=16'h96f;
17'h86cc:	data_out=16'h8a00;
17'h86cd:	data_out=16'h89e9;
17'h86ce:	data_out=16'h6c2;
17'h86cf:	data_out=16'h8a00;
17'h86d0:	data_out=16'h89ef;
17'h86d1:	data_out=16'h8a00;
17'h86d2:	data_out=16'h8a00;
17'h86d3:	data_out=16'h9f1;
17'h86d4:	data_out=16'h9e1;
17'h86d5:	data_out=16'h82e6;
17'h86d6:	data_out=16'h8a00;
17'h86d7:	data_out=16'h8a00;
17'h86d8:	data_out=16'h89f9;
17'h86d9:	data_out=16'h8a00;
17'h86da:	data_out=16'h9fd;
17'h86db:	data_out=16'h9d7;
17'h86dc:	data_out=16'h99f;
17'h86dd:	data_out=16'h85a9;
17'h86de:	data_out=16'ha00;
17'h86df:	data_out=16'h9f1;
17'h86e0:	data_out=16'h9a1;
17'h86e1:	data_out=16'h8a00;
17'h86e2:	data_out=16'h9e9;
17'h86e3:	data_out=16'ha00;
17'h86e4:	data_out=16'ha00;
17'h86e5:	data_out=16'h9cc;
17'h86e6:	data_out=16'h89ed;
17'h86e7:	data_out=16'h8a00;
17'h86e8:	data_out=16'h89fb;
17'h86e9:	data_out=16'h8772;
17'h86ea:	data_out=16'h89f6;
17'h86eb:	data_out=16'h89ee;
17'h86ec:	data_out=16'h985;
17'h86ed:	data_out=16'ha00;
17'h86ee:	data_out=16'h89f6;
17'h86ef:	data_out=16'h8a00;
17'h86f0:	data_out=16'h89f9;
17'h86f1:	data_out=16'h8e4;
17'h86f2:	data_out=16'h8a00;
17'h86f3:	data_out=16'h8a00;
17'h86f4:	data_out=16'h8a00;
17'h86f5:	data_out=16'h8a00;
17'h86f6:	data_out=16'h9f2;
17'h86f7:	data_out=16'h8a00;
17'h86f8:	data_out=16'h8a00;
17'h86f9:	data_out=16'hfd;
17'h86fa:	data_out=16'h9fd;
17'h86fb:	data_out=16'h89f7;
17'h86fc:	data_out=16'h89f8;
17'h86fd:	data_out=16'h8511;
17'h86fe:	data_out=16'ha00;
17'h86ff:	data_out=16'h8a00;
17'h8700:	data_out=16'h82f9;
17'h8701:	data_out=16'ha00;
17'h8702:	data_out=16'h89ed;
17'h8703:	data_out=16'h8733;
17'h8704:	data_out=16'h89d8;
17'h8705:	data_out=16'h89fc;
17'h8706:	data_out=16'h9ff;
17'h8707:	data_out=16'h8a00;
17'h8708:	data_out=16'h894a;
17'h8709:	data_out=16'h8783;
17'h870a:	data_out=16'ha00;
17'h870b:	data_out=16'h9fe;
17'h870c:	data_out=16'h89fd;
17'h870d:	data_out=16'h8a00;
17'h870e:	data_out=16'h65d;
17'h870f:	data_out=16'h89e9;
17'h8710:	data_out=16'h88db;
17'h8711:	data_out=16'ha00;
17'h8712:	data_out=16'h59f;
17'h8713:	data_out=16'h61f;
17'h8714:	data_out=16'h9e9;
17'h8715:	data_out=16'h89fc;
17'h8716:	data_out=16'h89fa;
17'h8717:	data_out=16'h9e2;
17'h8718:	data_out=16'h8a00;
17'h8719:	data_out=16'h89fe;
17'h871a:	data_out=16'h89fe;
17'h871b:	data_out=16'h8048;
17'h871c:	data_out=16'h870b;
17'h871d:	data_out=16'ha00;
17'h871e:	data_out=16'h9e5;
17'h871f:	data_out=16'h9f7;
17'h8720:	data_out=16'h956;
17'h8721:	data_out=16'h5e7;
17'h8722:	data_out=16'h88dc;
17'h8723:	data_out=16'h89d6;
17'h8724:	data_out=16'h89d7;
17'h8725:	data_out=16'h89e0;
17'h8726:	data_out=16'h9df;
17'h8727:	data_out=16'ha00;
17'h8728:	data_out=16'h693;
17'h8729:	data_out=16'h89d4;
17'h872a:	data_out=16'h778;
17'h872b:	data_out=16'h9fc;
17'h872c:	data_out=16'h89f9;
17'h872d:	data_out=16'ha00;
17'h872e:	data_out=16'h9f0;
17'h872f:	data_out=16'h5d6;
17'h8730:	data_out=16'h8a00;
17'h8731:	data_out=16'ha00;
17'h8732:	data_out=16'h89fc;
17'h8733:	data_out=16'h9f9;
17'h8734:	data_out=16'ha00;
17'h8735:	data_out=16'h9fb;
17'h8736:	data_out=16'h83b0;
17'h8737:	data_out=16'h585;
17'h8738:	data_out=16'ha00;
17'h8739:	data_out=16'h9fa;
17'h873a:	data_out=16'h80fb;
17'h873b:	data_out=16'h8247;
17'h873c:	data_out=16'h9f1;
17'h873d:	data_out=16'h8180;
17'h873e:	data_out=16'h6a0;
17'h873f:	data_out=16'h89fb;
17'h8740:	data_out=16'h89ed;
17'h8741:	data_out=16'h8a00;
17'h8742:	data_out=16'h89df;
17'h8743:	data_out=16'h8a00;
17'h8744:	data_out=16'h9eb;
17'h8745:	data_out=16'h89fc;
17'h8746:	data_out=16'h9f9;
17'h8747:	data_out=16'h97f;
17'h8748:	data_out=16'h9b2;
17'h8749:	data_out=16'h89b8;
17'h874a:	data_out=16'h8593;
17'h874b:	data_out=16'h2;
17'h874c:	data_out=16'h89fd;
17'h874d:	data_out=16'h8809;
17'h874e:	data_out=16'h5a6;
17'h874f:	data_out=16'h89a8;
17'h8750:	data_out=16'h89f9;
17'h8751:	data_out=16'h8a00;
17'h8752:	data_out=16'h89ee;
17'h8753:	data_out=16'h9d5;
17'h8754:	data_out=16'h9ef;
17'h8755:	data_out=16'h190;
17'h8756:	data_out=16'h89a0;
17'h8757:	data_out=16'h8962;
17'h8758:	data_out=16'h89fd;
17'h8759:	data_out=16'h89c4;
17'h875a:	data_out=16'h9d0;
17'h875b:	data_out=16'ha00;
17'h875c:	data_out=16'h971;
17'h875d:	data_out=16'h8447;
17'h875e:	data_out=16'ha00;
17'h875f:	data_out=16'h84f1;
17'h8760:	data_out=16'h9ef;
17'h8761:	data_out=16'h16;
17'h8762:	data_out=16'h9eb;
17'h8763:	data_out=16'h9f8;
17'h8764:	data_out=16'ha00;
17'h8765:	data_out=16'h9f6;
17'h8766:	data_out=16'h8a00;
17'h8767:	data_out=16'h89e9;
17'h8768:	data_out=16'h619;
17'h8769:	data_out=16'h89e7;
17'h876a:	data_out=16'h69f;
17'h876b:	data_out=16'h8989;
17'h876c:	data_out=16'h8738;
17'h876d:	data_out=16'h9f9;
17'h876e:	data_out=16'h69a;
17'h876f:	data_out=16'h89ff;
17'h8770:	data_out=16'h670;
17'h8771:	data_out=16'h855;
17'h8772:	data_out=16'h88f5;
17'h8773:	data_out=16'h8918;
17'h8774:	data_out=16'h8a00;
17'h8775:	data_out=16'h89fc;
17'h8776:	data_out=16'h9f2;
17'h8777:	data_out=16'h8a00;
17'h8778:	data_out=16'h8a00;
17'h8779:	data_out=16'h8788;
17'h877a:	data_out=16'h9f4;
17'h877b:	data_out=16'h6a0;
17'h877c:	data_out=16'h8a00;
17'h877d:	data_out=16'h819c;
17'h877e:	data_out=16'ha00;
17'h877f:	data_out=16'h8a00;
17'h8780:	data_out=16'h89ea;
17'h8781:	data_out=16'ha00;
17'h8782:	data_out=16'h86a2;
17'h8783:	data_out=16'h89fa;
17'h8784:	data_out=16'h898a;
17'h8785:	data_out=16'h89f6;
17'h8786:	data_out=16'ha00;
17'h8787:	data_out=16'h8a00;
17'h8788:	data_out=16'h89b5;
17'h8789:	data_out=16'h8795;
17'h878a:	data_out=16'ha00;
17'h878b:	data_out=16'h9f3;
17'h878c:	data_out=16'h89ee;
17'h878d:	data_out=16'h8a00;
17'h878e:	data_out=16'h9f7;
17'h878f:	data_out=16'h89c4;
17'h8790:	data_out=16'h89d1;
17'h8791:	data_out=16'ha00;
17'h8792:	data_out=16'h232;
17'h8793:	data_out=16'h713;
17'h8794:	data_out=16'h937;
17'h8795:	data_out=16'h8a00;
17'h8796:	data_out=16'h8a00;
17'h8797:	data_out=16'h9de;
17'h8798:	data_out=16'h8a00;
17'h8799:	data_out=16'h89af;
17'h879a:	data_out=16'h89f5;
17'h879b:	data_out=16'h88b3;
17'h879c:	data_out=16'h89fb;
17'h879d:	data_out=16'ha00;
17'h879e:	data_out=16'h572;
17'h879f:	data_out=16'h9e5;
17'h87a0:	data_out=16'h832c;
17'h87a1:	data_out=16'h9f6;
17'h87a2:	data_out=16'h867a;
17'h87a3:	data_out=16'ha00;
17'h87a4:	data_out=16'ha00;
17'h87a5:	data_out=16'h8933;
17'h87a6:	data_out=16'h8609;
17'h87a7:	data_out=16'h9fd;
17'h87a8:	data_out=16'h9f5;
17'h87a9:	data_out=16'h89e2;
17'h87aa:	data_out=16'h890d;
17'h87ab:	data_out=16'h9f0;
17'h87ac:	data_out=16'h8a00;
17'h87ad:	data_out=16'ha00;
17'h87ae:	data_out=16'h9fe;
17'h87af:	data_out=16'h8217;
17'h87b0:	data_out=16'h89ff;
17'h87b1:	data_out=16'ha00;
17'h87b2:	data_out=16'h8802;
17'h87b3:	data_out=16'h9e4;
17'h87b4:	data_out=16'ha00;
17'h87b5:	data_out=16'hba;
17'h87b6:	data_out=16'h86d8;
17'h87b7:	data_out=16'h9c7;
17'h87b8:	data_out=16'ha00;
17'h87b9:	data_out=16'h7db;
17'h87ba:	data_out=16'h89bc;
17'h87bb:	data_out=16'h8294;
17'h87bc:	data_out=16'h9f9;
17'h87bd:	data_out=16'h86b8;
17'h87be:	data_out=16'h9f5;
17'h87bf:	data_out=16'h89f6;
17'h87c0:	data_out=16'h8899;
17'h87c1:	data_out=16'h8a00;
17'h87c2:	data_out=16'h89db;
17'h87c3:	data_out=16'h8a00;
17'h87c4:	data_out=16'h693;
17'h87c5:	data_out=16'h8a00;
17'h87c6:	data_out=16'h9ff;
17'h87c7:	data_out=16'h8384;
17'h87c8:	data_out=16'h9f8;
17'h87c9:	data_out=16'h88e7;
17'h87ca:	data_out=16'h8809;
17'h87cb:	data_out=16'h89d5;
17'h87cc:	data_out=16'h89f5;
17'h87cd:	data_out=16'h83e8;
17'h87ce:	data_out=16'h753;
17'h87cf:	data_out=16'h871e;
17'h87d0:	data_out=16'h8a00;
17'h87d1:	data_out=16'h8a00;
17'h87d2:	data_out=16'h8609;
17'h87d3:	data_out=16'h9f7;
17'h87d4:	data_out=16'h80b9;
17'h87d5:	data_out=16'h83cb;
17'h87d6:	data_out=16'h88d6;
17'h87d7:	data_out=16'h4;
17'h87d8:	data_out=16'h8a00;
17'h87d9:	data_out=16'h888c;
17'h87da:	data_out=16'h87a;
17'h87db:	data_out=16'ha00;
17'h87dc:	data_out=16'h9af;
17'h87dd:	data_out=16'h879c;
17'h87de:	data_out=16'hc7;
17'h87df:	data_out=16'h8760;
17'h87e0:	data_out=16'h9f1;
17'h87e1:	data_out=16'h9a1;
17'h87e2:	data_out=16'h9ef;
17'h87e3:	data_out=16'h9eb;
17'h87e4:	data_out=16'h9fe;
17'h87e5:	data_out=16'h9f9;
17'h87e6:	data_out=16'h89df;
17'h87e7:	data_out=16'h89f8;
17'h87e8:	data_out=16'h9f6;
17'h87e9:	data_out=16'h8a00;
17'h87ea:	data_out=16'h9f7;
17'h87eb:	data_out=16'h895c;
17'h87ec:	data_out=16'h89f0;
17'h87ed:	data_out=16'h9eb;
17'h87ee:	data_out=16'h9f7;
17'h87ef:	data_out=16'h89fc;
17'h87f0:	data_out=16'h9f7;
17'h87f1:	data_out=16'h5f8;
17'h87f2:	data_out=16'h86f0;
17'h87f3:	data_out=16'h85b0;
17'h87f4:	data_out=16'h89e6;
17'h87f5:	data_out=16'h89f7;
17'h87f6:	data_out=16'h9f1;
17'h87f7:	data_out=16'h8a00;
17'h87f8:	data_out=16'h8a00;
17'h87f9:	data_out=16'h8a00;
17'h87fa:	data_out=16'h9ea;
17'h87fb:	data_out=16'h9f5;
17'h87fc:	data_out=16'h8a00;
17'h87fd:	data_out=16'h80b6;
17'h87fe:	data_out=16'ha00;
17'h87ff:	data_out=16'h8a00;
17'h8800:	data_out=16'h89bd;
17'h8801:	data_out=16'ha00;
17'h8802:	data_out=16'h443;
17'h8803:	data_out=16'h89ea;
17'h8804:	data_out=16'h8968;
17'h8805:	data_out=16'h89bb;
17'h8806:	data_out=16'ha00;
17'h8807:	data_out=16'h8a00;
17'h8808:	data_out=16'h887f;
17'h8809:	data_out=16'h89f1;
17'h880a:	data_out=16'ha00;
17'h880b:	data_out=16'h681;
17'h880c:	data_out=16'h89c3;
17'h880d:	data_out=16'h8a00;
17'h880e:	data_out=16'h9f5;
17'h880f:	data_out=16'h899f;
17'h8810:	data_out=16'h89e1;
17'h8811:	data_out=16'ha00;
17'h8812:	data_out=16'h823d;
17'h8813:	data_out=16'h892;
17'h8814:	data_out=16'h82a5;
17'h8815:	data_out=16'h8a00;
17'h8816:	data_out=16'h8a00;
17'h8817:	data_out=16'h1bf;
17'h8818:	data_out=16'h8a00;
17'h8819:	data_out=16'h89aa;
17'h881a:	data_out=16'h89b8;
17'h881b:	data_out=16'h82;
17'h881c:	data_out=16'h89c0;
17'h881d:	data_out=16'ha00;
17'h881e:	data_out=16'h8934;
17'h881f:	data_out=16'h9d7;
17'h8820:	data_out=16'h87af;
17'h8821:	data_out=16'h9f5;
17'h8822:	data_out=16'h896e;
17'h8823:	data_out=16'ha00;
17'h8824:	data_out=16'ha00;
17'h8825:	data_out=16'h89fc;
17'h8826:	data_out=16'h88e4;
17'h8827:	data_out=16'h56f;
17'h8828:	data_out=16'h9f5;
17'h8829:	data_out=16'h8a00;
17'h882a:	data_out=16'h8828;
17'h882b:	data_out=16'h9f2;
17'h882c:	data_out=16'h8a00;
17'h882d:	data_out=16'ha00;
17'h882e:	data_out=16'ha00;
17'h882f:	data_out=16'h8628;
17'h8830:	data_out=16'h89cf;
17'h8831:	data_out=16'ha00;
17'h8832:	data_out=16'h8603;
17'h8833:	data_out=16'h81af;
17'h8834:	data_out=16'ha00;
17'h8835:	data_out=16'h8561;
17'h8836:	data_out=16'h8699;
17'h8837:	data_out=16'h9f0;
17'h8838:	data_out=16'ha00;
17'h8839:	data_out=16'h89c2;
17'h883a:	data_out=16'h8a00;
17'h883b:	data_out=16'h84aa;
17'h883c:	data_out=16'h9ff;
17'h883d:	data_out=16'h893d;
17'h883e:	data_out=16'h9f5;
17'h883f:	data_out=16'h89be;
17'h8840:	data_out=16'h886e;
17'h8841:	data_out=16'h89b3;
17'h8842:	data_out=16'h89ab;
17'h8843:	data_out=16'h8a00;
17'h8844:	data_out=16'h8404;
17'h8845:	data_out=16'h8a00;
17'h8846:	data_out=16'h9fe;
17'h8847:	data_out=16'h89e6;
17'h8848:	data_out=16'h9ff;
17'h8849:	data_out=16'h89ef;
17'h884a:	data_out=16'h837b;
17'h884b:	data_out=16'h8977;
17'h884c:	data_out=16'h89fc;
17'h884d:	data_out=16'h87e8;
17'h884e:	data_out=16'h9e8;
17'h884f:	data_out=16'h896b;
17'h8850:	data_out=16'h8a00;
17'h8851:	data_out=16'h89ff;
17'h8852:	data_out=16'h86f1;
17'h8853:	data_out=16'h9fd;
17'h8854:	data_out=16'h8591;
17'h8855:	data_out=16'h85b5;
17'h8856:	data_out=16'h889b;
17'h8857:	data_out=16'h89a3;
17'h8858:	data_out=16'h89fb;
17'h8859:	data_out=16'h8980;
17'h885a:	data_out=16'h9e4;
17'h885b:	data_out=16'ha00;
17'h885c:	data_out=16'h9fe;
17'h885d:	data_out=16'h892d;
17'h885e:	data_out=16'h8516;
17'h885f:	data_out=16'h8931;
17'h8860:	data_out=16'h4b8;
17'h8861:	data_out=16'h8055;
17'h8862:	data_out=16'hf9;
17'h8863:	data_out=16'h9b1;
17'h8864:	data_out=16'ha00;
17'h8865:	data_out=16'h9fb;
17'h8866:	data_out=16'h89c0;
17'h8867:	data_out=16'h89fc;
17'h8868:	data_out=16'h9f5;
17'h8869:	data_out=16'h89da;
17'h886a:	data_out=16'h9f5;
17'h886b:	data_out=16'h8988;
17'h886c:	data_out=16'h89d5;
17'h886d:	data_out=16'h8b9;
17'h886e:	data_out=16'h9f5;
17'h886f:	data_out=16'h89c2;
17'h8870:	data_out=16'h9f5;
17'h8871:	data_out=16'h8333;
17'h8872:	data_out=16'h88fa;
17'h8873:	data_out=16'h87bc;
17'h8874:	data_out=16'h8963;
17'h8875:	data_out=16'h858;
17'h8876:	data_out=16'h9f6;
17'h8877:	data_out=16'h89ff;
17'h8878:	data_out=16'h8a00;
17'h8879:	data_out=16'h8a00;
17'h887a:	data_out=16'h66c;
17'h887b:	data_out=16'h9f5;
17'h887c:	data_out=16'h8a00;
17'h887d:	data_out=16'h89ff;
17'h887e:	data_out=16'ha00;
17'h887f:	data_out=16'h8a00;
17'h8880:	data_out=16'h8998;
17'h8881:	data_out=16'ha00;
17'h8882:	data_out=16'h6bc;
17'h8883:	data_out=16'h89fe;
17'h8884:	data_out=16'h8988;
17'h8885:	data_out=16'h89db;
17'h8886:	data_out=16'ha00;
17'h8887:	data_out=16'h89da;
17'h8888:	data_out=16'h876d;
17'h8889:	data_out=16'h89fe;
17'h888a:	data_out=16'h76b;
17'h888b:	data_out=16'h88f7;
17'h888c:	data_out=16'h8997;
17'h888d:	data_out=16'h8a00;
17'h888e:	data_out=16'h9f5;
17'h888f:	data_out=16'h8975;
17'h8890:	data_out=16'h8a00;
17'h8891:	data_out=16'ha00;
17'h8892:	data_out=16'h301;
17'h8893:	data_out=16'h5fb;
17'h8894:	data_out=16'h89d0;
17'h8895:	data_out=16'h8a00;
17'h8896:	data_out=16'h8a00;
17'h8897:	data_out=16'h89a3;
17'h8898:	data_out=16'h89ff;
17'h8899:	data_out=16'h89e5;
17'h889a:	data_out=16'h89d0;
17'h889b:	data_out=16'h89a9;
17'h889c:	data_out=16'h89ef;
17'h889d:	data_out=16'ha00;
17'h889e:	data_out=16'h89d1;
17'h889f:	data_out=16'h8968;
17'h88a0:	data_out=16'h896c;
17'h88a1:	data_out=16'h9f5;
17'h88a2:	data_out=16'h89ff;
17'h88a3:	data_out=16'ha00;
17'h88a4:	data_out=16'ha00;
17'h88a5:	data_out=16'h8a00;
17'h88a6:	data_out=16'h830b;
17'h88a7:	data_out=16'h831e;
17'h88a8:	data_out=16'h9f5;
17'h88a9:	data_out=16'h8a00;
17'h88aa:	data_out=16'h87a5;
17'h88ab:	data_out=16'h8916;
17'h88ac:	data_out=16'h8a00;
17'h88ad:	data_out=16'ha00;
17'h88ae:	data_out=16'ha00;
17'h88af:	data_out=16'h8900;
17'h88b0:	data_out=16'h89de;
17'h88b1:	data_out=16'h8016;
17'h88b2:	data_out=16'h8666;
17'h88b3:	data_out=16'h89db;
17'h88b4:	data_out=16'ha00;
17'h88b5:	data_out=16'h88d0;
17'h88b6:	data_out=16'h8718;
17'h88b7:	data_out=16'h9c6;
17'h88b8:	data_out=16'ha00;
17'h88b9:	data_out=16'h89ed;
17'h88ba:	data_out=16'h8a00;
17'h88bb:	data_out=16'h887e;
17'h88bc:	data_out=16'h9ed;
17'h88bd:	data_out=16'h89b0;
17'h88be:	data_out=16'h9f5;
17'h88bf:	data_out=16'h89dd;
17'h88c0:	data_out=16'h89a6;
17'h88c1:	data_out=16'h89b6;
17'h88c2:	data_out=16'h88c7;
17'h88c3:	data_out=16'h8a00;
17'h88c4:	data_out=16'h87c4;
17'h88c5:	data_out=16'h8a00;
17'h88c6:	data_out=16'h9fd;
17'h88c7:	data_out=16'h89e9;
17'h88c8:	data_out=16'ha00;
17'h88c9:	data_out=16'h8a00;
17'h88ca:	data_out=16'h810f;
17'h88cb:	data_out=16'h87d1;
17'h88cc:	data_out=16'h89ff;
17'h88cd:	data_out=16'h89f2;
17'h88ce:	data_out=16'h9df;
17'h88cf:	data_out=16'h89ee;
17'h88d0:	data_out=16'h8a00;
17'h88d1:	data_out=16'h89ff;
17'h88d2:	data_out=16'h2eb;
17'h88d3:	data_out=16'ha00;
17'h88d4:	data_out=16'h8826;
17'h88d5:	data_out=16'h89fc;
17'h88d6:	data_out=16'h8931;
17'h88d7:	data_out=16'h89fb;
17'h88d8:	data_out=16'h89fe;
17'h88d9:	data_out=16'h89c7;
17'h88da:	data_out=16'h9f3;
17'h88db:	data_out=16'ha00;
17'h88dc:	data_out=16'h9fd;
17'h88dd:	data_out=16'h8997;
17'h88de:	data_out=16'h8873;
17'h88df:	data_out=16'h897e;
17'h88e0:	data_out=16'h704;
17'h88e1:	data_out=16'hf5;
17'h88e2:	data_out=16'h8978;
17'h88e3:	data_out=16'h899e;
17'h88e4:	data_out=16'ha00;
17'h88e5:	data_out=16'h8996;
17'h88e6:	data_out=16'h89e4;
17'h88e7:	data_out=16'h89f8;
17'h88e8:	data_out=16'h9f4;
17'h88e9:	data_out=16'h89ba;
17'h88ea:	data_out=16'h9f4;
17'h88eb:	data_out=16'h89cd;
17'h88ec:	data_out=16'h89b4;
17'h88ed:	data_out=16'h89ab;
17'h88ee:	data_out=16'h9f4;
17'h88ef:	data_out=16'h89e2;
17'h88f0:	data_out=16'h9f4;
17'h88f1:	data_out=16'h14f;
17'h88f2:	data_out=16'h89d6;
17'h88f3:	data_out=16'h88d1;
17'h88f4:	data_out=16'h88b4;
17'h88f5:	data_out=16'h83d;
17'h88f6:	data_out=16'h87c9;
17'h88f7:	data_out=16'h8a00;
17'h88f8:	data_out=16'h8a00;
17'h88f9:	data_out=16'h8a00;
17'h88fa:	data_out=16'h8997;
17'h88fb:	data_out=16'h9f5;
17'h88fc:	data_out=16'h89fb;
17'h88fd:	data_out=16'h89f7;
17'h88fe:	data_out=16'ha00;
17'h88ff:	data_out=16'h8a00;
17'h8900:	data_out=16'h87c1;
17'h8901:	data_out=16'ha00;
17'h8902:	data_out=16'h89e;
17'h8903:	data_out=16'h8a00;
17'h8904:	data_out=16'h8941;
17'h8905:	data_out=16'h89fe;
17'h8906:	data_out=16'ha00;
17'h8907:	data_out=16'h89e1;
17'h8908:	data_out=16'h6f3;
17'h8909:	data_out=16'h8a00;
17'h890a:	data_out=16'h9ff;
17'h890b:	data_out=16'h89a8;
17'h890c:	data_out=16'h89ce;
17'h890d:	data_out=16'h8a00;
17'h890e:	data_out=16'h9f9;
17'h890f:	data_out=16'h894b;
17'h8910:	data_out=16'h8a00;
17'h8911:	data_out=16'ha00;
17'h8912:	data_out=16'h5da;
17'h8913:	data_out=16'h879c;
17'h8914:	data_out=16'h89fd;
17'h8915:	data_out=16'h89fe;
17'h8916:	data_out=16'h8a00;
17'h8917:	data_out=16'h89fa;
17'h8918:	data_out=16'h89fd;
17'h8919:	data_out=16'h8a00;
17'h891a:	data_out=16'h89fc;
17'h891b:	data_out=16'h89b4;
17'h891c:	data_out=16'h89ff;
17'h891d:	data_out=16'ha00;
17'h891e:	data_out=16'h89f9;
17'h891f:	data_out=16'h89f2;
17'h8920:	data_out=16'h89e2;
17'h8921:	data_out=16'h9f9;
17'h8922:	data_out=16'h8a00;
17'h8923:	data_out=16'ha00;
17'h8924:	data_out=16'ha00;
17'h8925:	data_out=16'h8a00;
17'h8926:	data_out=16'h9ff;
17'h8927:	data_out=16'h8795;
17'h8928:	data_out=16'h9f8;
17'h8929:	data_out=16'h8a00;
17'h892a:	data_out=16'h8700;
17'h892b:	data_out=16'h89c7;
17'h892c:	data_out=16'h8a00;
17'h892d:	data_out=16'ha00;
17'h892e:	data_out=16'h8305;
17'h892f:	data_out=16'h89c6;
17'h8930:	data_out=16'h88a8;
17'h8931:	data_out=16'h8368;
17'h8932:	data_out=16'h89c3;
17'h8933:	data_out=16'h89fa;
17'h8934:	data_out=16'ha00;
17'h8935:	data_out=16'h391;
17'h8936:	data_out=16'h87ae;
17'h8937:	data_out=16'h8c3;
17'h8938:	data_out=16'ha00;
17'h8939:	data_out=16'h89fa;
17'h893a:	data_out=16'h8a00;
17'h893b:	data_out=16'h7c7;
17'h893c:	data_out=16'h8991;
17'h893d:	data_out=16'h89f2;
17'h893e:	data_out=16'h9f8;
17'h893f:	data_out=16'h89fe;
17'h8940:	data_out=16'h89f3;
17'h8941:	data_out=16'h89aa;
17'h8942:	data_out=16'h80f;
17'h8943:	data_out=16'h8a00;
17'h8944:	data_out=16'h8919;
17'h8945:	data_out=16'h89fe;
17'h8946:	data_out=16'ha00;
17'h8947:	data_out=16'h89ff;
17'h8948:	data_out=16'h851a;
17'h8949:	data_out=16'h89fd;
17'h894a:	data_out=16'h88c6;
17'h894b:	data_out=16'h86df;
17'h894c:	data_out=16'h8a00;
17'h894d:	data_out=16'h89ff;
17'h894e:	data_out=16'h4e5;
17'h894f:	data_out=16'h89fe;
17'h8950:	data_out=16'h8a00;
17'h8951:	data_out=16'h8a00;
17'h8952:	data_out=16'h9f8;
17'h8953:	data_out=16'h8856;
17'h8954:	data_out=16'h8995;
17'h8955:	data_out=16'h89fd;
17'h8956:	data_out=16'ha00;
17'h8957:	data_out=16'h8716;
17'h8958:	data_out=16'h89dd;
17'h8959:	data_out=16'h89f9;
17'h895a:	data_out=16'h789;
17'h895b:	data_out=16'ha00;
17'h895c:	data_out=16'h897e;
17'h895d:	data_out=16'h89e5;
17'h895e:	data_out=16'h89ba;
17'h895f:	data_out=16'h89c7;
17'h8960:	data_out=16'h9fc;
17'h8961:	data_out=16'h3c5;
17'h8962:	data_out=16'h89cb;
17'h8963:	data_out=16'h89f7;
17'h8964:	data_out=16'ha00;
17'h8965:	data_out=16'h89f5;
17'h8966:	data_out=16'h8a00;
17'h8967:	data_out=16'h89ff;
17'h8968:	data_out=16'h9f8;
17'h8969:	data_out=16'hbb;
17'h896a:	data_out=16'h9f9;
17'h896b:	data_out=16'h89ff;
17'h896c:	data_out=16'h85a8;
17'h896d:	data_out=16'h89f9;
17'h896e:	data_out=16'h9f9;
17'h896f:	data_out=16'h89ff;
17'h8970:	data_out=16'h9f9;
17'h8971:	data_out=16'h2e3;
17'h8972:	data_out=16'h89fe;
17'h8973:	data_out=16'h89ec;
17'h8974:	data_out=16'h8498;
17'h8975:	data_out=16'h876d;
17'h8976:	data_out=16'h89f0;
17'h8977:	data_out=16'h8a00;
17'h8978:	data_out=16'h8a00;
17'h8979:	data_out=16'h89af;
17'h897a:	data_out=16'h89ee;
17'h897b:	data_out=16'h9f8;
17'h897c:	data_out=16'h8873;
17'h897d:	data_out=16'h89fc;
17'h897e:	data_out=16'h675;
17'h897f:	data_out=16'h8a00;
17'h8980:	data_out=16'ha00;
17'h8981:	data_out=16'ha00;
17'h8982:	data_out=16'ha00;
17'h8983:	data_out=16'h8a00;
17'h8984:	data_out=16'ha00;
17'h8985:	data_out=16'h89fb;
17'h8986:	data_out=16'h9f0;
17'h8987:	data_out=16'h89fd;
17'h8988:	data_out=16'ha00;
17'h8989:	data_out=16'h8a00;
17'h898a:	data_out=16'ha00;
17'h898b:	data_out=16'h89f6;
17'h898c:	data_out=16'h8a00;
17'h898d:	data_out=16'h8a00;
17'h898e:	data_out=16'ha00;
17'h898f:	data_out=16'h3f7;
17'h8990:	data_out=16'h8a00;
17'h8991:	data_out=16'h6b6;
17'h8992:	data_out=16'h3f9;
17'h8993:	data_out=16'h89f5;
17'h8994:	data_out=16'h8a00;
17'h8995:	data_out=16'h86a;
17'h8996:	data_out=16'h89ff;
17'h8997:	data_out=16'h8a00;
17'h8998:	data_out=16'h9fe;
17'h8999:	data_out=16'h8a00;
17'h899a:	data_out=16'h89f9;
17'h899b:	data_out=16'h8a00;
17'h899c:	data_out=16'h8a00;
17'h899d:	data_out=16'ha00;
17'h899e:	data_out=16'h89fe;
17'h899f:	data_out=16'h89fe;
17'h89a0:	data_out=16'h89e3;
17'h89a1:	data_out=16'ha00;
17'h89a2:	data_out=16'h8a00;
17'h89a3:	data_out=16'ha00;
17'h89a4:	data_out=16'ha00;
17'h89a5:	data_out=16'h885a;
17'h89a6:	data_out=16'ha00;
17'h89a7:	data_out=16'h341;
17'h89a8:	data_out=16'h9fd;
17'h89a9:	data_out=16'h8a00;
17'h89aa:	data_out=16'ha00;
17'h89ab:	data_out=16'h8a00;
17'h89ac:	data_out=16'h89ff;
17'h89ad:	data_out=16'ha00;
17'h89ae:	data_out=16'h89cf;
17'h89af:	data_out=16'h89fb;
17'h89b0:	data_out=16'ha00;
17'h89b1:	data_out=16'h2ac;
17'h89b2:	data_out=16'ha00;
17'h89b3:	data_out=16'h8a00;
17'h89b4:	data_out=16'ha00;
17'h89b5:	data_out=16'ha00;
17'h89b6:	data_out=16'h6dc;
17'h89b7:	data_out=16'h9ff;
17'h89b8:	data_out=16'ha00;
17'h89b9:	data_out=16'h8a00;
17'h89ba:	data_out=16'h89ff;
17'h89bb:	data_out=16'ha00;
17'h89bc:	data_out=16'h89dc;
17'h89bd:	data_out=16'h8911;
17'h89be:	data_out=16'h9fd;
17'h89bf:	data_out=16'h89fa;
17'h89c0:	data_out=16'h8941;
17'h89c1:	data_out=16'h886f;
17'h89c2:	data_out=16'ha00;
17'h89c3:	data_out=16'h8a00;
17'h89c4:	data_out=16'h7;
17'h89c5:	data_out=16'h7a0;
17'h89c6:	data_out=16'ha00;
17'h89c7:	data_out=16'h89fe;
17'h89c8:	data_out=16'h893b;
17'h89c9:	data_out=16'h816a;
17'h89ca:	data_out=16'h89e5;
17'h89cb:	data_out=16'h87f1;
17'h89cc:	data_out=16'h72e;
17'h89cd:	data_out=16'h8a00;
17'h89ce:	data_out=16'h579;
17'h89cf:	data_out=16'h9f9;
17'h89d0:	data_out=16'h8a00;
17'h89d1:	data_out=16'h89fe;
17'h89d2:	data_out=16'ha00;
17'h89d3:	data_out=16'h89d0;
17'h89d4:	data_out=16'h8996;
17'h89d5:	data_out=16'h89ff;
17'h89d6:	data_out=16'ha00;
17'h89d7:	data_out=16'h9f7;
17'h89d8:	data_out=16'h45f;
17'h89d9:	data_out=16'h9f3;
17'h89da:	data_out=16'h8a00;
17'h89db:	data_out=16'ha00;
17'h89dc:	data_out=16'h89fe;
17'h89dd:	data_out=16'he2;
17'h89de:	data_out=16'h89f7;
17'h89df:	data_out=16'h820;
17'h89e0:	data_out=16'ha00;
17'h89e1:	data_out=16'ha00;
17'h89e2:	data_out=16'h8a00;
17'h89e3:	data_out=16'h8a00;
17'h89e4:	data_out=16'h8f2;
17'h89e5:	data_out=16'h8a00;
17'h89e6:	data_out=16'h8a00;
17'h89e7:	data_out=16'h8a00;
17'h89e8:	data_out=16'h9ff;
17'h89e9:	data_out=16'ha00;
17'h89ea:	data_out=16'ha00;
17'h89eb:	data_out=16'h89fe;
17'h89ec:	data_out=16'ha00;
17'h89ed:	data_out=16'h8a00;
17'h89ee:	data_out=16'ha00;
17'h89ef:	data_out=16'h8a00;
17'h89f0:	data_out=16'ha00;
17'h89f1:	data_out=16'h10a;
17'h89f2:	data_out=16'h10f;
17'h89f3:	data_out=16'h630;
17'h89f4:	data_out=16'ha00;
17'h89f5:	data_out=16'hac;
17'h89f6:	data_out=16'h8a00;
17'h89f7:	data_out=16'h8a00;
17'h89f8:	data_out=16'h8a00;
17'h89f9:	data_out=16'h8578;
17'h89fa:	data_out=16'h8a00;
17'h89fb:	data_out=16'h9fd;
17'h89fc:	data_out=16'ha00;
17'h89fd:	data_out=16'h8a00;
17'h89fe:	data_out=16'h876f;
17'h89ff:	data_out=16'h8a00;
17'h8a00:	data_out=16'ha00;
17'h8a01:	data_out=16'ha00;
17'h8a02:	data_out=16'ha00;
17'h8a03:	data_out=16'h89fe;
17'h8a04:	data_out=16'ha00;
17'h8a05:	data_out=16'ha00;
17'h8a06:	data_out=16'h8a00;
17'h8a07:	data_out=16'h8a00;
17'h8a08:	data_out=16'ha00;
17'h8a09:	data_out=16'h8a00;
17'h8a0a:	data_out=16'ha00;
17'h8a0b:	data_out=16'h8a00;
17'h8a0c:	data_out=16'h86d7;
17'h8a0d:	data_out=16'ha00;
17'h8a0e:	data_out=16'ha00;
17'h8a0f:	data_out=16'ha00;
17'h8a10:	data_out=16'h8a00;
17'h8a11:	data_out=16'h973;
17'h8a12:	data_out=16'h85b6;
17'h8a13:	data_out=16'h87bf;
17'h8a14:	data_out=16'h89ff;
17'h8a15:	data_out=16'ha00;
17'h8a16:	data_out=16'ha00;
17'h8a17:	data_out=16'h8a00;
17'h8a18:	data_out=16'ha00;
17'h8a19:	data_out=16'h8a00;
17'h8a1a:	data_out=16'ha00;
17'h8a1b:	data_out=16'h89ac;
17'h8a1c:	data_out=16'ha00;
17'h8a1d:	data_out=16'ha00;
17'h8a1e:	data_out=16'h82cd;
17'h8a1f:	data_out=16'h89ff;
17'h8a20:	data_out=16'ha00;
17'h8a21:	data_out=16'ha00;
17'h8a22:	data_out=16'h8a00;
17'h8a23:	data_out=16'ha00;
17'h8a24:	data_out=16'ha00;
17'h8a25:	data_out=16'h8093;
17'h8a26:	data_out=16'ha00;
17'h8a27:	data_out=16'ha00;
17'h8a28:	data_out=16'ha00;
17'h8a29:	data_out=16'h8a00;
17'h8a2a:	data_out=16'ha00;
17'h8a2b:	data_out=16'h8a00;
17'h8a2c:	data_out=16'ha00;
17'h8a2d:	data_out=16'h8989;
17'h8a2e:	data_out=16'h88aa;
17'h8a2f:	data_out=16'h89ad;
17'h8a30:	data_out=16'ha00;
17'h8a31:	data_out=16'h984;
17'h8a32:	data_out=16'ha00;
17'h8a33:	data_out=16'h8a00;
17'h8a34:	data_out=16'ha00;
17'h8a35:	data_out=16'ha00;
17'h8a36:	data_out=16'ha00;
17'h8a37:	data_out=16'ha00;
17'h8a38:	data_out=16'h8f6;
17'h8a39:	data_out=16'h8a00;
17'h8a3a:	data_out=16'h8a00;
17'h8a3b:	data_out=16'ha00;
17'h8a3c:	data_out=16'h9af;
17'h8a3d:	data_out=16'ha00;
17'h8a3e:	data_out=16'ha00;
17'h8a3f:	data_out=16'ha00;
17'h8a40:	data_out=16'ha00;
17'h8a41:	data_out=16'ha00;
17'h8a42:	data_out=16'h73f;
17'h8a43:	data_out=16'h8a00;
17'h8a44:	data_out=16'ha00;
17'h8a45:	data_out=16'ha00;
17'h8a46:	data_out=16'ha00;
17'h8a47:	data_out=16'h8a00;
17'h8a48:	data_out=16'h89d7;
17'h8a49:	data_out=16'h73e;
17'h8a4a:	data_out=16'h87e9;
17'h8a4b:	data_out=16'h89c3;
17'h8a4c:	data_out=16'h438;
17'h8a4d:	data_out=16'h8a00;
17'h8a4e:	data_out=16'ha00;
17'h8a4f:	data_out=16'ha00;
17'h8a50:	data_out=16'h8a00;
17'h8a51:	data_out=16'ha00;
17'h8a52:	data_out=16'ha00;
17'h8a53:	data_out=16'h89c1;
17'h8a54:	data_out=16'ha00;
17'h8a55:	data_out=16'h85c1;
17'h8a56:	data_out=16'ha00;
17'h8a57:	data_out=16'ha00;
17'h8a58:	data_out=16'ha00;
17'h8a59:	data_out=16'ha00;
17'h8a5a:	data_out=16'h89fd;
17'h8a5b:	data_out=16'ha00;
17'h8a5c:	data_out=16'h887f;
17'h8a5d:	data_out=16'ha00;
17'h8a5e:	data_out=16'h89c7;
17'h8a5f:	data_out=16'ha00;
17'h8a60:	data_out=16'ha00;
17'h8a61:	data_out=16'ha00;
17'h8a62:	data_out=16'h89fe;
17'h8a63:	data_out=16'h8a00;
17'h8a64:	data_out=16'h87fe;
17'h8a65:	data_out=16'h8a00;
17'h8a66:	data_out=16'h8a00;
17'h8a67:	data_out=16'h8a00;
17'h8a68:	data_out=16'ha00;
17'h8a69:	data_out=16'ha00;
17'h8a6a:	data_out=16'ha00;
17'h8a6b:	data_out=16'h43c;
17'h8a6c:	data_out=16'ha00;
17'h8a6d:	data_out=16'h8a00;
17'h8a6e:	data_out=16'ha00;
17'h8a6f:	data_out=16'h89fe;
17'h8a70:	data_out=16'ha00;
17'h8a71:	data_out=16'ha00;
17'h8a72:	data_out=16'ha00;
17'h8a73:	data_out=16'ha00;
17'h8a74:	data_out=16'ha00;
17'h8a75:	data_out=16'ha00;
17'h8a76:	data_out=16'h8a00;
17'h8a77:	data_out=16'h81b9;
17'h8a78:	data_out=16'h8a00;
17'h8a79:	data_out=16'ha00;
17'h8a7a:	data_out=16'h89ff;
17'h8a7b:	data_out=16'ha00;
17'h8a7c:	data_out=16'ha00;
17'h8a7d:	data_out=16'h8a00;
17'h8a7e:	data_out=16'h8a00;
17'h8a7f:	data_out=16'ha00;
17'h8a80:	data_out=16'ha00;
17'h8a81:	data_out=16'ha00;
17'h8a82:	data_out=16'ha00;
17'h8a83:	data_out=16'h972;
17'h8a84:	data_out=16'ha00;
17'h8a85:	data_out=16'ha00;
17'h8a86:	data_out=16'h8a00;
17'h8a87:	data_out=16'h89ff;
17'h8a88:	data_out=16'ha00;
17'h8a89:	data_out=16'h8a00;
17'h8a8a:	data_out=16'ha00;
17'h8a8b:	data_out=16'h8a00;
17'h8a8c:	data_out=16'h428;
17'h8a8d:	data_out=16'ha00;
17'h8a8e:	data_out=16'ha00;
17'h8a8f:	data_out=16'ha00;
17'h8a90:	data_out=16'h8944;
17'h8a91:	data_out=16'ha00;
17'h8a92:	data_out=16'h82a3;
17'h8a93:	data_out=16'h84d;
17'h8a94:	data_out=16'h442;
17'h8a95:	data_out=16'ha00;
17'h8a96:	data_out=16'ha00;
17'h8a97:	data_out=16'h8a00;
17'h8a98:	data_out=16'ha00;
17'h8a99:	data_out=16'h8a00;
17'h8a9a:	data_out=16'ha00;
17'h8a9b:	data_out=16'h5bf;
17'h8a9c:	data_out=16'ha00;
17'h8a9d:	data_out=16'ha00;
17'h8a9e:	data_out=16'ha00;
17'h8a9f:	data_out=16'h80bf;
17'h8aa0:	data_out=16'ha00;
17'h8aa1:	data_out=16'ha00;
17'h8aa2:	data_out=16'h8a00;
17'h8aa3:	data_out=16'ha00;
17'h8aa4:	data_out=16'ha00;
17'h8aa5:	data_out=16'h8296;
17'h8aa6:	data_out=16'ha00;
17'h8aa7:	data_out=16'ha00;
17'h8aa8:	data_out=16'ha00;
17'h8aa9:	data_out=16'h8a00;
17'h8aaa:	data_out=16'ha00;
17'h8aab:	data_out=16'h8a00;
17'h8aac:	data_out=16'ha00;
17'h8aad:	data_out=16'h8a00;
17'h8aae:	data_out=16'h625;
17'h8aaf:	data_out=16'ha00;
17'h8ab0:	data_out=16'ha00;
17'h8ab1:	data_out=16'h73b;
17'h8ab2:	data_out=16'ha00;
17'h8ab3:	data_out=16'h51a;
17'h8ab4:	data_out=16'h23c;
17'h8ab5:	data_out=16'ha00;
17'h8ab6:	data_out=16'ha00;
17'h8ab7:	data_out=16'ha00;
17'h8ab8:	data_out=16'h92a;
17'h8ab9:	data_out=16'h981;
17'h8aba:	data_out=16'h8a00;
17'h8abb:	data_out=16'ha00;
17'h8abc:	data_out=16'h9fe;
17'h8abd:	data_out=16'ha00;
17'h8abe:	data_out=16'ha00;
17'h8abf:	data_out=16'ha00;
17'h8ac0:	data_out=16'ha00;
17'h8ac1:	data_out=16'ha00;
17'h8ac2:	data_out=16'h8593;
17'h8ac3:	data_out=16'h8a00;
17'h8ac4:	data_out=16'ha00;
17'h8ac5:	data_out=16'ha00;
17'h8ac6:	data_out=16'ha00;
17'h8ac7:	data_out=16'h8972;
17'h8ac8:	data_out=16'h89b8;
17'h8ac9:	data_out=16'h18c;
17'h8aca:	data_out=16'h93e;
17'h8acb:	data_out=16'h89fa;
17'h8acc:	data_out=16'h2b0;
17'h8acd:	data_out=16'h8a00;
17'h8ace:	data_out=16'ha00;
17'h8acf:	data_out=16'h940;
17'h8ad0:	data_out=16'h62a;
17'h8ad1:	data_out=16'ha00;
17'h8ad2:	data_out=16'ha00;
17'h8ad3:	data_out=16'ha00;
17'h8ad4:	data_out=16'ha00;
17'h8ad5:	data_out=16'h9bc;
17'h8ad6:	data_out=16'ha00;
17'h8ad7:	data_out=16'ha00;
17'h8ad8:	data_out=16'ha00;
17'h8ad9:	data_out=16'ha00;
17'h8ada:	data_out=16'h89fa;
17'h8adb:	data_out=16'ha00;
17'h8adc:	data_out=16'ha00;
17'h8add:	data_out=16'ha00;
17'h8ade:	data_out=16'ha00;
17'h8adf:	data_out=16'ha00;
17'h8ae0:	data_out=16'h9fe;
17'h8ae1:	data_out=16'ha00;
17'h8ae2:	data_out=16'h89ff;
17'h8ae3:	data_out=16'h3dc;
17'h8ae4:	data_out=16'h88a1;
17'h8ae5:	data_out=16'h8a00;
17'h8ae6:	data_out=16'h8a00;
17'h8ae7:	data_out=16'h8a00;
17'h8ae8:	data_out=16'ha00;
17'h8ae9:	data_out=16'ha00;
17'h8aea:	data_out=16'ha00;
17'h8aeb:	data_out=16'ha00;
17'h8aec:	data_out=16'ha00;
17'h8aed:	data_out=16'h4a5;
17'h8aee:	data_out=16'ha00;
17'h8aef:	data_out=16'h4c1;
17'h8af0:	data_out=16'ha00;
17'h8af1:	data_out=16'ha00;
17'h8af2:	data_out=16'ha00;
17'h8af3:	data_out=16'ha00;
17'h8af4:	data_out=16'ha00;
17'h8af5:	data_out=16'ha00;
17'h8af6:	data_out=16'h8a00;
17'h8af7:	data_out=16'h9f9;
17'h8af8:	data_out=16'h8a00;
17'h8af9:	data_out=16'ha00;
17'h8afa:	data_out=16'h819;
17'h8afb:	data_out=16'ha00;
17'h8afc:	data_out=16'ha00;
17'h8afd:	data_out=16'h87cb;
17'h8afe:	data_out=16'h8a00;
17'h8aff:	data_out=16'ha00;
17'h8b00:	data_out=16'ha00;
17'h8b01:	data_out=16'ha00;
17'h8b02:	data_out=16'ha00;
17'h8b03:	data_out=16'h848f;
17'h8b04:	data_out=16'ha00;
17'h8b05:	data_out=16'ha00;
17'h8b06:	data_out=16'h863c;
17'h8b07:	data_out=16'h8a00;
17'h8b08:	data_out=16'ha00;
17'h8b09:	data_out=16'h8a00;
17'h8b0a:	data_out=16'ha00;
17'h8b0b:	data_out=16'h8a00;
17'h8b0c:	data_out=16'h82cd;
17'h8b0d:	data_out=16'h85a5;
17'h8b0e:	data_out=16'h832;
17'h8b0f:	data_out=16'ha00;
17'h8b10:	data_out=16'h8a00;
17'h8b11:	data_out=16'h708;
17'h8b12:	data_out=16'h8971;
17'h8b13:	data_out=16'h8558;
17'h8b14:	data_out=16'h80bb;
17'h8b15:	data_out=16'ha00;
17'h8b16:	data_out=16'ha00;
17'h8b17:	data_out=16'h86ef;
17'h8b18:	data_out=16'h959;
17'h8b19:	data_out=16'h8a00;
17'h8b1a:	data_out=16'ha00;
17'h8b1b:	data_out=16'h88ae;
17'h8b1c:	data_out=16'ha00;
17'h8b1d:	data_out=16'h7c3;
17'h8b1e:	data_out=16'h15a;
17'h8b1f:	data_out=16'h5da;
17'h8b20:	data_out=16'h6d6;
17'h8b21:	data_out=16'h801;
17'h8b22:	data_out=16'h8a00;
17'h8b23:	data_out=16'h806;
17'h8b24:	data_out=16'h80d;
17'h8b25:	data_out=16'h8900;
17'h8b26:	data_out=16'h8543;
17'h8b27:	data_out=16'h55f;
17'h8b28:	data_out=16'h7b3;
17'h8b29:	data_out=16'h8916;
17'h8b2a:	data_out=16'h8172;
17'h8b2b:	data_out=16'h8a00;
17'h8b2c:	data_out=16'ha00;
17'h8b2d:	data_out=16'h8a00;
17'h8b2e:	data_out=16'h5b7;
17'h8b2f:	data_out=16'h8489;
17'h8b30:	data_out=16'ha00;
17'h8b31:	data_out=16'h8182;
17'h8b32:	data_out=16'ha00;
17'h8b33:	data_out=16'ha0;
17'h8b34:	data_out=16'h80a9;
17'h8b35:	data_out=16'ha00;
17'h8b36:	data_out=16'ha00;
17'h8b37:	data_out=16'ha00;
17'h8b38:	data_out=16'ha00;
17'h8b39:	data_out=16'h24a;
17'h8b3a:	data_out=16'h8a00;
17'h8b3b:	data_out=16'h9ff;
17'h8b3c:	data_out=16'ha00;
17'h8b3d:	data_out=16'ha00;
17'h8b3e:	data_out=16'h7b1;
17'h8b3f:	data_out=16'ha00;
17'h8b40:	data_out=16'h455;
17'h8b41:	data_out=16'ha00;
17'h8b42:	data_out=16'h8848;
17'h8b43:	data_out=16'h8a00;
17'h8b44:	data_out=16'ha00;
17'h8b45:	data_out=16'ha00;
17'h8b46:	data_out=16'h150;
17'h8b47:	data_out=16'h8a00;
17'h8b48:	data_out=16'h89fc;
17'h8b49:	data_out=16'h885c;
17'h8b4a:	data_out=16'h8157;
17'h8b4b:	data_out=16'h8a00;
17'h8b4c:	data_out=16'h891d;
17'h8b4d:	data_out=16'h8a00;
17'h8b4e:	data_out=16'h4fc;
17'h8b4f:	data_out=16'h89c9;
17'h8b50:	data_out=16'h449;
17'h8b51:	data_out=16'ha00;
17'h8b52:	data_out=16'h903;
17'h8b53:	data_out=16'h85d1;
17'h8b54:	data_out=16'ha00;
17'h8b55:	data_out=16'h8a4;
17'h8b56:	data_out=16'ha00;
17'h8b57:	data_out=16'ha00;
17'h8b58:	data_out=16'ha00;
17'h8b59:	data_out=16'ha00;
17'h8b5a:	data_out=16'h867e;
17'h8b5b:	data_out=16'ha00;
17'h8b5c:	data_out=16'h3da;
17'h8b5d:	data_out=16'ha00;
17'h8b5e:	data_out=16'h85c9;
17'h8b5f:	data_out=16'h523;
17'h8b60:	data_out=16'h8089;
17'h8b61:	data_out=16'ha00;
17'h8b62:	data_out=16'h8a00;
17'h8b63:	data_out=16'h16;
17'h8b64:	data_out=16'h88c6;
17'h8b65:	data_out=16'h8a00;
17'h8b66:	data_out=16'h8a00;
17'h8b67:	data_out=16'h8a00;
17'h8b68:	data_out=16'h7e0;
17'h8b69:	data_out=16'ha00;
17'h8b6a:	data_out=16'h84e;
17'h8b6b:	data_out=16'h9ff;
17'h8b6c:	data_out=16'ha00;
17'h8b6d:	data_out=16'h61;
17'h8b6e:	data_out=16'h84e;
17'h8b6f:	data_out=16'h83d0;
17'h8b70:	data_out=16'h840;
17'h8b71:	data_out=16'h9fe;
17'h8b72:	data_out=16'ha00;
17'h8b73:	data_out=16'ha00;
17'h8b74:	data_out=16'ha00;
17'h8b75:	data_out=16'ha00;
17'h8b76:	data_out=16'h8a00;
17'h8b77:	data_out=16'h8053;
17'h8b78:	data_out=16'h8a00;
17'h8b79:	data_out=16'ha00;
17'h8b7a:	data_out=16'h8077;
17'h8b7b:	data_out=16'h7b0;
17'h8b7c:	data_out=16'h7a9;
17'h8b7d:	data_out=16'h89fb;
17'h8b7e:	data_out=16'h8a00;
17'h8b7f:	data_out=16'ha00;
17'h8b80:	data_out=16'h20c;
17'h8b81:	data_out=16'h31f;
17'h8b82:	data_out=16'h249;
17'h8b83:	data_out=16'h88;
17'h8b84:	data_out=16'h81d8;
17'h8b85:	data_out=16'h80d5;
17'h8b86:	data_out=16'h80de;
17'h8b87:	data_out=16'h827b;
17'h8b88:	data_out=16'h25a;
17'h8b89:	data_out=16'h8287;
17'h8b8a:	data_out=16'hc1;
17'h8b8b:	data_out=16'h81c0;
17'h8b8c:	data_out=16'h825e;
17'h8b8d:	data_out=16'h14;
17'h8b8e:	data_out=16'h1b;
17'h8b8f:	data_out=16'h15f;
17'h8b90:	data_out=16'heb;
17'h8b91:	data_out=16'h8218;
17'h8b92:	data_out=16'h1a3;
17'h8b93:	data_out=16'h80f3;
17'h8b94:	data_out=16'h152;
17'h8b95:	data_out=16'h8018;
17'h8b96:	data_out=16'h8060;
17'h8b97:	data_out=16'h167;
17'h8b98:	data_out=16'h1e;
17'h8b99:	data_out=16'h84ca;
17'h8b9a:	data_out=16'h82eb;
17'h8b9b:	data_out=16'h154;
17'h8b9c:	data_out=16'h16;
17'h8b9d:	data_out=16'h1fd;
17'h8b9e:	data_out=16'h1d9;
17'h8b9f:	data_out=16'h81dc;
17'h8ba0:	data_out=16'h2a2;
17'h8ba1:	data_out=16'h17;
17'h8ba2:	data_out=16'h8102;
17'h8ba3:	data_out=16'h39;
17'h8ba4:	data_out=16'h39;
17'h8ba5:	data_out=16'h80d8;
17'h8ba6:	data_out=16'h81e8;
17'h8ba7:	data_out=16'h1f8;
17'h8ba8:	data_out=16'ha;
17'h8ba9:	data_out=16'h16;
17'h8baa:	data_out=16'h113;
17'h8bab:	data_out=16'h8189;
17'h8bac:	data_out=16'h8056;
17'h8bad:	data_out=16'h803d;
17'h8bae:	data_out=16'h1c3;
17'h8baf:	data_out=16'h2a2;
17'h8bb0:	data_out=16'h81d7;
17'h8bb1:	data_out=16'h811c;
17'h8bb2:	data_out=16'h8213;
17'h8bb3:	data_out=16'h193;
17'h8bb4:	data_out=16'h8118;
17'h8bb5:	data_out=16'h81a9;
17'h8bb6:	data_out=16'h4ae;
17'h8bb7:	data_out=16'h205;
17'h8bb8:	data_out=16'h128;
17'h8bb9:	data_out=16'h79;
17'h8bba:	data_out=16'h161;
17'h8bbb:	data_out=16'h815d;
17'h8bbc:	data_out=16'h329;
17'h8bbd:	data_out=16'h8084;
17'h8bbe:	data_out=16'h6;
17'h8bbf:	data_out=16'h8162;
17'h8bc0:	data_out=16'h80a2;
17'h8bc1:	data_out=16'h389;
17'h8bc2:	data_out=16'h802c;
17'h8bc3:	data_out=16'h81f0;
17'h8bc4:	data_out=16'h8139;
17'h8bc5:	data_out=16'h804e;
17'h8bc6:	data_out=16'h251;
17'h8bc7:	data_out=16'h804a;
17'h8bc8:	data_out=16'h801d;
17'h8bc9:	data_out=16'h8090;
17'h8bca:	data_out=16'h817c;
17'h8bcb:	data_out=16'h80;
17'h8bcc:	data_out=16'h80ba;
17'h8bcd:	data_out=16'h80c8;
17'h8bce:	data_out=16'h27e;
17'h8bcf:	data_out=16'h816d;
17'h8bd0:	data_out=16'h80c9;
17'h8bd1:	data_out=16'h8004;
17'h8bd2:	data_out=16'h20;
17'h8bd3:	data_out=16'h2a6;
17'h8bd4:	data_out=16'h35f;
17'h8bd5:	data_out=16'h123;
17'h8bd6:	data_out=16'h19a;
17'h8bd7:	data_out=16'h154;
17'h8bd8:	data_out=16'h213;
17'h8bd9:	data_out=16'h9a;
17'h8bda:	data_out=16'h271;
17'h8bdb:	data_out=16'h1bc;
17'h8bdc:	data_out=16'h103;
17'h8bdd:	data_out=16'h1e4;
17'h8bde:	data_out=16'h1ee;
17'h8bdf:	data_out=16'h169;
17'h8be0:	data_out=16'h8174;
17'h8be1:	data_out=16'h80bd;
17'h8be2:	data_out=16'hde;
17'h8be3:	data_out=16'h1a3;
17'h8be4:	data_out=16'h827c;
17'h8be5:	data_out=16'h8357;
17'h8be6:	data_out=16'h854f;
17'h8be7:	data_out=16'h8076;
17'h8be8:	data_out=16'hb;
17'h8be9:	data_out=16'h382;
17'h8bea:	data_out=16'h33;
17'h8beb:	data_out=16'h82de;
17'h8bec:	data_out=16'h4a1;
17'h8bed:	data_out=16'h19b;
17'h8bee:	data_out=16'h2e;
17'h8bef:	data_out=16'h80cf;
17'h8bf0:	data_out=16'h1d;
17'h8bf1:	data_out=16'h8017;
17'h8bf2:	data_out=16'h8114;
17'h8bf3:	data_out=16'h81bf;
17'h8bf4:	data_out=16'h81d8;
17'h8bf5:	data_out=16'h816f;
17'h8bf6:	data_out=16'h832f;
17'h8bf7:	data_out=16'h81de;
17'h8bf8:	data_out=16'h8394;
17'h8bf9:	data_out=16'h245;
17'h8bfa:	data_out=16'h18d;
17'h8bfb:	data_out=16'h8;
17'h8bfc:	data_out=16'hf0;
17'h8bfd:	data_out=16'h81e7;
17'h8bfe:	data_out=16'h829a;
17'h8bff:	data_out=16'h81c1;
17'h8c00:	data_out=16'h5f;
17'h8c01:	data_out=16'h9a;
17'h8c02:	data_out=16'h74;
17'h8c03:	data_out=16'h75;
17'h8c04:	data_out=16'h96;
17'h8c05:	data_out=16'h9a;
17'h8c06:	data_out=16'h2;
17'h8c07:	data_out=16'h6b;
17'h8c08:	data_out=16'h3a;
17'h8c09:	data_out=16'h8008;
17'h8c0a:	data_out=16'hb2;
17'h8c0b:	data_out=16'h4;
17'h8c0c:	data_out=16'h9e;
17'h8c0d:	data_out=16'h53;
17'h8c0e:	data_out=16'h7;
17'h8c0f:	data_out=16'h5f;
17'h8c10:	data_out=16'h8007;
17'h8c11:	data_out=16'h94;
17'h8c12:	data_out=16'h6d;
17'h8c13:	data_out=16'h49;
17'h8c14:	data_out=16'h8a;
17'h8c15:	data_out=16'h38;
17'h8c16:	data_out=16'h5e;
17'h8c17:	data_out=16'h8f;
17'h8c18:	data_out=16'ha;
17'h8c19:	data_out=16'h2b;
17'h8c1a:	data_out=16'h7f;
17'h8c1b:	data_out=16'h39;
17'h8c1c:	data_out=16'hae;
17'h8c1d:	data_out=16'hfd;
17'h8c1e:	data_out=16'h85;
17'h8c1f:	data_out=16'h3b;
17'h8c20:	data_out=16'hd8;
17'h8c21:	data_out=16'hd;
17'h8c22:	data_out=16'h53;
17'h8c23:	data_out=16'h13;
17'h8c24:	data_out=16'h15;
17'h8c25:	data_out=16'h5a;
17'h8c26:	data_out=16'h801f;
17'h8c27:	data_out=16'he9;
17'h8c28:	data_out=16'h16;
17'h8c29:	data_out=16'h41;
17'h8c2a:	data_out=16'h3d;
17'h8c2b:	data_out=16'h4d;
17'h8c2c:	data_out=16'h6f;
17'h8c2d:	data_out=16'h33;
17'h8c2e:	data_out=16'h42;
17'h8c2f:	data_out=16'h98;
17'h8c30:	data_out=16'h9d;
17'h8c31:	data_out=16'h9e;
17'h8c32:	data_out=16'hac;
17'h8c33:	data_out=16'h98;
17'h8c34:	data_out=16'h58;
17'h8c35:	data_out=16'ha1;
17'h8c36:	data_out=16'h4c;
17'h8c37:	data_out=16'h95;
17'h8c38:	data_out=16'h67;
17'h8c39:	data_out=16'h29;
17'h8c3a:	data_out=16'h84;
17'h8c3b:	data_out=16'h65;
17'h8c3c:	data_out=16'h90;
17'h8c3d:	data_out=16'h65;
17'h8c3e:	data_out=16'h16;
17'h8c3f:	data_out=16'h6a;
17'h8c40:	data_out=16'h8d;
17'h8c41:	data_out=16'h66;
17'h8c42:	data_out=16'h51;
17'h8c43:	data_out=16'h8009;
17'h8c44:	data_out=16'h57;
17'h8c45:	data_out=16'h16;
17'h8c46:	data_out=16'h6d;
17'h8c47:	data_out=16'h5b;
17'h8c48:	data_out=16'h2d;
17'h8c49:	data_out=16'h67;
17'h8c4a:	data_out=16'h72;
17'h8c4b:	data_out=16'ha3;
17'h8c4c:	data_out=16'h60;
17'h8c4d:	data_out=16'h6e;
17'h8c4e:	data_out=16'h6c;
17'h8c4f:	data_out=16'h69;
17'h8c50:	data_out=16'h68;
17'h8c51:	data_out=16'h35;
17'h8c52:	data_out=16'h25;
17'h8c53:	data_out=16'h100;
17'h8c54:	data_out=16'hac;
17'h8c55:	data_out=16'h28;
17'h8c56:	data_out=16'h81;
17'h8c57:	data_out=16'h3e;
17'h8c58:	data_out=16'h6d;
17'h8c59:	data_out=16'h67;
17'h8c5a:	data_out=16'h4d;
17'h8c5b:	data_out=16'h68;
17'h8c5c:	data_out=16'h96;
17'h8c5d:	data_out=16'h83;
17'h8c5e:	data_out=16'h93;
17'h8c5f:	data_out=16'h33;
17'h8c60:	data_out=16'h26;
17'h8c61:	data_out=16'h97;
17'h8c62:	data_out=16'h2d;
17'h8c63:	data_out=16'h92;
17'h8c64:	data_out=16'h5a;
17'h8c65:	data_out=16'h79;
17'h8c66:	data_out=16'h24;
17'h8c67:	data_out=16'h35;
17'h8c68:	data_out=16'he;
17'h8c69:	data_out=16'h51;
17'h8c6a:	data_out=16'h4;
17'h8c6b:	data_out=16'h7f;
17'h8c6c:	data_out=16'h11a;
17'h8c6d:	data_out=16'h88;
17'h8c6e:	data_out=16'h11;
17'h8c6f:	data_out=16'hae;
17'h8c70:	data_out=16'h6;
17'h8c71:	data_out=16'h2b;
17'h8c72:	data_out=16'h6e;
17'h8c73:	data_out=16'h76;
17'h8c74:	data_out=16'h98;
17'h8c75:	data_out=16'h52;
17'h8c76:	data_out=16'h2f;
17'h8c77:	data_out=16'h2d;
17'h8c78:	data_out=16'h0;
17'h8c79:	data_out=16'h4b;
17'h8c7a:	data_out=16'h8a;
17'h8c7b:	data_out=16'ha;
17'h8c7c:	data_out=16'h15;
17'h8c7d:	data_out=16'h7;
17'h8c7e:	data_out=16'h801d;
17'h8c7f:	data_out=16'h59;
17'h8c80:	data_out=16'h5f7;
17'h8c81:	data_out=16'h758;
17'h8c82:	data_out=16'h25f;
17'h8c83:	data_out=16'h42c;
17'h8c84:	data_out=16'h80d6;
17'h8c85:	data_out=16'h8013;
17'h8c86:	data_out=16'h8303;
17'h8c87:	data_out=16'h1cf;
17'h8c88:	data_out=16'h2e7;
17'h8c89:	data_out=16'h99;
17'h8c8a:	data_out=16'h2ab;
17'h8c8b:	data_out=16'ha1;
17'h8c8c:	data_out=16'h8075;
17'h8c8d:	data_out=16'h3b1;
17'h8c8e:	data_out=16'h10;
17'h8c8f:	data_out=16'h42d;
17'h8c90:	data_out=16'h33a;
17'h8c91:	data_out=16'h810e;
17'h8c92:	data_out=16'h553;
17'h8c93:	data_out=16'h38b;
17'h8c94:	data_out=16'h2cf;
17'h8c95:	data_out=16'heb;
17'h8c96:	data_out=16'h221;
17'h8c97:	data_out=16'h40f;
17'h8c98:	data_out=16'ha7;
17'h8c99:	data_out=16'h8110;
17'h8c9a:	data_out=16'h80a1;
17'h8c9b:	data_out=16'h58c;
17'h8c9c:	data_out=16'h8038;
17'h8c9d:	data_out=16'h5da;
17'h8c9e:	data_out=16'h4fc;
17'h8c9f:	data_out=16'h82a5;
17'h8ca0:	data_out=16'h8c9;
17'h8ca1:	data_out=16'h20;
17'h8ca2:	data_out=16'h51e;
17'h8ca3:	data_out=16'h80e2;
17'h8ca4:	data_out=16'h80d8;
17'h8ca5:	data_out=16'h22e;
17'h8ca6:	data_out=16'h810e;
17'h8ca7:	data_out=16'h606;
17'h8ca8:	data_out=16'h16;
17'h8ca9:	data_out=16'h4d7;
17'h8caa:	data_out=16'h7cf;
17'h8cab:	data_out=16'h121;
17'h8cac:	data_out=16'h187;
17'h8cad:	data_out=16'h650;
17'h8cae:	data_out=16'h652;
17'h8caf:	data_out=16'ha00;
17'h8cb0:	data_out=16'h8084;
17'h8cb1:	data_out=16'h2ed;
17'h8cb2:	data_out=16'h8045;
17'h8cb3:	data_out=16'h325;
17'h8cb4:	data_out=16'h37f;
17'h8cb5:	data_out=16'h816d;
17'h8cb6:	data_out=16'h65d;
17'h8cb7:	data_out=16'h258;
17'h8cb8:	data_out=16'h8035;
17'h8cb9:	data_out=16'h3ae;
17'h8cba:	data_out=16'h73a;
17'h8cbb:	data_out=16'h813c;
17'h8cbc:	data_out=16'h410;
17'h8cbd:	data_out=16'h1e8;
17'h8cbe:	data_out=16'h1d;
17'h8cbf:	data_out=16'h80b9;
17'h8cc0:	data_out=16'h801c;
17'h8cc1:	data_out=16'h259;
17'h8cc2:	data_out=16'h7a4;
17'h8cc3:	data_out=16'h8486;
17'h8cc4:	data_out=16'h8083;
17'h8cc5:	data_out=16'h8020;
17'h8cc6:	data_out=16'h2c3;
17'h8cc7:	data_out=16'h355;
17'h8cc8:	data_out=16'h56e;
17'h8cc9:	data_out=16'h194;
17'h8cca:	data_out=16'h384;
17'h8ccb:	data_out=16'h816;
17'h8ccc:	data_out=16'h5cd;
17'h8ccd:	data_out=16'h58d;
17'h8cce:	data_out=16'h6a8;
17'h8ccf:	data_out=16'h4b7;
17'h8cd0:	data_out=16'h80de;
17'h8cd1:	data_out=16'h81a2;
17'h8cd2:	data_out=16'h80ee;
17'h8cd3:	data_out=16'h7c4;
17'h8cd4:	data_out=16'ha00;
17'h8cd5:	data_out=16'h801d;
17'h8cd6:	data_out=16'h804d;
17'h8cd7:	data_out=16'h8016;
17'h8cd8:	data_out=16'h84;
17'h8cd9:	data_out=16'hac;
17'h8cda:	data_out=16'h443;
17'h8cdb:	data_out=16'h82aa;
17'h8cdc:	data_out=16'h38d;
17'h8cdd:	data_out=16'h86e;
17'h8cde:	data_out=16'ha00;
17'h8cdf:	data_out=16'h439;
17'h8ce0:	data_out=16'h1ab;
17'h8ce1:	data_out=16'h8128;
17'h8ce2:	data_out=16'h22b;
17'h8ce3:	data_out=16'h325;
17'h8ce4:	data_out=16'h12a;
17'h8ce5:	data_out=16'h1a3;
17'h8ce6:	data_out=16'h8140;
17'h8ce7:	data_out=16'h325;
17'h8ce8:	data_out=16'h12;
17'h8ce9:	data_out=16'h35c;
17'h8cea:	data_out=16'hd;
17'h8ceb:	data_out=16'h8074;
17'h8cec:	data_out=16'ha00;
17'h8ced:	data_out=16'h342;
17'h8cee:	data_out=16'h4;
17'h8cef:	data_out=16'h25f;
17'h8cf0:	data_out=16'h17;
17'h8cf1:	data_out=16'h2d8;
17'h8cf2:	data_out=16'h802b;
17'h8cf3:	data_out=16'hbe;
17'h8cf4:	data_out=16'h8088;
17'h8cf5:	data_out=16'h8389;
17'h8cf6:	data_out=16'h96;
17'h8cf7:	data_out=16'h8116;
17'h8cf8:	data_out=16'h83fc;
17'h8cf9:	data_out=16'h714;
17'h8cfa:	data_out=16'h313;
17'h8cfb:	data_out=16'h1c;
17'h8cfc:	data_out=16'h1b4;
17'h8cfd:	data_out=16'h83b5;
17'h8cfe:	data_out=16'h8181;
17'h8cff:	data_out=16'h8033;
17'h8d00:	data_out=16'ha00;
17'h8d01:	data_out=16'ha00;
17'h8d02:	data_out=16'h6e9;
17'h8d03:	data_out=16'ha00;
17'h8d04:	data_out=16'h2d;
17'h8d05:	data_out=16'h293;
17'h8d06:	data_out=16'h8700;
17'h8d07:	data_out=16'h948;
17'h8d08:	data_out=16'ha00;
17'h8d09:	data_out=16'h675;
17'h8d0a:	data_out=16'h9f6;
17'h8d0b:	data_out=16'h576;
17'h8d0c:	data_out=16'h259;
17'h8d0d:	data_out=16'h98f;
17'h8d0e:	data_out=16'h808f;
17'h8d0f:	data_out=16'ha00;
17'h8d10:	data_out=16'ha00;
17'h8d11:	data_out=16'h1fa;
17'h8d12:	data_out=16'ha00;
17'h8d13:	data_out=16'ha00;
17'h8d14:	data_out=16'h70c;
17'h8d15:	data_out=16'h202;
17'h8d16:	data_out=16'h79f;
17'h8d17:	data_out=16'ha00;
17'h8d18:	data_out=16'he4;
17'h8d19:	data_out=16'h80ed;
17'h8d1a:	data_out=16'h18;
17'h8d1b:	data_out=16'ha00;
17'h8d1c:	data_out=16'h20b;
17'h8d1d:	data_out=16'ha00;
17'h8d1e:	data_out=16'ha00;
17'h8d1f:	data_out=16'h8756;
17'h8d20:	data_out=16'ha00;
17'h8d21:	data_out=16'h8091;
17'h8d22:	data_out=16'ha00;
17'h8d23:	data_out=16'h8316;
17'h8d24:	data_out=16'h8333;
17'h8d25:	data_out=16'h927;
17'h8d26:	data_out=16'h403;
17'h8d27:	data_out=16'ha00;
17'h8d28:	data_out=16'h8098;
17'h8d29:	data_out=16'ha00;
17'h8d2a:	data_out=16'ha00;
17'h8d2b:	data_out=16'h990;
17'h8d2c:	data_out=16'h572;
17'h8d2d:	data_out=16'ha00;
17'h8d2e:	data_out=16'ha00;
17'h8d2f:	data_out=16'ha00;
17'h8d30:	data_out=16'h182;
17'h8d31:	data_out=16'h9f6;
17'h8d32:	data_out=16'h257;
17'h8d33:	data_out=16'h8b9;
17'h8d34:	data_out=16'ha00;
17'h8d35:	data_out=16'h12b;
17'h8d36:	data_out=16'ha00;
17'h8d37:	data_out=16'h6c4;
17'h8d38:	data_out=16'h40c;
17'h8d39:	data_out=16'ha00;
17'h8d3a:	data_out=16'ha00;
17'h8d3b:	data_out=16'h17b;
17'h8d3c:	data_out=16'h9cd;
17'h8d3d:	data_out=16'ha00;
17'h8d3e:	data_out=16'h8098;
17'h8d3f:	data_out=16'h290;
17'h8d40:	data_out=16'h2ce;
17'h8d41:	data_out=16'h4d8;
17'h8d42:	data_out=16'ha00;
17'h8d43:	data_out=16'h8a00;
17'h8d44:	data_out=16'h367;
17'h8d45:	data_out=16'h22f;
17'h8d46:	data_out=16'h885;
17'h8d47:	data_out=16'ha00;
17'h8d48:	data_out=16'ha00;
17'h8d49:	data_out=16'h7d2;
17'h8d4a:	data_out=16'ha00;
17'h8d4b:	data_out=16'ha00;
17'h8d4c:	data_out=16'ha00;
17'h8d4d:	data_out=16'ha00;
17'h8d4e:	data_out=16'ha00;
17'h8d4f:	data_out=16'ha00;
17'h8d50:	data_out=16'h8255;
17'h8d51:	data_out=16'h8644;
17'h8d52:	data_out=16'h83ae;
17'h8d53:	data_out=16'ha00;
17'h8d54:	data_out=16'ha00;
17'h8d55:	data_out=16'h81f3;
17'h8d56:	data_out=16'h112;
17'h8d57:	data_out=16'h1d0;
17'h8d58:	data_out=16'h14f;
17'h8d59:	data_out=16'h520;
17'h8d5a:	data_out=16'h9ed;
17'h8d5b:	data_out=16'h8531;
17'h8d5c:	data_out=16'h9fb;
17'h8d5d:	data_out=16'ha00;
17'h8d5e:	data_out=16'ha00;
17'h8d5f:	data_out=16'ha00;
17'h8d60:	data_out=16'h79c;
17'h8d61:	data_out=16'h6;
17'h8d62:	data_out=16'h445;
17'h8d63:	data_out=16'h8a9;
17'h8d64:	data_out=16'h71b;
17'h8d65:	data_out=16'h9ff;
17'h8d66:	data_out=16'h8315;
17'h8d67:	data_out=16'h90c;
17'h8d68:	data_out=16'h8095;
17'h8d69:	data_out=16'ha00;
17'h8d6a:	data_out=16'h8094;
17'h8d6b:	data_out=16'h184;
17'h8d6c:	data_out=16'ha00;
17'h8d6d:	data_out=16'h90e;
17'h8d6e:	data_out=16'h8094;
17'h8d6f:	data_out=16'h9f8;
17'h8d70:	data_out=16'h8092;
17'h8d71:	data_out=16'h65c;
17'h8d72:	data_out=16'h3bb;
17'h8d73:	data_out=16'h57e;
17'h8d74:	data_out=16'h16c;
17'h8d75:	data_out=16'h8927;
17'h8d76:	data_out=16'h188;
17'h8d77:	data_out=16'h813d;
17'h8d78:	data_out=16'h8a00;
17'h8d79:	data_out=16'ha00;
17'h8d7a:	data_out=16'h806;
17'h8d7b:	data_out=16'h8098;
17'h8d7c:	data_out=16'h397;
17'h8d7d:	data_out=16'h893f;
17'h8d7e:	data_out=16'h228;
17'h8d7f:	data_out=16'h1af;
17'h8d80:	data_out=16'h9f5;
17'h8d81:	data_out=16'ha00;
17'h8d82:	data_out=16'h9fa;
17'h8d83:	data_out=16'h94c;
17'h8d84:	data_out=16'h87a5;
17'h8d85:	data_out=16'h9f7;
17'h8d86:	data_out=16'h864d;
17'h8d87:	data_out=16'h13e;
17'h8d88:	data_out=16'ha00;
17'h8d89:	data_out=16'h89f5;
17'h8d8a:	data_out=16'h272;
17'h8d8b:	data_out=16'ha00;
17'h8d8c:	data_out=16'h206;
17'h8d8d:	data_out=16'h878;
17'h8d8e:	data_out=16'h83a5;
17'h8d8f:	data_out=16'ha00;
17'h8d90:	data_out=16'h989;
17'h8d91:	data_out=16'h2fd;
17'h8d92:	data_out=16'ha00;
17'h8d93:	data_out=16'h91f;
17'h8d94:	data_out=16'ha00;
17'h8d95:	data_out=16'h8746;
17'h8d96:	data_out=16'h8138;
17'h8d97:	data_out=16'ha00;
17'h8d98:	data_out=16'h8033;
17'h8d99:	data_out=16'h44d;
17'h8d9a:	data_out=16'h8182;
17'h8d9b:	data_out=16'h9fb;
17'h8d9c:	data_out=16'h9b4;
17'h8d9d:	data_out=16'ha00;
17'h8d9e:	data_out=16'ha00;
17'h8d9f:	data_out=16'h886b;
17'h8da0:	data_out=16'ha00;
17'h8da1:	data_out=16'h8382;
17'h8da2:	data_out=16'h9c5;
17'h8da3:	data_out=16'h8a00;
17'h8da4:	data_out=16'h8a00;
17'h8da5:	data_out=16'h81e4;
17'h8da6:	data_out=16'h8a00;
17'h8da7:	data_out=16'ha00;
17'h8da8:	data_out=16'h8334;
17'h8da9:	data_out=16'h9e8;
17'h8daa:	data_out=16'ha00;
17'h8dab:	data_out=16'ha00;
17'h8dac:	data_out=16'h844c;
17'h8dad:	data_out=16'h9fb;
17'h8dae:	data_out=16'ha00;
17'h8daf:	data_out=16'ha00;
17'h8db0:	data_out=16'h8528;
17'h8db1:	data_out=16'h9ff;
17'h8db2:	data_out=16'h856e;
17'h8db3:	data_out=16'ha00;
17'h8db4:	data_out=16'ha00;
17'h8db5:	data_out=16'h97a;
17'h8db6:	data_out=16'ha00;
17'h8db7:	data_out=16'h9fc;
17'h8db8:	data_out=16'ha00;
17'h8db9:	data_out=16'ha00;
17'h8dba:	data_out=16'h93d;
17'h8dbb:	data_out=16'h84fe;
17'h8dbc:	data_out=16'h9fa;
17'h8dbd:	data_out=16'h68d;
17'h8dbe:	data_out=16'h8331;
17'h8dbf:	data_out=16'h9f6;
17'h8dc0:	data_out=16'h84e3;
17'h8dc1:	data_out=16'h9f7;
17'h8dc2:	data_out=16'h93e;
17'h8dc3:	data_out=16'h89fd;
17'h8dc4:	data_out=16'h65a;
17'h8dc5:	data_out=16'h8782;
17'h8dc6:	data_out=16'h9ea;
17'h8dc7:	data_out=16'h8e;
17'h8dc8:	data_out=16'ha00;
17'h8dc9:	data_out=16'h845f;
17'h8dca:	data_out=16'ha00;
17'h8dcb:	data_out=16'h9ff;
17'h8dcc:	data_out=16'h818;
17'h8dcd:	data_out=16'ha00;
17'h8dce:	data_out=16'ha00;
17'h8dcf:	data_out=16'h573;
17'h8dd0:	data_out=16'h8898;
17'h8dd1:	data_out=16'h89f7;
17'h8dd2:	data_out=16'h8a00;
17'h8dd3:	data_out=16'ha00;
17'h8dd4:	data_out=16'ha00;
17'h8dd5:	data_out=16'h429;
17'h8dd6:	data_out=16'h8a00;
17'h8dd7:	data_out=16'h8a00;
17'h8dd8:	data_out=16'h709;
17'h8dd9:	data_out=16'h89f2;
17'h8dda:	data_out=16'h9ff;
17'h8ddb:	data_out=16'h80b1;
17'h8ddc:	data_out=16'ha00;
17'h8ddd:	data_out=16'ha00;
17'h8dde:	data_out=16'ha00;
17'h8ddf:	data_out=16'ha00;
17'h8de0:	data_out=16'h89fe;
17'h8de1:	data_out=16'hbd;
17'h8de2:	data_out=16'h9f8;
17'h8de3:	data_out=16'ha00;
17'h8de4:	data_out=16'h914;
17'h8de5:	data_out=16'ha00;
17'h8de6:	data_out=16'h26b;
17'h8de7:	data_out=16'ha00;
17'h8de8:	data_out=16'h8376;
17'h8de9:	data_out=16'h9b9;
17'h8dea:	data_out=16'h83ce;
17'h8deb:	data_out=16'h40;
17'h8dec:	data_out=16'h9f6;
17'h8ded:	data_out=16'ha00;
17'h8dee:	data_out=16'h83ce;
17'h8def:	data_out=16'h9fc;
17'h8df0:	data_out=16'h83b8;
17'h8df1:	data_out=16'ha00;
17'h8df2:	data_out=16'h89f2;
17'h8df3:	data_out=16'hb3;
17'h8df4:	data_out=16'h8567;
17'h8df5:	data_out=16'h8d8;
17'h8df6:	data_out=16'ha00;
17'h8df7:	data_out=16'h87e2;
17'h8df8:	data_out=16'h89ff;
17'h8df9:	data_out=16'h9fe;
17'h8dfa:	data_out=16'ha00;
17'h8dfb:	data_out=16'h832f;
17'h8dfc:	data_out=16'h94e;
17'h8dfd:	data_out=16'h81b5;
17'h8dfe:	data_out=16'h89fb;
17'h8dff:	data_out=16'h89fe;
17'h8e00:	data_out=16'h176;
17'h8e01:	data_out=16'h9fc;
17'h8e02:	data_out=16'h7ed;
17'h8e03:	data_out=16'h8a00;
17'h8e04:	data_out=16'h88d0;
17'h8e05:	data_out=16'h80a7;
17'h8e06:	data_out=16'h89e9;
17'h8e07:	data_out=16'h8501;
17'h8e08:	data_out=16'h83e2;
17'h8e09:	data_out=16'h89ef;
17'h8e0a:	data_out=16'h89ef;
17'h8e0b:	data_out=16'h19c;
17'h8e0c:	data_out=16'h88c0;
17'h8e0d:	data_out=16'h82f8;
17'h8e0e:	data_out=16'h8272;
17'h8e0f:	data_out=16'h9ea;
17'h8e10:	data_out=16'h89ff;
17'h8e11:	data_out=16'h8501;
17'h8e12:	data_out=16'h9ed;
17'h8e13:	data_out=16'h8a00;
17'h8e14:	data_out=16'h6fd;
17'h8e15:	data_out=16'h8a00;
17'h8e16:	data_out=16'h8a00;
17'h8e17:	data_out=16'h877;
17'h8e18:	data_out=16'h81b2;
17'h8e19:	data_out=16'h8dd;
17'h8e1a:	data_out=16'h3e8;
17'h8e1b:	data_out=16'h7dc;
17'h8e1c:	data_out=16'h8043;
17'h8e1d:	data_out=16'ha00;
17'h8e1e:	data_out=16'h928;
17'h8e1f:	data_out=16'h89e1;
17'h8e20:	data_out=16'h9f8;
17'h8e21:	data_out=16'h822c;
17'h8e22:	data_out=16'h9fc;
17'h8e23:	data_out=16'h89fe;
17'h8e24:	data_out=16'h89fe;
17'h8e25:	data_out=16'h89f6;
17'h8e26:	data_out=16'h8a00;
17'h8e27:	data_out=16'h9f4;
17'h8e28:	data_out=16'h81e5;
17'h8e29:	data_out=16'h7b3;
17'h8e2a:	data_out=16'h9d6;
17'h8e2b:	data_out=16'ha00;
17'h8e2c:	data_out=16'h8a00;
17'h8e2d:	data_out=16'h9fb;
17'h8e2e:	data_out=16'h9f6;
17'h8e2f:	data_out=16'h9f3;
17'h8e30:	data_out=16'h4b2;
17'h8e31:	data_out=16'h47a;
17'h8e32:	data_out=16'h311;
17'h8e33:	data_out=16'h9e8;
17'h8e34:	data_out=16'h9f9;
17'h8e35:	data_out=16'h86eb;
17'h8e36:	data_out=16'h9de;
17'h8e37:	data_out=16'h7ef;
17'h8e38:	data_out=16'ha00;
17'h8e39:	data_out=16'h9e5;
17'h8e3a:	data_out=16'h4d6;
17'h8e3b:	data_out=16'h89f4;
17'h8e3c:	data_out=16'h8bd;
17'h8e3d:	data_out=16'h85a3;
17'h8e3e:	data_out=16'h81e4;
17'h8e3f:	data_out=16'h80fa;
17'h8e40:	data_out=16'h884d;
17'h8e41:	data_out=16'h34d;
17'h8e42:	data_out=16'h8a00;
17'h8e43:	data_out=16'h89fc;
17'h8e44:	data_out=16'h89af;
17'h8e45:	data_out=16'h8a00;
17'h8e46:	data_out=16'h9dd;
17'h8e47:	data_out=16'h8725;
17'h8e48:	data_out=16'h9fd;
17'h8e49:	data_out=16'h89fd;
17'h8e4a:	data_out=16'h9fb;
17'h8e4b:	data_out=16'h496;
17'h8e4c:	data_out=16'h2e1;
17'h8e4d:	data_out=16'h9ff;
17'h8e4e:	data_out=16'h9fd;
17'h8e4f:	data_out=16'h84b3;
17'h8e50:	data_out=16'h89f7;
17'h8e51:	data_out=16'h8a00;
17'h8e52:	data_out=16'h89fb;
17'h8e53:	data_out=16'ha00;
17'h8e54:	data_out=16'h9f1;
17'h8e55:	data_out=16'h8a00;
17'h8e56:	data_out=16'h8a00;
17'h8e57:	data_out=16'h89fe;
17'h8e58:	data_out=16'h8767;
17'h8e59:	data_out=16'h89dd;
17'h8e5a:	data_out=16'h9e6;
17'h8e5b:	data_out=16'h8186;
17'h8e5c:	data_out=16'h9e7;
17'h8e5d:	data_out=16'h9f3;
17'h8e5e:	data_out=16'h9f1;
17'h8e5f:	data_out=16'h9ff;
17'h8e60:	data_out=16'h8a00;
17'h8e61:	data_out=16'h8644;
17'h8e62:	data_out=16'h8ca;
17'h8e63:	data_out=16'h9f0;
17'h8e64:	data_out=16'hcd;
17'h8e65:	data_out=16'h85ad;
17'h8e66:	data_out=16'h84e6;
17'h8e67:	data_out=16'ha00;
17'h8e68:	data_out=16'h8210;
17'h8e69:	data_out=16'h89e7;
17'h8e6a:	data_out=16'h82c2;
17'h8e6b:	data_out=16'h8446;
17'h8e6c:	data_out=16'h9cf;
17'h8e6d:	data_out=16'h9ed;
17'h8e6e:	data_out=16'h82c0;
17'h8e6f:	data_out=16'h8c;
17'h8e70:	data_out=16'h8292;
17'h8e71:	data_out=16'h9f9;
17'h8e72:	data_out=16'h85f2;
17'h8e73:	data_out=16'h148;
17'h8e74:	data_out=16'h4b3;
17'h8e75:	data_out=16'h64e;
17'h8e76:	data_out=16'h5bd;
17'h8e77:	data_out=16'h89fd;
17'h8e78:	data_out=16'h89ea;
17'h8e79:	data_out=16'h969;
17'h8e7a:	data_out=16'h9e9;
17'h8e7b:	data_out=16'h81e3;
17'h8e7c:	data_out=16'ha00;
17'h8e7d:	data_out=16'h8954;
17'h8e7e:	data_out=16'h89fb;
17'h8e7f:	data_out=16'h871d;
17'h8e80:	data_out=16'h12;
17'h8e81:	data_out=16'h9d1;
17'h8e82:	data_out=16'h89ff;
17'h8e83:	data_out=16'h8a00;
17'h8e84:	data_out=16'h101;
17'h8e85:	data_out=16'h89ff;
17'h8e86:	data_out=16'h89ea;
17'h8e87:	data_out=16'h89fc;
17'h8e88:	data_out=16'h8083;
17'h8e89:	data_out=16'h89df;
17'h8e8a:	data_out=16'h89e0;
17'h8e8b:	data_out=16'h857d;
17'h8e8c:	data_out=16'h89f1;
17'h8e8d:	data_out=16'h8a00;
17'h8e8e:	data_out=16'h8153;
17'h8e8f:	data_out=16'h899b;
17'h8e90:	data_out=16'h315;
17'h8e91:	data_out=16'h8509;
17'h8e92:	data_out=16'h812a;
17'h8e93:	data_out=16'h8a00;
17'h8e94:	data_out=16'h858d;
17'h8e95:	data_out=16'h89ff;
17'h8e96:	data_out=16'h89ff;
17'h8e97:	data_out=16'h8573;
17'h8e98:	data_out=16'h848e;
17'h8e99:	data_out=16'ha00;
17'h8e9a:	data_out=16'h82e9;
17'h8e9b:	data_out=16'h87c8;
17'h8e9c:	data_out=16'h8a00;
17'h8e9d:	data_out=16'h68c;
17'h8e9e:	data_out=16'h8111;
17'h8e9f:	data_out=16'h89f2;
17'h8ea0:	data_out=16'h9d0;
17'h8ea1:	data_out=16'h810b;
17'h8ea2:	data_out=16'h9fe;
17'h8ea3:	data_out=16'h89ed;
17'h8ea4:	data_out=16'h89ed;
17'h8ea5:	data_out=16'h89e7;
17'h8ea6:	data_out=16'h8a00;
17'h8ea7:	data_out=16'h9ba;
17'h8ea8:	data_out=16'h80c8;
17'h8ea9:	data_out=16'h8278;
17'h8eaa:	data_out=16'h832c;
17'h8eab:	data_out=16'ha00;
17'h8eac:	data_out=16'h89ff;
17'h8ead:	data_out=16'h9f2;
17'h8eae:	data_out=16'h8f3;
17'h8eaf:	data_out=16'h9c9;
17'h8eb0:	data_out=16'h8121;
17'h8eb1:	data_out=16'h8a00;
17'h8eb2:	data_out=16'h825f;
17'h8eb3:	data_out=16'h146;
17'h8eb4:	data_out=16'h2a5;
17'h8eb5:	data_out=16'h88e5;
17'h8eb6:	data_out=16'h9c4;
17'h8eb7:	data_out=16'h8a00;
17'h8eb8:	data_out=16'h9f4;
17'h8eb9:	data_out=16'h5a9;
17'h8eba:	data_out=16'hf5;
17'h8ebb:	data_out=16'h89fd;
17'h8ebc:	data_out=16'h4c4;
17'h8ebd:	data_out=16'h8415;
17'h8ebe:	data_out=16'h80c9;
17'h8ebf:	data_out=16'h89ff;
17'h8ec0:	data_out=16'h872c;
17'h8ec1:	data_out=16'h89ff;
17'h8ec2:	data_out=16'h8a00;
17'h8ec3:	data_out=16'h8a00;
17'h8ec4:	data_out=16'h89f5;
17'h8ec5:	data_out=16'h89ff;
17'h8ec6:	data_out=16'h9c5;
17'h8ec7:	data_out=16'h829b;
17'h8ec8:	data_out=16'h9d5;
17'h8ec9:	data_out=16'h89e8;
17'h8eca:	data_out=16'h965;
17'h8ecb:	data_out=16'h332;
17'h8ecc:	data_out=16'h8060;
17'h8ecd:	data_out=16'ha00;
17'h8ece:	data_out=16'ha00;
17'h8ecf:	data_out=16'h88a8;
17'h8ed0:	data_out=16'h88d4;
17'h8ed1:	data_out=16'h8a00;
17'h8ed2:	data_out=16'h89e7;
17'h8ed3:	data_out=16'h9d2;
17'h8ed4:	data_out=16'h9d2;
17'h8ed5:	data_out=16'h8a00;
17'h8ed6:	data_out=16'h8a00;
17'h8ed7:	data_out=16'h89e4;
17'h8ed8:	data_out=16'h8a00;
17'h8ed9:	data_out=16'h85c3;
17'h8eda:	data_out=16'h3d1;
17'h8edb:	data_out=16'h897d;
17'h8edc:	data_out=16'h53a;
17'h8edd:	data_out=16'h9d3;
17'h8ede:	data_out=16'h9b1;
17'h8edf:	data_out=16'h9fc;
17'h8ee0:	data_out=16'h8a00;
17'h8ee1:	data_out=16'h89ea;
17'h8ee2:	data_out=16'h8a00;
17'h8ee3:	data_out=16'h173;
17'h8ee4:	data_out=16'h9d8;
17'h8ee5:	data_out=16'h8882;
17'h8ee6:	data_out=16'hf0;
17'h8ee7:	data_out=16'ha00;
17'h8ee8:	data_out=16'h80e4;
17'h8ee9:	data_out=16'h8554;
17'h8eea:	data_out=16'h81a2;
17'h8eeb:	data_out=16'h89f6;
17'h8eec:	data_out=16'h9be;
17'h8eed:	data_out=16'h235;
17'h8eee:	data_out=16'h81a0;
17'h8eef:	data_out=16'h89ff;
17'h8ef0:	data_out=16'h8171;
17'h8ef1:	data_out=16'h831f;
17'h8ef2:	data_out=16'h89d9;
17'h8ef3:	data_out=16'h873b;
17'h8ef4:	data_out=16'h81d8;
17'h8ef5:	data_out=16'h8a00;
17'h8ef6:	data_out=16'ha00;
17'h8ef7:	data_out=16'h89dd;
17'h8ef8:	data_out=16'h8431;
17'h8ef9:	data_out=16'h9ef;
17'h8efa:	data_out=16'h819e;
17'h8efb:	data_out=16'h80c9;
17'h8efc:	data_out=16'h9fc;
17'h8efd:	data_out=16'h89b7;
17'h8efe:	data_out=16'h89ed;
17'h8eff:	data_out=16'h8696;
17'h8f00:	data_out=16'h825f;
17'h8f01:	data_out=16'h853f;
17'h8f02:	data_out=16'h89fd;
17'h8f03:	data_out=16'h89fe;
17'h8f04:	data_out=16'h9ae;
17'h8f05:	data_out=16'h89fe;
17'h8f06:	data_out=16'h89fb;
17'h8f07:	data_out=16'h88d6;
17'h8f08:	data_out=16'h71;
17'h8f09:	data_out=16'h89ea;
17'h8f0a:	data_out=16'h8495;
17'h8f0b:	data_out=16'h8814;
17'h8f0c:	data_out=16'h8955;
17'h8f0d:	data_out=16'h89fe;
17'h8f0e:	data_out=16'h9b2;
17'h8f0f:	data_out=16'h899b;
17'h8f10:	data_out=16'h89f8;
17'h8f11:	data_out=16'h85ff;
17'h8f12:	data_out=16'h898c;
17'h8f13:	data_out=16'h89fd;
17'h8f14:	data_out=16'h89fe;
17'h8f15:	data_out=16'h89fc;
17'h8f16:	data_out=16'h89fd;
17'h8f17:	data_out=16'h89fe;
17'h8f18:	data_out=16'h89ce;
17'h8f19:	data_out=16'ha00;
17'h8f1a:	data_out=16'h84cc;
17'h8f1b:	data_out=16'h89fc;
17'h8f1c:	data_out=16'h8a00;
17'h8f1d:	data_out=16'h87c4;
17'h8f1e:	data_out=16'h89fc;
17'h8f1f:	data_out=16'h89fe;
17'h8f20:	data_out=16'h8950;
17'h8f21:	data_out=16'h9b1;
17'h8f22:	data_out=16'h9fb;
17'h8f23:	data_out=16'h940;
17'h8f24:	data_out=16'h93b;
17'h8f25:	data_out=16'h89e7;
17'h8f26:	data_out=16'h8619;
17'h8f27:	data_out=16'h880a;
17'h8f28:	data_out=16'h9a5;
17'h8f29:	data_out=16'h86f6;
17'h8f2a:	data_out=16'h8974;
17'h8f2b:	data_out=16'ha00;
17'h8f2c:	data_out=16'h89fe;
17'h8f2d:	data_out=16'h9f1;
17'h8f2e:	data_out=16'h89ff;
17'h8f2f:	data_out=16'h89fa;
17'h8f30:	data_out=16'h9ed;
17'h8f31:	data_out=16'h8a00;
17'h8f32:	data_out=16'h604;
17'h8f33:	data_out=16'h89fc;
17'h8f34:	data_out=16'h85b6;
17'h8f35:	data_out=16'h89f5;
17'h8f36:	data_out=16'h8972;
17'h8f37:	data_out=16'h89fe;
17'h8f38:	data_out=16'h432;
17'h8f39:	data_out=16'h89fb;
17'h8f3a:	data_out=16'h892d;
17'h8f3b:	data_out=16'h89fa;
17'h8f3c:	data_out=16'h8a00;
17'h8f3d:	data_out=16'h89d4;
17'h8f3e:	data_out=16'h9a3;
17'h8f3f:	data_out=16'h89fe;
17'h8f40:	data_out=16'h8296;
17'h8f41:	data_out=16'h89fb;
17'h8f42:	data_out=16'h8540;
17'h8f43:	data_out=16'h8a00;
17'h8f44:	data_out=16'h89eb;
17'h8f45:	data_out=16'h89fd;
17'h8f46:	data_out=16'h9ed;
17'h8f47:	data_out=16'h831e;
17'h8f48:	data_out=16'h89fb;
17'h8f49:	data_out=16'h89e6;
17'h8f4a:	data_out=16'h81c4;
17'h8f4b:	data_out=16'h818c;
17'h8f4c:	data_out=16'h4b4;
17'h8f4d:	data_out=16'h9f9;
17'h8f4e:	data_out=16'h485;
17'h8f4f:	data_out=16'h8401;
17'h8f50:	data_out=16'h89fe;
17'h8f51:	data_out=16'h8a00;
17'h8f52:	data_out=16'h8a9;
17'h8f53:	data_out=16'h89f5;
17'h8f54:	data_out=16'h8415;
17'h8f55:	data_out=16'h89ff;
17'h8f56:	data_out=16'h89fe;
17'h8f57:	data_out=16'h89d9;
17'h8f58:	data_out=16'h8159;
17'h8f59:	data_out=16'h32c;
17'h8f5a:	data_out=16'h89fd;
17'h8f5b:	data_out=16'h8935;
17'h8f5c:	data_out=16'h89ff;
17'h8f5d:	data_out=16'h873c;
17'h8f5e:	data_out=16'h89fd;
17'h8f5f:	data_out=16'h884;
17'h8f60:	data_out=16'h9a4;
17'h8f61:	data_out=16'h8630;
17'h8f62:	data_out=16'h8a00;
17'h8f63:	data_out=16'h89fc;
17'h8f64:	data_out=16'h809f;
17'h8f65:	data_out=16'h89ef;
17'h8f66:	data_out=16'h9ff;
17'h8f67:	data_out=16'ha00;
17'h8f68:	data_out=16'h9b0;
17'h8f69:	data_out=16'h6e;
17'h8f6a:	data_out=16'h9ab;
17'h8f6b:	data_out=16'h89f6;
17'h8f6c:	data_out=16'h39a;
17'h8f6d:	data_out=16'h89fc;
17'h8f6e:	data_out=16'h9ab;
17'h8f6f:	data_out=16'h89fd;
17'h8f70:	data_out=16'h9b0;
17'h8f71:	data_out=16'h899d;
17'h8f72:	data_out=16'h845d;
17'h8f73:	data_out=16'h80ba;
17'h8f74:	data_out=16'h973;
17'h8f75:	data_out=16'h8a00;
17'h8f76:	data_out=16'ha00;
17'h8f77:	data_out=16'h8966;
17'h8f78:	data_out=16'h80c3;
17'h8f79:	data_out=16'h2ed;
17'h8f7a:	data_out=16'h89fd;
17'h8f7b:	data_out=16'h9a3;
17'h8f7c:	data_out=16'h8090;
17'h8f7d:	data_out=16'h89e5;
17'h8f7e:	data_out=16'h89ef;
17'h8f7f:	data_out=16'h88bd;
17'h8f80:	data_out=16'h8325;
17'h8f81:	data_out=16'h89f9;
17'h8f82:	data_out=16'h530;
17'h8f83:	data_out=16'h89d6;
17'h8f84:	data_out=16'h89c5;
17'h8f85:	data_out=16'h89fe;
17'h8f86:	data_out=16'h8a00;
17'h8f87:	data_out=16'h85e1;
17'h8f88:	data_out=16'h850f;
17'h8f89:	data_out=16'h89c3;
17'h8f8a:	data_out=16'h854f;
17'h8f8b:	data_out=16'h87b8;
17'h8f8c:	data_out=16'h869c;
17'h8f8d:	data_out=16'h89fc;
17'h8f8e:	data_out=16'h9fd;
17'h8f8f:	data_out=16'h8253;
17'h8f90:	data_out=16'h89e4;
17'h8f91:	data_out=16'h89ef;
17'h8f92:	data_out=16'h89db;
17'h8f93:	data_out=16'h89c9;
17'h8f94:	data_out=16'h89fe;
17'h8f95:	data_out=16'h89fc;
17'h8f96:	data_out=16'h89fa;
17'h8f97:	data_out=16'h89fd;
17'h8f98:	data_out=16'h89f8;
17'h8f99:	data_out=16'ha00;
17'h8f9a:	data_out=16'h89f6;
17'h8f9b:	data_out=16'h89fa;
17'h8f9c:	data_out=16'h89fc;
17'h8f9d:	data_out=16'h89f9;
17'h8f9e:	data_out=16'h89f8;
17'h8f9f:	data_out=16'h8a00;
17'h8fa0:	data_out=16'h89ed;
17'h8fa1:	data_out=16'h9f7;
17'h8fa2:	data_out=16'ha00;
17'h8fa3:	data_out=16'h9ee;
17'h8fa4:	data_out=16'h9ef;
17'h8fa5:	data_out=16'h89c1;
17'h8fa6:	data_out=16'h9f9;
17'h8fa7:	data_out=16'h89f3;
17'h8fa8:	data_out=16'h9dc;
17'h8fa9:	data_out=16'h292;
17'h8faa:	data_out=16'h6de;
17'h8fab:	data_out=16'h9f9;
17'h8fac:	data_out=16'h89fb;
17'h8fad:	data_out=16'ha00;
17'h8fae:	data_out=16'h86c2;
17'h8faf:	data_out=16'h89f5;
17'h8fb0:	data_out=16'ha00;
17'h8fb1:	data_out=16'h8a00;
17'h8fb2:	data_out=16'h6b7;
17'h8fb3:	data_out=16'h89fe;
17'h8fb4:	data_out=16'h8949;
17'h8fb5:	data_out=16'h89f3;
17'h8fb6:	data_out=16'h8985;
17'h8fb7:	data_out=16'h8150;
17'h8fb8:	data_out=16'h8a00;
17'h8fb9:	data_out=16'h89fd;
17'h8fba:	data_out=16'h884b;
17'h8fbb:	data_out=16'h89fc;
17'h8fbc:	data_out=16'h8965;
17'h8fbd:	data_out=16'h89d2;
17'h8fbe:	data_out=16'h9db;
17'h8fbf:	data_out=16'h89fe;
17'h8fc0:	data_out=16'h89a6;
17'h8fc1:	data_out=16'h89f6;
17'h8fc2:	data_out=16'h9f3;
17'h8fc3:	data_out=16'h89fe;
17'h8fc4:	data_out=16'h89f9;
17'h8fc5:	data_out=16'h89fc;
17'h8fc6:	data_out=16'ha00;
17'h8fc7:	data_out=16'h6ff;
17'h8fc8:	data_out=16'h89fc;
17'h8fc9:	data_out=16'h89be;
17'h8fca:	data_out=16'h88d7;
17'h8fcb:	data_out=16'h8445;
17'h8fcc:	data_out=16'ha00;
17'h8fcd:	data_out=16'h9f6;
17'h8fce:	data_out=16'ha00;
17'h8fcf:	data_out=16'ha00;
17'h8fd0:	data_out=16'h89fb;
17'h8fd1:	data_out=16'h8a00;
17'h8fd2:	data_out=16'h9f6;
17'h8fd3:	data_out=16'h89fa;
17'h8fd4:	data_out=16'h89e6;
17'h8fd5:	data_out=16'h89f5;
17'h8fd6:	data_out=16'h101;
17'h8fd7:	data_out=16'h404;
17'h8fd8:	data_out=16'h8790;
17'h8fd9:	data_out=16'h8910;
17'h8fda:	data_out=16'h8a00;
17'h8fdb:	data_out=16'h89f6;
17'h8fdc:	data_out=16'h8a00;
17'h8fdd:	data_out=16'h89df;
17'h8fde:	data_out=16'h89fa;
17'h8fdf:	data_out=16'h15f;
17'h8fe0:	data_out=16'h9fa;
17'h8fe1:	data_out=16'h89e9;
17'h8fe2:	data_out=16'h89fe;
17'h8fe3:	data_out=16'h89fe;
17'h8fe4:	data_out=16'h86a4;
17'h8fe5:	data_out=16'h89f1;
17'h8fe6:	data_out=16'h9f8;
17'h8fe7:	data_out=16'ha00;
17'h8fe8:	data_out=16'h9f0;
17'h8fe9:	data_out=16'h13a;
17'h8fea:	data_out=16'h9fe;
17'h8feb:	data_out=16'h89fc;
17'h8fec:	data_out=16'h9e2;
17'h8fed:	data_out=16'h89fe;
17'h8fee:	data_out=16'h9fe;
17'h8fef:	data_out=16'h89f9;
17'h8ff0:	data_out=16'h9fd;
17'h8ff1:	data_out=16'h8668;
17'h8ff2:	data_out=16'h89b9;
17'h8ff3:	data_out=16'h89ba;
17'h8ff4:	data_out=16'ha00;
17'h8ff5:	data_out=16'h8a00;
17'h8ff6:	data_out=16'ha00;
17'h8ff7:	data_out=16'h87ad;
17'h8ff8:	data_out=16'h449;
17'h8ff9:	data_out=16'h9ee;
17'h8ffa:	data_out=16'h89fe;
17'h8ffb:	data_out=16'h9db;
17'h8ffc:	data_out=16'h89fb;
17'h8ffd:	data_out=16'h89fa;
17'h8ffe:	data_out=16'h89d7;
17'h8fff:	data_out=16'h89f8;
17'h9000:	data_out=16'h9f4;
17'h9001:	data_out=16'h89f3;
17'h9002:	data_out=16'h9ea;
17'h9003:	data_out=16'h84fa;
17'h9004:	data_out=16'h89ee;
17'h9005:	data_out=16'h8a00;
17'h9006:	data_out=16'h8a00;
17'h9007:	data_out=16'h89be;
17'h9008:	data_out=16'h2c9;
17'h9009:	data_out=16'h8850;
17'h900a:	data_out=16'h86aa;
17'h900b:	data_out=16'h87c7;
17'h900c:	data_out=16'h8115;
17'h900d:	data_out=16'h89b0;
17'h900e:	data_out=16'ha00;
17'h900f:	data_out=16'h9fb;
17'h9010:	data_out=16'h8915;
17'h9011:	data_out=16'h89ff;
17'h9012:	data_out=16'h88b3;
17'h9013:	data_out=16'h888e;
17'h9014:	data_out=16'h89e5;
17'h9015:	data_out=16'h89e8;
17'h9016:	data_out=16'h89bb;
17'h9017:	data_out=16'h89d8;
17'h9018:	data_out=16'h80c4;
17'h9019:	data_out=16'h9fc;
17'h901a:	data_out=16'h89fb;
17'h901b:	data_out=16'h89da;
17'h901c:	data_out=16'h89cd;
17'h901d:	data_out=16'h89f8;
17'h901e:	data_out=16'h894e;
17'h901f:	data_out=16'h8a00;
17'h9020:	data_out=16'h89ec;
17'h9021:	data_out=16'ha00;
17'h9022:	data_out=16'ha00;
17'h9023:	data_out=16'h9f6;
17'h9024:	data_out=16'h9f6;
17'h9025:	data_out=16'ha00;
17'h9026:	data_out=16'ha00;
17'h9027:	data_out=16'h89f0;
17'h9028:	data_out=16'h9ff;
17'h9029:	data_out=16'h9f8;
17'h902a:	data_out=16'ha00;
17'h902b:	data_out=16'h9c3;
17'h902c:	data_out=16'h89cc;
17'h902d:	data_out=16'ha00;
17'h902e:	data_out=16'h89a5;
17'h902f:	data_out=16'h89ef;
17'h9030:	data_out=16'ha00;
17'h9031:	data_out=16'h8a00;
17'h9032:	data_out=16'h3f3;
17'h9033:	data_out=16'h89fa;
17'h9034:	data_out=16'h89cf;
17'h9035:	data_out=16'h89e7;
17'h9036:	data_out=16'h155;
17'h9037:	data_out=16'h9c3;
17'h9038:	data_out=16'h8a00;
17'h9039:	data_out=16'h89f4;
17'h903a:	data_out=16'h8492;
17'h903b:	data_out=16'h89fe;
17'h903c:	data_out=16'h287;
17'h903d:	data_out=16'h888a;
17'h903e:	data_out=16'h9ff;
17'h903f:	data_out=16'h8a00;
17'h9040:	data_out=16'h88dd;
17'h9041:	data_out=16'h89de;
17'h9042:	data_out=16'ha00;
17'h9043:	data_out=16'h89e0;
17'h9044:	data_out=16'h89fb;
17'h9045:	data_out=16'h89e7;
17'h9046:	data_out=16'ha00;
17'h9047:	data_out=16'ha00;
17'h9048:	data_out=16'h89fb;
17'h9049:	data_out=16'ha00;
17'h904a:	data_out=16'h89f8;
17'h904b:	data_out=16'h83a8;
17'h904c:	data_out=16'ha00;
17'h904d:	data_out=16'ha00;
17'h904e:	data_out=16'ha00;
17'h904f:	data_out=16'ha00;
17'h9050:	data_out=16'h89d6;
17'h9051:	data_out=16'h89ea;
17'h9052:	data_out=16'h9ff;
17'h9053:	data_out=16'h89f8;
17'h9054:	data_out=16'h89b2;
17'h9055:	data_out=16'h89af;
17'h9056:	data_out=16'h9e0;
17'h9057:	data_out=16'ha00;
17'h9058:	data_out=16'h844c;
17'h9059:	data_out=16'h878;
17'h905a:	data_out=16'h89ff;
17'h905b:	data_out=16'h89f3;
17'h905c:	data_out=16'h8a00;
17'h905d:	data_out=16'ha00;
17'h905e:	data_out=16'h89f2;
17'h905f:	data_out=16'h281;
17'h9060:	data_out=16'ha00;
17'h9061:	data_out=16'h89f1;
17'h9062:	data_out=16'h89c6;
17'h9063:	data_out=16'h89fb;
17'h9064:	data_out=16'h87b2;
17'h9065:	data_out=16'h89fc;
17'h9066:	data_out=16'h9f7;
17'h9067:	data_out=16'ha00;
17'h9068:	data_out=16'ha00;
17'h9069:	data_out=16'h81e;
17'h906a:	data_out=16'ha00;
17'h906b:	data_out=16'h89f4;
17'h906c:	data_out=16'ha00;
17'h906d:	data_out=16'h89fa;
17'h906e:	data_out=16'ha00;
17'h906f:	data_out=16'h89f6;
17'h9070:	data_out=16'ha00;
17'h9071:	data_out=16'h831d;
17'h9072:	data_out=16'h8992;
17'h9073:	data_out=16'h8980;
17'h9074:	data_out=16'ha00;
17'h9075:	data_out=16'h8a00;
17'h9076:	data_out=16'ha00;
17'h9077:	data_out=16'ha00;
17'h9078:	data_out=16'h781;
17'h9079:	data_out=16'h9d9;
17'h907a:	data_out=16'h89f8;
17'h907b:	data_out=16'h9ff;
17'h907c:	data_out=16'h89fe;
17'h907d:	data_out=16'h8a00;
17'h907e:	data_out=16'h89b9;
17'h907f:	data_out=16'h8a00;
17'h9080:	data_out=16'h9fd;
17'h9081:	data_out=16'h89c3;
17'h9082:	data_out=16'h9f7;
17'h9083:	data_out=16'h413;
17'h9084:	data_out=16'h89fa;
17'h9085:	data_out=16'h8a00;
17'h9086:	data_out=16'h8a00;
17'h9087:	data_out=16'h89da;
17'h9088:	data_out=16'h829;
17'h9089:	data_out=16'h705;
17'h908a:	data_out=16'h99a;
17'h908b:	data_out=16'h89bf;
17'h908c:	data_out=16'h7ca;
17'h908d:	data_out=16'h1f2;
17'h908e:	data_out=16'ha00;
17'h908f:	data_out=16'h9fd;
17'h9090:	data_out=16'h8782;
17'h9091:	data_out=16'h89fd;
17'h9092:	data_out=16'h8757;
17'h9093:	data_out=16'h84dd;
17'h9094:	data_out=16'h89ec;
17'h9095:	data_out=16'h854a;
17'h9096:	data_out=16'h113;
17'h9097:	data_out=16'h89cc;
17'h9098:	data_out=16'h98f;
17'h9099:	data_out=16'h9f1;
17'h909a:	data_out=16'h8a00;
17'h909b:	data_out=16'h89c7;
17'h909c:	data_out=16'h89c3;
17'h909d:	data_out=16'h89f7;
17'h909e:	data_out=16'h86c0;
17'h909f:	data_out=16'h8a00;
17'h90a0:	data_out=16'h89f5;
17'h90a1:	data_out=16'ha00;
17'h90a2:	data_out=16'ha00;
17'h90a3:	data_out=16'h9ff;
17'h90a4:	data_out=16'h9ff;
17'h90a5:	data_out=16'ha00;
17'h90a6:	data_out=16'ha00;
17'h90a7:	data_out=16'h89fa;
17'h90a8:	data_out=16'ha00;
17'h90a9:	data_out=16'ha00;
17'h90aa:	data_out=16'ha00;
17'h90ab:	data_out=16'h89ea;
17'h90ac:	data_out=16'h89ba;
17'h90ad:	data_out=16'ha00;
17'h90ae:	data_out=16'h89ce;
17'h90af:	data_out=16'h89cf;
17'h90b0:	data_out=16'ha00;
17'h90b1:	data_out=16'h8a00;
17'h90b2:	data_out=16'hc1;
17'h90b3:	data_out=16'h89fc;
17'h90b4:	data_out=16'h895b;
17'h90b5:	data_out=16'h89ec;
17'h90b6:	data_out=16'h9ee;
17'h90b7:	data_out=16'h9f6;
17'h90b8:	data_out=16'h8a00;
17'h90b9:	data_out=16'h89f4;
17'h90ba:	data_out=16'ha00;
17'h90bb:	data_out=16'h8a00;
17'h90bc:	data_out=16'h8908;
17'h90bd:	data_out=16'h8118;
17'h90be:	data_out=16'ha00;
17'h90bf:	data_out=16'h8a00;
17'h90c0:	data_out=16'h376;
17'h90c1:	data_out=16'h41f;
17'h90c2:	data_out=16'ha00;
17'h90c3:	data_out=16'h89f3;
17'h90c4:	data_out=16'h8a00;
17'h90c5:	data_out=16'h842b;
17'h90c6:	data_out=16'ha00;
17'h90c7:	data_out=16'ha00;
17'h90c8:	data_out=16'h89d9;
17'h90c9:	data_out=16'ha00;
17'h90ca:	data_out=16'h89ff;
17'h90cb:	data_out=16'ha00;
17'h90cc:	data_out=16'ha00;
17'h90cd:	data_out=16'h9ff;
17'h90ce:	data_out=16'h9f8;
17'h90cf:	data_out=16'ha00;
17'h90d0:	data_out=16'h89e3;
17'h90d1:	data_out=16'h89d5;
17'h90d2:	data_out=16'ha00;
17'h90d3:	data_out=16'h89ff;
17'h90d4:	data_out=16'h8995;
17'h90d5:	data_out=16'h870d;
17'h90d6:	data_out=16'ha00;
17'h90d7:	data_out=16'ha00;
17'h90d8:	data_out=16'h168;
17'h90d9:	data_out=16'h9fe;
17'h90da:	data_out=16'h8a00;
17'h90db:	data_out=16'h89fa;
17'h90dc:	data_out=16'h8a00;
17'h90dd:	data_out=16'ha00;
17'h90de:	data_out=16'h89ac;
17'h90df:	data_out=16'h9fd;
17'h90e0:	data_out=16'ha00;
17'h90e1:	data_out=16'h89dd;
17'h90e2:	data_out=16'h89aa;
17'h90e3:	data_out=16'h89ff;
17'h90e4:	data_out=16'h88cf;
17'h90e5:	data_out=16'h8a00;
17'h90e6:	data_out=16'h9f6;
17'h90e7:	data_out=16'ha00;
17'h90e8:	data_out=16'ha00;
17'h90e9:	data_out=16'h9cb;
17'h90ea:	data_out=16'ha00;
17'h90eb:	data_out=16'h8a00;
17'h90ec:	data_out=16'ha00;
17'h90ed:	data_out=16'h89fd;
17'h90ee:	data_out=16'ha00;
17'h90ef:	data_out=16'h8a00;
17'h90f0:	data_out=16'ha00;
17'h90f1:	data_out=16'h8b2;
17'h90f2:	data_out=16'h8863;
17'h90f3:	data_out=16'h88fc;
17'h90f4:	data_out=16'ha00;
17'h90f5:	data_out=16'h8a00;
17'h90f6:	data_out=16'ha00;
17'h90f7:	data_out=16'ha00;
17'h90f8:	data_out=16'h89fb;
17'h90f9:	data_out=16'h9fa;
17'h90fa:	data_out=16'h89f4;
17'h90fb:	data_out=16'ha00;
17'h90fc:	data_out=16'h88b1;
17'h90fd:	data_out=16'h8a00;
17'h90fe:	data_out=16'h89da;
17'h90ff:	data_out=16'h8a00;
17'h9100:	data_out=16'ha00;
17'h9101:	data_out=16'h92;
17'h9102:	data_out=16'h9f7;
17'h9103:	data_out=16'ha00;
17'h9104:	data_out=16'h89aa;
17'h9105:	data_out=16'h8a00;
17'h9106:	data_out=16'h8a00;
17'h9107:	data_out=16'h89fa;
17'h9108:	data_out=16'h53a;
17'h9109:	data_out=16'h2f2;
17'h910a:	data_out=16'h9f7;
17'h910b:	data_out=16'h89fc;
17'h910c:	data_out=16'h84a8;
17'h910d:	data_out=16'h8de;
17'h910e:	data_out=16'ha00;
17'h910f:	data_out=16'h9d7;
17'h9110:	data_out=16'h1ab;
17'h9111:	data_out=16'h89fe;
17'h9112:	data_out=16'h89d4;
17'h9113:	data_out=16'h461;
17'h9114:	data_out=16'h8a00;
17'h9115:	data_out=16'h9df;
17'h9116:	data_out=16'h9c5;
17'h9117:	data_out=16'h8a00;
17'h9118:	data_out=16'h8be;
17'h9119:	data_out=16'h849a;
17'h911a:	data_out=16'h8a00;
17'h911b:	data_out=16'h89e8;
17'h911c:	data_out=16'h85aa;
17'h911d:	data_out=16'h8a00;
17'h911e:	data_out=16'hbd;
17'h911f:	data_out=16'h8a00;
17'h9120:	data_out=16'h89e2;
17'h9121:	data_out=16'ha00;
17'h9122:	data_out=16'h9fc;
17'h9123:	data_out=16'ha00;
17'h9124:	data_out=16'ha00;
17'h9125:	data_out=16'ha00;
17'h9126:	data_out=16'ha00;
17'h9127:	data_out=16'h8a00;
17'h9128:	data_out=16'ha00;
17'h9129:	data_out=16'h9fe;
17'h912a:	data_out=16'h9c5;
17'h912b:	data_out=16'h89fb;
17'h912c:	data_out=16'h96a;
17'h912d:	data_out=16'h9e1;
17'h912e:	data_out=16'h8a00;
17'h912f:	data_out=16'h89b9;
17'h9130:	data_out=16'ha00;
17'h9131:	data_out=16'h8a00;
17'h9132:	data_out=16'h59a;
17'h9133:	data_out=16'h8a00;
17'h9134:	data_out=16'h899a;
17'h9135:	data_out=16'h89a3;
17'h9136:	data_out=16'h8e2;
17'h9137:	data_out=16'h9f2;
17'h9138:	data_out=16'h8a00;
17'h9139:	data_out=16'h8a00;
17'h913a:	data_out=16'h9ae;
17'h913b:	data_out=16'h8a00;
17'h913c:	data_out=16'h922;
17'h913d:	data_out=16'h9cf;
17'h913e:	data_out=16'ha00;
17'h913f:	data_out=16'h8a00;
17'h9140:	data_out=16'h788;
17'h9141:	data_out=16'h9ef;
17'h9142:	data_out=16'ha00;
17'h9143:	data_out=16'h8a00;
17'h9144:	data_out=16'h8a00;
17'h9145:	data_out=16'h9dd;
17'h9146:	data_out=16'h9eb;
17'h9147:	data_out=16'h8d4;
17'h9148:	data_out=16'h89dc;
17'h9149:	data_out=16'ha00;
17'h914a:	data_out=16'h89ff;
17'h914b:	data_out=16'h9fc;
17'h914c:	data_out=16'ha00;
17'h914d:	data_out=16'h9fa;
17'h914e:	data_out=16'h851;
17'h914f:	data_out=16'ha00;
17'h9150:	data_out=16'h89df;
17'h9151:	data_out=16'h77e;
17'h9152:	data_out=16'ha00;
17'h9153:	data_out=16'h8a00;
17'h9154:	data_out=16'h8982;
17'h9155:	data_out=16'h987;
17'h9156:	data_out=16'ha00;
17'h9157:	data_out=16'h9da;
17'h9158:	data_out=16'h735;
17'h9159:	data_out=16'h9ff;
17'h915a:	data_out=16'h8a00;
17'h915b:	data_out=16'h8a00;
17'h915c:	data_out=16'h8a00;
17'h915d:	data_out=16'ha00;
17'h915e:	data_out=16'h8460;
17'h915f:	data_out=16'h9c1;
17'h9160:	data_out=16'ha00;
17'h9161:	data_out=16'h89d3;
17'h9162:	data_out=16'h89f6;
17'h9163:	data_out=16'h8a00;
17'h9164:	data_out=16'h89d0;
17'h9165:	data_out=16'h8a00;
17'h9166:	data_out=16'h8fd;
17'h9167:	data_out=16'ha00;
17'h9168:	data_out=16'ha00;
17'h9169:	data_out=16'h97f;
17'h916a:	data_out=16'ha00;
17'h916b:	data_out=16'h8a00;
17'h916c:	data_out=16'ha00;
17'h916d:	data_out=16'h8a00;
17'h916e:	data_out=16'ha00;
17'h916f:	data_out=16'h89e3;
17'h9170:	data_out=16'ha00;
17'h9171:	data_out=16'h23d;
17'h9172:	data_out=16'h987;
17'h9173:	data_out=16'h84;
17'h9174:	data_out=16'ha00;
17'h9175:	data_out=16'h8a00;
17'h9176:	data_out=16'h9dd;
17'h9177:	data_out=16'h9fc;
17'h9178:	data_out=16'h8a00;
17'h9179:	data_out=16'ha00;
17'h917a:	data_out=16'h8a00;
17'h917b:	data_out=16'ha00;
17'h917c:	data_out=16'h87bc;
17'h917d:	data_out=16'h8a00;
17'h917e:	data_out=16'h8a00;
17'h917f:	data_out=16'h8a00;
17'h9180:	data_out=16'h9f6;
17'h9181:	data_out=16'h91c;
17'h9182:	data_out=16'h9ac;
17'h9183:	data_out=16'h9f0;
17'h9184:	data_out=16'h89a9;
17'h9185:	data_out=16'h8a00;
17'h9186:	data_out=16'h8a00;
17'h9187:	data_out=16'h89f7;
17'h9188:	data_out=16'h323;
17'h9189:	data_out=16'h89e5;
17'h918a:	data_out=16'h9ef;
17'h918b:	data_out=16'h8a00;
17'h918c:	data_out=16'h89ff;
17'h918d:	data_out=16'h939;
17'h918e:	data_out=16'ha00;
17'h918f:	data_out=16'h935;
17'h9190:	data_out=16'h89ee;
17'h9191:	data_out=16'h8319;
17'h9192:	data_out=16'h89fa;
17'h9193:	data_out=16'h6be;
17'h9194:	data_out=16'h8a00;
17'h9195:	data_out=16'h9d9;
17'h9196:	data_out=16'h978;
17'h9197:	data_out=16'h8a00;
17'h9198:	data_out=16'h83a;
17'h9199:	data_out=16'h89e3;
17'h919a:	data_out=16'h8a00;
17'h919b:	data_out=16'h89f1;
17'h919c:	data_out=16'hd2;
17'h919d:	data_out=16'h8778;
17'h919e:	data_out=16'hd2;
17'h919f:	data_out=16'h8a00;
17'h91a0:	data_out=16'h8a00;
17'h91a1:	data_out=16'ha00;
17'h91a2:	data_out=16'h8515;
17'h91a3:	data_out=16'ha00;
17'h91a4:	data_out=16'ha00;
17'h91a5:	data_out=16'h9fc;
17'h91a6:	data_out=16'ha00;
17'h91a7:	data_out=16'h8a00;
17'h91a8:	data_out=16'ha00;
17'h91a9:	data_out=16'h9fe;
17'h91aa:	data_out=16'h83a;
17'h91ab:	data_out=16'h8a00;
17'h91ac:	data_out=16'h956;
17'h91ad:	data_out=16'h88db;
17'h91ae:	data_out=16'h8a00;
17'h91af:	data_out=16'h896b;
17'h91b0:	data_out=16'h37;
17'h91b1:	data_out=16'h89ce;
17'h91b2:	data_out=16'h8914;
17'h91b3:	data_out=16'h8a00;
17'h91b4:	data_out=16'h98f;
17'h91b5:	data_out=16'h8559;
17'h91b6:	data_out=16'h6af;
17'h91b7:	data_out=16'h999;
17'h91b8:	data_out=16'h8a00;
17'h91b9:	data_out=16'h8a00;
17'h91ba:	data_out=16'h7d8;
17'h91bb:	data_out=16'h8a00;
17'h91bc:	data_out=16'h9d0;
17'h91bd:	data_out=16'h8fa;
17'h91be:	data_out=16'ha00;
17'h91bf:	data_out=16'h8a00;
17'h91c0:	data_out=16'h628;
17'h91c1:	data_out=16'h9f5;
17'h91c2:	data_out=16'ha00;
17'h91c3:	data_out=16'h8a00;
17'h91c4:	data_out=16'h8a00;
17'h91c5:	data_out=16'h9d8;
17'h91c6:	data_out=16'h9e2;
17'h91c7:	data_out=16'h5ca;
17'h91c8:	data_out=16'h8a00;
17'h91c9:	data_out=16'ha00;
17'h91ca:	data_out=16'h89ff;
17'h91cb:	data_out=16'h966;
17'h91cc:	data_out=16'ha00;
17'h91cd:	data_out=16'h89ee;
17'h91ce:	data_out=16'h4bb;
17'h91cf:	data_out=16'ha00;
17'h91d0:	data_out=16'h8a00;
17'h91d1:	data_out=16'h92e;
17'h91d2:	data_out=16'ha00;
17'h91d3:	data_out=16'h8a00;
17'h91d4:	data_out=16'h8a00;
17'h91d5:	data_out=16'h987;
17'h91d6:	data_out=16'ha00;
17'h91d7:	data_out=16'h9df;
17'h91d8:	data_out=16'h912;
17'h91d9:	data_out=16'h9ae;
17'h91da:	data_out=16'h8a00;
17'h91db:	data_out=16'h8a00;
17'h91dc:	data_out=16'h89f3;
17'h91dd:	data_out=16'h9fe;
17'h91de:	data_out=16'h247;
17'h91df:	data_out=16'h8da;
17'h91e0:	data_out=16'h9ec;
17'h91e1:	data_out=16'h89da;
17'h91e2:	data_out=16'h8a00;
17'h91e3:	data_out=16'h8a00;
17'h91e4:	data_out=16'h8a00;
17'h91e5:	data_out=16'h89fe;
17'h91e6:	data_out=16'h89fc;
17'h91e7:	data_out=16'ha00;
17'h91e8:	data_out=16'ha00;
17'h91e9:	data_out=16'h966;
17'h91ea:	data_out=16'ha00;
17'h91eb:	data_out=16'h89ec;
17'h91ec:	data_out=16'h9f5;
17'h91ed:	data_out=16'h8a00;
17'h91ee:	data_out=16'ha00;
17'h91ef:	data_out=16'h89e5;
17'h91f0:	data_out=16'ha00;
17'h91f1:	data_out=16'h8033;
17'h91f2:	data_out=16'h973;
17'h91f3:	data_out=16'h85a1;
17'h91f4:	data_out=16'h823b;
17'h91f5:	data_out=16'h8a00;
17'h91f6:	data_out=16'h89ff;
17'h91f7:	data_out=16'h905;
17'h91f8:	data_out=16'h8a00;
17'h91f9:	data_out=16'ha00;
17'h91fa:	data_out=16'h8a00;
17'h91fb:	data_out=16'ha00;
17'h91fc:	data_out=16'h82d4;
17'h91fd:	data_out=16'h8a00;
17'h91fe:	data_out=16'h8a00;
17'h91ff:	data_out=16'h8a00;
17'h9200:	data_out=16'h9f3;
17'h9201:	data_out=16'h378;
17'h9202:	data_out=16'h986;
17'h9203:	data_out=16'h86ca;
17'h9204:	data_out=16'h89af;
17'h9205:	data_out=16'h89ed;
17'h9206:	data_out=16'h8a00;
17'h9207:	data_out=16'h8470;
17'h9208:	data_out=16'h350;
17'h9209:	data_out=16'h89e6;
17'h920a:	data_out=16'h665;
17'h920b:	data_out=16'h8a00;
17'h920c:	data_out=16'h8294;
17'h920d:	data_out=16'h94b;
17'h920e:	data_out=16'h9fe;
17'h920f:	data_out=16'h8a9;
17'h9210:	data_out=16'h8a00;
17'h9211:	data_out=16'h2fa;
17'h9212:	data_out=16'h89fb;
17'h9213:	data_out=16'h84c1;
17'h9214:	data_out=16'h8a00;
17'h9215:	data_out=16'h823;
17'h9216:	data_out=16'h92d;
17'h9217:	data_out=16'h8a00;
17'h9218:	data_out=16'h7cf;
17'h9219:	data_out=16'h8a00;
17'h921a:	data_out=16'h8a00;
17'h921b:	data_out=16'h89f9;
17'h921c:	data_out=16'h89d6;
17'h921d:	data_out=16'h8720;
17'h921e:	data_out=16'h8a00;
17'h921f:	data_out=16'h8a00;
17'h9220:	data_out=16'h89ee;
17'h9221:	data_out=16'h9fb;
17'h9222:	data_out=16'h8a00;
17'h9223:	data_out=16'ha00;
17'h9224:	data_out=16'ha00;
17'h9225:	data_out=16'h80aa;
17'h9226:	data_out=16'h9fd;
17'h9227:	data_out=16'h8a00;
17'h9228:	data_out=16'h9f6;
17'h9229:	data_out=16'h9f4;
17'h922a:	data_out=16'h6d9;
17'h922b:	data_out=16'h8a00;
17'h922c:	data_out=16'h91a;
17'h922d:	data_out=16'h8a00;
17'h922e:	data_out=16'h89ff;
17'h922f:	data_out=16'h88cd;
17'h9230:	data_out=16'h897e;
17'h9231:	data_out=16'h52e;
17'h9232:	data_out=16'h8a00;
17'h9233:	data_out=16'h8a00;
17'h9234:	data_out=16'h9e6;
17'h9235:	data_out=16'h89bc;
17'h9236:	data_out=16'h65c;
17'h9237:	data_out=16'h8536;
17'h9238:	data_out=16'h89b6;
17'h9239:	data_out=16'h8a00;
17'h923a:	data_out=16'h89ef;
17'h923b:	data_out=16'h8a00;
17'h923c:	data_out=16'h176;
17'h923d:	data_out=16'h898d;
17'h923e:	data_out=16'h9f5;
17'h923f:	data_out=16'h89eb;
17'h9240:	data_out=16'h89e5;
17'h9241:	data_out=16'h9fa;
17'h9242:	data_out=16'h9ff;
17'h9243:	data_out=16'h8a00;
17'h9244:	data_out=16'h8a00;
17'h9245:	data_out=16'h9af;
17'h9246:	data_out=16'h995;
17'h9247:	data_out=16'h83de;
17'h9248:	data_out=16'h89da;
17'h9249:	data_out=16'h3f;
17'h924a:	data_out=16'h8a00;
17'h924b:	data_out=16'h962;
17'h924c:	data_out=16'h9fb;
17'h924d:	data_out=16'h8a00;
17'h924e:	data_out=16'h4df;
17'h924f:	data_out=16'h9dd;
17'h9250:	data_out=16'h89f4;
17'h9251:	data_out=16'h8880;
17'h9252:	data_out=16'ha00;
17'h9253:	data_out=16'h8a00;
17'h9254:	data_out=16'h89e2;
17'h9255:	data_out=16'h89db;
17'h9256:	data_out=16'h9ff;
17'h9257:	data_out=16'h821d;
17'h9258:	data_out=16'h8fb;
17'h9259:	data_out=16'h838c;
17'h925a:	data_out=16'h8a00;
17'h925b:	data_out=16'h8a00;
17'h925c:	data_out=16'h9f2;
17'h925d:	data_out=16'h9f2;
17'h925e:	data_out=16'h8263;
17'h925f:	data_out=16'h3d1;
17'h9260:	data_out=16'h81d;
17'h9261:	data_out=16'h8a00;
17'h9262:	data_out=16'h8a00;
17'h9263:	data_out=16'h8a00;
17'h9264:	data_out=16'h89e7;
17'h9265:	data_out=16'h89e7;
17'h9266:	data_out=16'h8a00;
17'h9267:	data_out=16'h56;
17'h9268:	data_out=16'h9f9;
17'h9269:	data_out=16'h959;
17'h926a:	data_out=16'h9fe;
17'h926b:	data_out=16'h89a7;
17'h926c:	data_out=16'h9f7;
17'h926d:	data_out=16'h8a00;
17'h926e:	data_out=16'h9fe;
17'h926f:	data_out=16'h89e8;
17'h9270:	data_out=16'h9fe;
17'h9271:	data_out=16'h82f9;
17'h9272:	data_out=16'h868c;
17'h9273:	data_out=16'h884a;
17'h9274:	data_out=16'h8971;
17'h9275:	data_out=16'h81a8;
17'h9276:	data_out=16'h8a00;
17'h9277:	data_out=16'h83a0;
17'h9278:	data_out=16'h8a00;
17'h9279:	data_out=16'ha00;
17'h927a:	data_out=16'h8a00;
17'h927b:	data_out=16'h9f5;
17'h927c:	data_out=16'h8269;
17'h927d:	data_out=16'h8a00;
17'h927e:	data_out=16'h8a00;
17'h927f:	data_out=16'h8a00;
17'h9280:	data_out=16'ha00;
17'h9281:	data_out=16'h9f8;
17'h9282:	data_out=16'h8a00;
17'h9283:	data_out=16'h897b;
17'h9284:	data_out=16'h89ea;
17'h9285:	data_out=16'h89c3;
17'h9286:	data_out=16'h89f9;
17'h9287:	data_out=16'h6b9;
17'h9288:	data_out=16'h817;
17'h9289:	data_out=16'h8a00;
17'h928a:	data_out=16'h8c3;
17'h928b:	data_out=16'h8a00;
17'h928c:	data_out=16'h983;
17'h928d:	data_out=16'h6c5;
17'h928e:	data_out=16'h81ec;
17'h928f:	data_out=16'h8a00;
17'h9290:	data_out=16'h8a00;
17'h9291:	data_out=16'h2ed;
17'h9292:	data_out=16'h8a00;
17'h9293:	data_out=16'h89c0;
17'h9294:	data_out=16'h8a00;
17'h9295:	data_out=16'h89ec;
17'h9296:	data_out=16'h716;
17'h9297:	data_out=16'h89b8;
17'h9298:	data_out=16'h8a00;
17'h9299:	data_out=16'h8a00;
17'h929a:	data_out=16'h8a00;
17'h929b:	data_out=16'h8996;
17'h929c:	data_out=16'h89ad;
17'h929d:	data_out=16'h9ff;
17'h929e:	data_out=16'h8a00;
17'h929f:	data_out=16'h8a00;
17'h92a0:	data_out=16'h89ba;
17'h92a1:	data_out=16'h82b8;
17'h92a2:	data_out=16'h8a00;
17'h92a3:	data_out=16'h85d2;
17'h92a4:	data_out=16'h85a6;
17'h92a5:	data_out=16'h8a00;
17'h92a6:	data_out=16'h89c7;
17'h92a7:	data_out=16'h89f8;
17'h92a8:	data_out=16'h84be;
17'h92a9:	data_out=16'h8447;
17'h92aa:	data_out=16'h89fa;
17'h92ab:	data_out=16'h89ff;
17'h92ac:	data_out=16'h4c6;
17'h92ad:	data_out=16'h8a00;
17'h92ae:	data_out=16'h8a00;
17'h92af:	data_out=16'h673;
17'h92b0:	data_out=16'h8962;
17'h92b1:	data_out=16'h9fc;
17'h92b2:	data_out=16'h8a00;
17'h92b3:	data_out=16'h8a00;
17'h92b4:	data_out=16'ha00;
17'h92b5:	data_out=16'h8a00;
17'h92b6:	data_out=16'h49c;
17'h92b7:	data_out=16'h8a00;
17'h92b8:	data_out=16'ha00;
17'h92b9:	data_out=16'h8a00;
17'h92ba:	data_out=16'h8a00;
17'h92bb:	data_out=16'h869c;
17'h92bc:	data_out=16'h8079;
17'h92bd:	data_out=16'h8a00;
17'h92be:	data_out=16'h84c7;
17'h92bf:	data_out=16'h89c2;
17'h92c0:	data_out=16'h8a00;
17'h92c1:	data_out=16'h9fe;
17'h92c2:	data_out=16'ha00;
17'h92c3:	data_out=16'h8a00;
17'h92c4:	data_out=16'h89cb;
17'h92c5:	data_out=16'h89ea;
17'h92c6:	data_out=16'h592;
17'h92c7:	data_out=16'h8a00;
17'h92c8:	data_out=16'h8773;
17'h92c9:	data_out=16'h8a00;
17'h92ca:	data_out=16'h8234;
17'h92cb:	data_out=16'h9fd;
17'h92cc:	data_out=16'h609;
17'h92cd:	data_out=16'h8a00;
17'h92ce:	data_out=16'h898b;
17'h92cf:	data_out=16'h8a00;
17'h92d0:	data_out=16'h89e2;
17'h92d1:	data_out=16'h8a00;
17'h92d2:	data_out=16'h718;
17'h92d3:	data_out=16'h88f4;
17'h92d4:	data_out=16'h897e;
17'h92d5:	data_out=16'h8a00;
17'h92d6:	data_out=16'h9de;
17'h92d7:	data_out=16'h8a00;
17'h92d8:	data_out=16'h8c4;
17'h92d9:	data_out=16'h8a00;
17'h92da:	data_out=16'h9e7;
17'h92db:	data_out=16'h8a00;
17'h92dc:	data_out=16'ha00;
17'h92dd:	data_out=16'h9ec;
17'h92de:	data_out=16'h77d;
17'h92df:	data_out=16'h89fb;
17'h92e0:	data_out=16'h8a00;
17'h92e1:	data_out=16'h8a00;
17'h92e2:	data_out=16'h89a7;
17'h92e3:	data_out=16'h8a00;
17'h92e4:	data_out=16'h1f4;
17'h92e5:	data_out=16'h8983;
17'h92e6:	data_out=16'h8a00;
17'h92e7:	data_out=16'h8a00;
17'h92e8:	data_out=16'h83a1;
17'h92e9:	data_out=16'h5c3;
17'h92ea:	data_out=16'h819b;
17'h92eb:	data_out=16'h89bf;
17'h92ec:	data_out=16'h9fe;
17'h92ed:	data_out=16'h8a00;
17'h92ee:	data_out=16'h8198;
17'h92ef:	data_out=16'h89ce;
17'h92f0:	data_out=16'h81b7;
17'h92f1:	data_out=16'h8a00;
17'h92f2:	data_out=16'h89cc;
17'h92f3:	data_out=16'h89db;
17'h92f4:	data_out=16'h88bd;
17'h92f5:	data_out=16'h9ff;
17'h92f6:	data_out=16'h8a00;
17'h92f7:	data_out=16'h8a00;
17'h92f8:	data_out=16'h8a00;
17'h92f9:	data_out=16'h9a8;
17'h92fa:	data_out=16'h89f7;
17'h92fb:	data_out=16'h84c2;
17'h92fc:	data_out=16'h8a00;
17'h92fd:	data_out=16'h8a00;
17'h92fe:	data_out=16'h8a00;
17'h92ff:	data_out=16'h89ed;
17'h9300:	data_out=16'ha00;
17'h9301:	data_out=16'ha00;
17'h9302:	data_out=16'h8a00;
17'h9303:	data_out=16'h4d0;
17'h9304:	data_out=16'h8a00;
17'h9305:	data_out=16'h9f3;
17'h9306:	data_out=16'h8963;
17'h9307:	data_out=16'h8a00;
17'h9308:	data_out=16'h8421;
17'h9309:	data_out=16'h8a00;
17'h930a:	data_out=16'h2ae;
17'h930b:	data_out=16'h8a00;
17'h930c:	data_out=16'h12c;
17'h930d:	data_out=16'h943;
17'h930e:	data_out=16'h8a00;
17'h930f:	data_out=16'h8a00;
17'h9310:	data_out=16'h8a00;
17'h9311:	data_out=16'h8354;
17'h9312:	data_out=16'h89f2;
17'h9313:	data_out=16'h67b;
17'h9314:	data_out=16'h89c2;
17'h9315:	data_out=16'h867a;
17'h9316:	data_out=16'h9ba;
17'h9317:	data_out=16'h946;
17'h9318:	data_out=16'h8a00;
17'h9319:	data_out=16'h8a00;
17'h931a:	data_out=16'h89fe;
17'h931b:	data_out=16'h83eb;
17'h931c:	data_out=16'h9f5;
17'h931d:	data_out=16'ha00;
17'h931e:	data_out=16'h89fb;
17'h931f:	data_out=16'h8a00;
17'h9320:	data_out=16'h28;
17'h9321:	data_out=16'h8a00;
17'h9322:	data_out=16'h8a00;
17'h9323:	data_out=16'h8a00;
17'h9324:	data_out=16'h8a00;
17'h9325:	data_out=16'h8a00;
17'h9326:	data_out=16'h8a00;
17'h9327:	data_out=16'h86df;
17'h9328:	data_out=16'h8a00;
17'h9329:	data_out=16'h89f3;
17'h932a:	data_out=16'h8a00;
17'h932b:	data_out=16'h8a00;
17'h932c:	data_out=16'h99f;
17'h932d:	data_out=16'h89fd;
17'h932e:	data_out=16'h8a00;
17'h932f:	data_out=16'h9ff;
17'h9330:	data_out=16'h89fc;
17'h9331:	data_out=16'h9fc;
17'h9332:	data_out=16'h8a00;
17'h9333:	data_out=16'h89c8;
17'h9334:	data_out=16'ha00;
17'h9335:	data_out=16'h8a00;
17'h9336:	data_out=16'h873e;
17'h9337:	data_out=16'h8a00;
17'h9338:	data_out=16'ha00;
17'h9339:	data_out=16'h89d6;
17'h933a:	data_out=16'h8a00;
17'h933b:	data_out=16'h8a00;
17'h933c:	data_out=16'h950;
17'h933d:	data_out=16'h8a00;
17'h933e:	data_out=16'h8a00;
17'h933f:	data_out=16'h9f4;
17'h9340:	data_out=16'h8a00;
17'h9341:	data_out=16'ha00;
17'h9342:	data_out=16'h9c1;
17'h9343:	data_out=16'h8a00;
17'h9344:	data_out=16'h635;
17'h9345:	data_out=16'h8461;
17'h9346:	data_out=16'h89bd;
17'h9347:	data_out=16'h8a00;
17'h9348:	data_out=16'h84ee;
17'h9349:	data_out=16'h8a00;
17'h934a:	data_out=16'h805d;
17'h934b:	data_out=16'h9f6;
17'h934c:	data_out=16'h8a00;
17'h934d:	data_out=16'h8a00;
17'h934e:	data_out=16'h8a00;
17'h934f:	data_out=16'h8a00;
17'h9350:	data_out=16'h2e9;
17'h9351:	data_out=16'h89fc;
17'h9352:	data_out=16'h8a00;
17'h9353:	data_out=16'ha00;
17'h9354:	data_out=16'h7ff;
17'h9355:	data_out=16'h89ff;
17'h9356:	data_out=16'h8a00;
17'h9357:	data_out=16'h8a00;
17'h9358:	data_out=16'h9d9;
17'h9359:	data_out=16'h8a00;
17'h935a:	data_out=16'ha00;
17'h935b:	data_out=16'h8a00;
17'h935c:	data_out=16'ha00;
17'h935d:	data_out=16'h851;
17'h935e:	data_out=16'ha00;
17'h935f:	data_out=16'h89fe;
17'h9360:	data_out=16'h8a00;
17'h9361:	data_out=16'h8a00;
17'h9362:	data_out=16'h85af;
17'h9363:	data_out=16'h89a2;
17'h9364:	data_out=16'ha00;
17'h9365:	data_out=16'h846e;
17'h9366:	data_out=16'h8a00;
17'h9367:	data_out=16'h8a00;
17'h9368:	data_out=16'h8a00;
17'h9369:	data_out=16'h89e2;
17'h936a:	data_out=16'h8a00;
17'h936b:	data_out=16'h898c;
17'h936c:	data_out=16'ha00;
17'h936d:	data_out=16'h89a9;
17'h936e:	data_out=16'h8a00;
17'h936f:	data_out=16'h89db;
17'h9370:	data_out=16'h8a00;
17'h9371:	data_out=16'h8a00;
17'h9372:	data_out=16'h89eb;
17'h9373:	data_out=16'h89c8;
17'h9374:	data_out=16'h89bb;
17'h9375:	data_out=16'ha00;
17'h9376:	data_out=16'h8a00;
17'h9377:	data_out=16'h8a00;
17'h9378:	data_out=16'h8a00;
17'h9379:	data_out=16'h8735;
17'h937a:	data_out=16'h89aa;
17'h937b:	data_out=16'h8a00;
17'h937c:	data_out=16'h8a00;
17'h937d:	data_out=16'h8a00;
17'h937e:	data_out=16'h8a00;
17'h937f:	data_out=16'h878f;
17'h9380:	data_out=16'ha00;
17'h9381:	data_out=16'h9f5;
17'h9382:	data_out=16'h8a00;
17'h9383:	data_out=16'h964;
17'h9384:	data_out=16'h8a00;
17'h9385:	data_out=16'h143;
17'h9386:	data_out=16'h4b3;
17'h9387:	data_out=16'h8a00;
17'h9388:	data_out=16'h9e3;
17'h9389:	data_out=16'h8a00;
17'h938a:	data_out=16'h8a00;
17'h938b:	data_out=16'h89d2;
17'h938c:	data_out=16'h89de;
17'h938d:	data_out=16'h9ed;
17'h938e:	data_out=16'h8a00;
17'h938f:	data_out=16'h89ff;
17'h9390:	data_out=16'h8a00;
17'h9391:	data_out=16'h89e0;
17'h9392:	data_out=16'ha00;
17'h9393:	data_out=16'h9cc;
17'h9394:	data_out=16'h9ff;
17'h9395:	data_out=16'h84d9;
17'h9396:	data_out=16'h9db;
17'h9397:	data_out=16'ha00;
17'h9398:	data_out=16'h8a00;
17'h9399:	data_out=16'h8a00;
17'h939a:	data_out=16'h8a00;
17'h939b:	data_out=16'h622;
17'h939c:	data_out=16'h9f6;
17'h939d:	data_out=16'ha00;
17'h939e:	data_out=16'h784;
17'h939f:	data_out=16'h8993;
17'h93a0:	data_out=16'h9ff;
17'h93a1:	data_out=16'h8a00;
17'h93a2:	data_out=16'h8a00;
17'h93a3:	data_out=16'h8a00;
17'h93a4:	data_out=16'h8a00;
17'h93a5:	data_out=16'h8a00;
17'h93a6:	data_out=16'h8a00;
17'h93a7:	data_out=16'h8141;
17'h93a8:	data_out=16'h8a00;
17'h93a9:	data_out=16'h8a00;
17'h93aa:	data_out=16'h89ff;
17'h93ab:	data_out=16'h72f;
17'h93ac:	data_out=16'h9df;
17'h93ad:	data_out=16'h89f8;
17'h93ae:	data_out=16'h898e;
17'h93af:	data_out=16'ha00;
17'h93b0:	data_out=16'h8a00;
17'h93b1:	data_out=16'h529;
17'h93b2:	data_out=16'h8a00;
17'h93b3:	data_out=16'ha00;
17'h93b4:	data_out=16'ha00;
17'h93b5:	data_out=16'h8a00;
17'h93b6:	data_out=16'h84c;
17'h93b7:	data_out=16'h8a00;
17'h93b8:	data_out=16'ha00;
17'h93b9:	data_out=16'ha00;
17'h93ba:	data_out=16'h8a00;
17'h93bb:	data_out=16'h8a00;
17'h93bc:	data_out=16'h8096;
17'h93bd:	data_out=16'h8a00;
17'h93be:	data_out=16'h8a00;
17'h93bf:	data_out=16'h11a;
17'h93c0:	data_out=16'h8a00;
17'h93c1:	data_out=16'ha00;
17'h93c2:	data_out=16'h2fa;
17'h93c3:	data_out=16'h8a00;
17'h93c4:	data_out=16'h35f;
17'h93c5:	data_out=16'h81fe;
17'h93c6:	data_out=16'h8a00;
17'h93c7:	data_out=16'h8a00;
17'h93c8:	data_out=16'ha00;
17'h93c9:	data_out=16'h8a00;
17'h93ca:	data_out=16'h9f5;
17'h93cb:	data_out=16'h95d;
17'h93cc:	data_out=16'h8a00;
17'h93cd:	data_out=16'h8a00;
17'h93ce:	data_out=16'h467;
17'h93cf:	data_out=16'h8a00;
17'h93d0:	data_out=16'h907;
17'h93d1:	data_out=16'h26f;
17'h93d2:	data_out=16'h8a00;
17'h93d3:	data_out=16'h9ff;
17'h93d4:	data_out=16'ha00;
17'h93d5:	data_out=16'h8a00;
17'h93d6:	data_out=16'h8a00;
17'h93d7:	data_out=16'h8a00;
17'h93d8:	data_out=16'h9d6;
17'h93d9:	data_out=16'h8a00;
17'h93da:	data_out=16'ha00;
17'h93db:	data_out=16'h8a00;
17'h93dc:	data_out=16'ha00;
17'h93dd:	data_out=16'h9e8;
17'h93de:	data_out=16'ha00;
17'h93df:	data_out=16'h9b2;
17'h93e0:	data_out=16'h8a00;
17'h93e1:	data_out=16'h8a00;
17'h93e2:	data_out=16'ha00;
17'h93e3:	data_out=16'ha00;
17'h93e4:	data_out=16'ha00;
17'h93e5:	data_out=16'h89ff;
17'h93e6:	data_out=16'h8a00;
17'h93e7:	data_out=16'h8a00;
17'h93e8:	data_out=16'h8a00;
17'h93e9:	data_out=16'h89f7;
17'h93ea:	data_out=16'h8a00;
17'h93eb:	data_out=16'h89bf;
17'h93ec:	data_out=16'ha00;
17'h93ed:	data_out=16'ha00;
17'h93ee:	data_out=16'h8a00;
17'h93ef:	data_out=16'h8a00;
17'h93f0:	data_out=16'h8a00;
17'h93f1:	data_out=16'h21d;
17'h93f2:	data_out=16'h8a00;
17'h93f3:	data_out=16'h8a00;
17'h93f4:	data_out=16'h8a00;
17'h93f5:	data_out=16'h97a;
17'h93f6:	data_out=16'h8a00;
17'h93f7:	data_out=16'h8a00;
17'h93f8:	data_out=16'h8a00;
17'h93f9:	data_out=16'h85a3;
17'h93fa:	data_out=16'ha00;
17'h93fb:	data_out=16'h8a00;
17'h93fc:	data_out=16'h89f6;
17'h93fd:	data_out=16'h89b8;
17'h93fe:	data_out=16'h89b7;
17'h93ff:	data_out=16'h871d;
17'h9400:	data_out=16'h9cd;
17'h9401:	data_out=16'h9ec;
17'h9402:	data_out=16'h8a00;
17'h9403:	data_out=16'h86f;
17'h9404:	data_out=16'h8a00;
17'h9405:	data_out=16'h8a00;
17'h9406:	data_out=16'ha00;
17'h9407:	data_out=16'h8a00;
17'h9408:	data_out=16'h9c4;
17'h9409:	data_out=16'h89e1;
17'h940a:	data_out=16'h8a00;
17'h940b:	data_out=16'ha00;
17'h940c:	data_out=16'h89db;
17'h940d:	data_out=16'h6ce;
17'h940e:	data_out=16'h8a00;
17'h940f:	data_out=16'h89f9;
17'h9410:	data_out=16'h8a00;
17'h9411:	data_out=16'h8502;
17'h9412:	data_out=16'ha00;
17'h9413:	data_out=16'h819;
17'h9414:	data_out=16'h9ed;
17'h9415:	data_out=16'h8a00;
17'h9416:	data_out=16'h662;
17'h9417:	data_out=16'ha00;
17'h9418:	data_out=16'h89fd;
17'h9419:	data_out=16'h8a00;
17'h941a:	data_out=16'h8a00;
17'h941b:	data_out=16'h7de;
17'h941c:	data_out=16'h986;
17'h941d:	data_out=16'ha00;
17'h941e:	data_out=16'h985;
17'h941f:	data_out=16'h812f;
17'h9420:	data_out=16'h9a3;
17'h9421:	data_out=16'h8a00;
17'h9422:	data_out=16'h8a00;
17'h9423:	data_out=16'h8a00;
17'h9424:	data_out=16'h8a00;
17'h9425:	data_out=16'h8a00;
17'h9426:	data_out=16'h8a00;
17'h9427:	data_out=16'h4b3;
17'h9428:	data_out=16'h8a00;
17'h9429:	data_out=16'h8a00;
17'h942a:	data_out=16'h844b;
17'h942b:	data_out=16'ha00;
17'h942c:	data_out=16'h630;
17'h942d:	data_out=16'h9e9;
17'h942e:	data_out=16'h9f0;
17'h942f:	data_out=16'ha00;
17'h9430:	data_out=16'h8a00;
17'h9431:	data_out=16'h8a00;
17'h9432:	data_out=16'h8a00;
17'h9433:	data_out=16'ha00;
17'h9434:	data_out=16'ha00;
17'h9435:	data_out=16'h8a00;
17'h9436:	data_out=16'h998;
17'h9437:	data_out=16'h8a00;
17'h9438:	data_out=16'ha00;
17'h9439:	data_out=16'ha00;
17'h943a:	data_out=16'h8a00;
17'h943b:	data_out=16'h8a00;
17'h943c:	data_out=16'h8a00;
17'h943d:	data_out=16'h8a00;
17'h943e:	data_out=16'h8a00;
17'h943f:	data_out=16'h8a00;
17'h9440:	data_out=16'h8a00;
17'h9441:	data_out=16'h9ec;
17'h9442:	data_out=16'h8a00;
17'h9443:	data_out=16'h8a00;
17'h9444:	data_out=16'h8787;
17'h9445:	data_out=16'h8a00;
17'h9446:	data_out=16'h8a00;
17'h9447:	data_out=16'h89ab;
17'h9448:	data_out=16'h9ff;
17'h9449:	data_out=16'h8a00;
17'h944a:	data_out=16'h9ef;
17'h944b:	data_out=16'h857;
17'h944c:	data_out=16'h8a00;
17'h944d:	data_out=16'h8a00;
17'h944e:	data_out=16'h8ba;
17'h944f:	data_out=16'h8a00;
17'h9450:	data_out=16'h89ed;
17'h9451:	data_out=16'h145;
17'h9452:	data_out=16'h8a00;
17'h9453:	data_out=16'h9fd;
17'h9454:	data_out=16'h9ff;
17'h9455:	data_out=16'h8a00;
17'h9456:	data_out=16'h8a00;
17'h9457:	data_out=16'h8a00;
17'h9458:	data_out=16'h141;
17'h9459:	data_out=16'h8a00;
17'h945a:	data_out=16'ha00;
17'h945b:	data_out=16'h8a00;
17'h945c:	data_out=16'h99c;
17'h945d:	data_out=16'h567;
17'h945e:	data_out=16'ha00;
17'h945f:	data_out=16'h9fd;
17'h9460:	data_out=16'h8a00;
17'h9461:	data_out=16'h8a00;
17'h9462:	data_out=16'h9db;
17'h9463:	data_out=16'ha00;
17'h9464:	data_out=16'h9ff;
17'h9465:	data_out=16'h89f1;
17'h9466:	data_out=16'h89ff;
17'h9467:	data_out=16'h8a00;
17'h9468:	data_out=16'h8a00;
17'h9469:	data_out=16'h89f3;
17'h946a:	data_out=16'h8a00;
17'h946b:	data_out=16'h8a00;
17'h946c:	data_out=16'h9ec;
17'h946d:	data_out=16'ha00;
17'h946e:	data_out=16'h8a00;
17'h946f:	data_out=16'h8a00;
17'h9470:	data_out=16'h8a00;
17'h9471:	data_out=16'h95f;
17'h9472:	data_out=16'h8a00;
17'h9473:	data_out=16'h8a00;
17'h9474:	data_out=16'h8a00;
17'h9475:	data_out=16'h8a00;
17'h9476:	data_out=16'h89cb;
17'h9477:	data_out=16'h8a00;
17'h9478:	data_out=16'h8a00;
17'h9479:	data_out=16'h99e;
17'h947a:	data_out=16'ha00;
17'h947b:	data_out=16'h8a00;
17'h947c:	data_out=16'h32c;
17'h947d:	data_out=16'h898b;
17'h947e:	data_out=16'ha00;
17'h947f:	data_out=16'h8a00;
17'h9480:	data_out=16'h8915;
17'h9481:	data_out=16'h9e2;
17'h9482:	data_out=16'h8a00;
17'h9483:	data_out=16'h8506;
17'h9484:	data_out=16'h8a00;
17'h9485:	data_out=16'h8a00;
17'h9486:	data_out=16'ha00;
17'h9487:	data_out=16'h8a00;
17'h9488:	data_out=16'h80f5;
17'h9489:	data_out=16'h8970;
17'h948a:	data_out=16'h89db;
17'h948b:	data_out=16'ha00;
17'h948c:	data_out=16'h89e2;
17'h948d:	data_out=16'h8a00;
17'h948e:	data_out=16'h89fd;
17'h948f:	data_out=16'h89f4;
17'h9490:	data_out=16'h8957;
17'h9491:	data_out=16'ha00;
17'h9492:	data_out=16'h99c;
17'h9493:	data_out=16'h1f7;
17'h9494:	data_out=16'h9f1;
17'h9495:	data_out=16'h8a00;
17'h9496:	data_out=16'h8a00;
17'h9497:	data_out=16'h9f8;
17'h9498:	data_out=16'h8a00;
17'h9499:	data_out=16'h89fe;
17'h949a:	data_out=16'h8a00;
17'h949b:	data_out=16'h6f7;
17'h949c:	data_out=16'h8909;
17'h949d:	data_out=16'ha00;
17'h949e:	data_out=16'h9a1;
17'h949f:	data_out=16'h9eb;
17'h94a0:	data_out=16'h81b5;
17'h94a1:	data_out=16'h89fd;
17'h94a2:	data_out=16'h899e;
17'h94a3:	data_out=16'h8a00;
17'h94a4:	data_out=16'h8a00;
17'h94a5:	data_out=16'h8a00;
17'h94a6:	data_out=16'h8a00;
17'h94a7:	data_out=16'h9dc;
17'h94a8:	data_out=16'h89fc;
17'h94a9:	data_out=16'h8a00;
17'h94aa:	data_out=16'h838e;
17'h94ab:	data_out=16'ha00;
17'h94ac:	data_out=16'h8a00;
17'h94ad:	data_out=16'ha00;
17'h94ae:	data_out=16'h9dc;
17'h94af:	data_out=16'h9e8;
17'h94b0:	data_out=16'h8a00;
17'h94b1:	data_out=16'h45a;
17'h94b2:	data_out=16'h8a00;
17'h94b3:	data_out=16'ha00;
17'h94b4:	data_out=16'ha00;
17'h94b5:	data_out=16'h8a00;
17'h94b6:	data_out=16'h816c;
17'h94b7:	data_out=16'h8a00;
17'h94b8:	data_out=16'ha00;
17'h94b9:	data_out=16'ha00;
17'h94ba:	data_out=16'h89d5;
17'h94bb:	data_out=16'h8a00;
17'h94bc:	data_out=16'h8a00;
17'h94bd:	data_out=16'h89ff;
17'h94be:	data_out=16'h89fc;
17'h94bf:	data_out=16'h8a00;
17'h94c0:	data_out=16'h8a00;
17'h94c1:	data_out=16'h89b4;
17'h94c2:	data_out=16'h8a00;
17'h94c3:	data_out=16'h8a00;
17'h94c4:	data_out=16'h86b6;
17'h94c5:	data_out=16'h8a00;
17'h94c6:	data_out=16'h8065;
17'h94c7:	data_out=16'h294;
17'h94c8:	data_out=16'h9ee;
17'h94c9:	data_out=16'h8a00;
17'h94ca:	data_out=16'h9bb;
17'h94cb:	data_out=16'h8dc;
17'h94cc:	data_out=16'h8a00;
17'h94cd:	data_out=16'h8984;
17'h94ce:	data_out=16'h865;
17'h94cf:	data_out=16'h89f9;
17'h94d0:	data_out=16'h89d9;
17'h94d1:	data_out=16'h8a00;
17'h94d2:	data_out=16'h8a00;
17'h94d3:	data_out=16'h9cb;
17'h94d4:	data_out=16'h9ce;
17'h94d5:	data_out=16'h8a00;
17'h94d6:	data_out=16'h8a00;
17'h94d7:	data_out=16'h8a00;
17'h94d8:	data_out=16'h89fc;
17'h94d9:	data_out=16'h8a00;
17'h94da:	data_out=16'h9fb;
17'h94db:	data_out=16'h89c7;
17'h94dc:	data_out=16'h919;
17'h94dd:	data_out=16'h897c;
17'h94de:	data_out=16'ha00;
17'h94df:	data_out=16'h6b5;
17'h94e0:	data_out=16'h2b8;
17'h94e1:	data_out=16'h8a00;
17'h94e2:	data_out=16'h9ce;
17'h94e3:	data_out=16'ha00;
17'h94e4:	data_out=16'h9f1;
17'h94e5:	data_out=16'h9d9;
17'h94e6:	data_out=16'h89f6;
17'h94e7:	data_out=16'h89f5;
17'h94e8:	data_out=16'h89fc;
17'h94e9:	data_out=16'h89ff;
17'h94ea:	data_out=16'h89fd;
17'h94eb:	data_out=16'h89ff;
17'h94ec:	data_out=16'h89f8;
17'h94ed:	data_out=16'ha00;
17'h94ee:	data_out=16'h89fd;
17'h94ef:	data_out=16'h8a00;
17'h94f0:	data_out=16'h89fd;
17'h94f1:	data_out=16'h8ba;
17'h94f2:	data_out=16'h8a00;
17'h94f3:	data_out=16'h8a00;
17'h94f4:	data_out=16'h8a00;
17'h94f5:	data_out=16'h8a00;
17'h94f6:	data_out=16'h9fc;
17'h94f7:	data_out=16'h8a00;
17'h94f8:	data_out=16'h8a00;
17'h94f9:	data_out=16'h26b;
17'h94fa:	data_out=16'h9fa;
17'h94fb:	data_out=16'h89fc;
17'h94fc:	data_out=16'h89ff;
17'h94fd:	data_out=16'h8489;
17'h94fe:	data_out=16'ha00;
17'h94ff:	data_out=16'h8a00;
17'h9500:	data_out=16'h89fc;
17'h9501:	data_out=16'h9fd;
17'h9502:	data_out=16'h8a00;
17'h9503:	data_out=16'h89e2;
17'h9504:	data_out=16'h8a00;
17'h9505:	data_out=16'h8a00;
17'h9506:	data_out=16'ha00;
17'h9507:	data_out=16'h8a00;
17'h9508:	data_out=16'h892a;
17'h9509:	data_out=16'h9f9;
17'h950a:	data_out=16'h761;
17'h950b:	data_out=16'ha00;
17'h950c:	data_out=16'h89f5;
17'h950d:	data_out=16'h8a00;
17'h950e:	data_out=16'h1f1;
17'h950f:	data_out=16'h89ff;
17'h9510:	data_out=16'he;
17'h9511:	data_out=16'ha00;
17'h9512:	data_out=16'h7ad;
17'h9513:	data_out=16'h5fb;
17'h9514:	data_out=16'h9eb;
17'h9515:	data_out=16'h8a00;
17'h9516:	data_out=16'h8a00;
17'h9517:	data_out=16'h9e8;
17'h9518:	data_out=16'h8a00;
17'h9519:	data_out=16'h8944;
17'h951a:	data_out=16'h8a00;
17'h951b:	data_out=16'h8929;
17'h951c:	data_out=16'h89ec;
17'h951d:	data_out=16'ha00;
17'h951e:	data_out=16'h9c9;
17'h951f:	data_out=16'h9e7;
17'h9520:	data_out=16'h810e;
17'h9521:	data_out=16'h1f0;
17'h9522:	data_out=16'h832f;
17'h9523:	data_out=16'h8a00;
17'h9524:	data_out=16'h89ff;
17'h9525:	data_out=16'h89e5;
17'h9526:	data_out=16'h874b;
17'h9527:	data_out=16'h9fc;
17'h9528:	data_out=16'h434;
17'h9529:	data_out=16'h89d5;
17'h952a:	data_out=16'h8a00;
17'h952b:	data_out=16'ha00;
17'h952c:	data_out=16'h8a00;
17'h952d:	data_out=16'ha00;
17'h952e:	data_out=16'h9ee;
17'h952f:	data_out=16'h45f;
17'h9530:	data_out=16'h8a00;
17'h9531:	data_out=16'h9c8;
17'h9532:	data_out=16'h89fb;
17'h9533:	data_out=16'h9fb;
17'h9534:	data_out=16'ha00;
17'h9535:	data_out=16'h85e9;
17'h9536:	data_out=16'h84d0;
17'h9537:	data_out=16'h89fe;
17'h9538:	data_out=16'ha00;
17'h9539:	data_out=16'h9fb;
17'h953a:	data_out=16'h2dc;
17'h953b:	data_out=16'h89b2;
17'h953c:	data_out=16'h83d8;
17'h953d:	data_out=16'h897d;
17'h953e:	data_out=16'h43e;
17'h953f:	data_out=16'h8a00;
17'h9540:	data_out=16'h89df;
17'h9541:	data_out=16'h8a00;
17'h9542:	data_out=16'h89d3;
17'h9543:	data_out=16'h8a00;
17'h9544:	data_out=16'h81dc;
17'h9545:	data_out=16'h8a00;
17'h9546:	data_out=16'h9ff;
17'h9547:	data_out=16'h9b4;
17'h9548:	data_out=16'h9ff;
17'h9549:	data_out=16'h89bd;
17'h954a:	data_out=16'h9c6;
17'h954b:	data_out=16'h3b7;
17'h954c:	data_out=16'h89ff;
17'h954d:	data_out=16'h8e9;
17'h954e:	data_out=16'h7cb;
17'h954f:	data_out=16'h896b;
17'h9550:	data_out=16'h89f7;
17'h9551:	data_out=16'h8a00;
17'h9552:	data_out=16'h8a00;
17'h9553:	data_out=16'h9e5;
17'h9554:	data_out=16'h9f2;
17'h9555:	data_out=16'h8a00;
17'h9556:	data_out=16'h8a00;
17'h9557:	data_out=16'h89f9;
17'h9558:	data_out=16'h8a00;
17'h9559:	data_out=16'h89cc;
17'h955a:	data_out=16'h994;
17'h955b:	data_out=16'h8360;
17'h955c:	data_out=16'hfe;
17'h955d:	data_out=16'h87ae;
17'h955e:	data_out=16'h793;
17'h955f:	data_out=16'h852f;
17'h9560:	data_out=16'h9e0;
17'h9561:	data_out=16'h89ff;
17'h9562:	data_out=16'h9f0;
17'h9563:	data_out=16'h9fb;
17'h9564:	data_out=16'ha00;
17'h9565:	data_out=16'h9fd;
17'h9566:	data_out=16'h89c0;
17'h9567:	data_out=16'h89d9;
17'h9568:	data_out=16'h2ce;
17'h9569:	data_out=16'h8a00;
17'h956a:	data_out=16'h1ad;
17'h956b:	data_out=16'h89f1;
17'h956c:	data_out=16'h89fe;
17'h956d:	data_out=16'h9fc;
17'h956e:	data_out=16'h1aa;
17'h956f:	data_out=16'h89ff;
17'h9570:	data_out=16'h1cf;
17'h9571:	data_out=16'h803a;
17'h9572:	data_out=16'h89d7;
17'h9573:	data_out=16'h8a00;
17'h9574:	data_out=16'h8a00;
17'h9575:	data_out=16'h8a00;
17'h9576:	data_out=16'h9fc;
17'h9577:	data_out=16'h89e2;
17'h9578:	data_out=16'h8a00;
17'h9579:	data_out=16'h8a00;
17'h957a:	data_out=16'h9f9;
17'h957b:	data_out=16'h43f;
17'h957c:	data_out=16'h8a00;
17'h957d:	data_out=16'h8227;
17'h957e:	data_out=16'ha00;
17'h957f:	data_out=16'h8a00;
17'h9580:	data_out=16'h89f9;
17'h9581:	data_out=16'ha00;
17'h9582:	data_out=16'h89ff;
17'h9583:	data_out=16'h89ed;
17'h9584:	data_out=16'h8a00;
17'h9585:	data_out=16'h8a00;
17'h9586:	data_out=16'ha00;
17'h9587:	data_out=16'h8a00;
17'h9588:	data_out=16'h89d0;
17'h9589:	data_out=16'h8c;
17'h958a:	data_out=16'h982;
17'h958b:	data_out=16'ha00;
17'h958c:	data_out=16'h89dc;
17'h958d:	data_out=16'h8a00;
17'h958e:	data_out=16'h80b;
17'h958f:	data_out=16'h89ff;
17'h9590:	data_out=16'h836d;
17'h9591:	data_out=16'ha00;
17'h9592:	data_out=16'h32d;
17'h9593:	data_out=16'h9ac;
17'h9594:	data_out=16'h9d9;
17'h9595:	data_out=16'h8a00;
17'h9596:	data_out=16'h8a00;
17'h9597:	data_out=16'h9e5;
17'h9598:	data_out=16'h8a00;
17'h9599:	data_out=16'h9f9;
17'h959a:	data_out=16'h8a00;
17'h959b:	data_out=16'h8967;
17'h959c:	data_out=16'h89fe;
17'h959d:	data_out=16'ha00;
17'h959e:	data_out=16'h869b;
17'h959f:	data_out=16'h9bb;
17'h95a0:	data_out=16'h8684;
17'h95a1:	data_out=16'h86d;
17'h95a2:	data_out=16'h9ff;
17'h95a3:	data_out=16'h511;
17'h95a4:	data_out=16'h4af;
17'h95a5:	data_out=16'h89ec;
17'h95a6:	data_out=16'h87f1;
17'h95a7:	data_out=16'h379;
17'h95a8:	data_out=16'h9e7;
17'h95a9:	data_out=16'h89d2;
17'h95aa:	data_out=16'h8950;
17'h95ab:	data_out=16'ha00;
17'h95ac:	data_out=16'h8a00;
17'h95ad:	data_out=16'ha00;
17'h95ae:	data_out=16'ha00;
17'h95af:	data_out=16'h82de;
17'h95b0:	data_out=16'h89ce;
17'h95b1:	data_out=16'h9f4;
17'h95b2:	data_out=16'h89aa;
17'h95b3:	data_out=16'h9ec;
17'h95b4:	data_out=16'ha00;
17'h95b5:	data_out=16'h86f7;
17'h95b6:	data_out=16'h870e;
17'h95b7:	data_out=16'h571;
17'h95b8:	data_out=16'ha00;
17'h95b9:	data_out=16'h9d5;
17'h95ba:	data_out=16'h8319;
17'h95bb:	data_out=16'h88c3;
17'h95bc:	data_out=16'h9f7;
17'h95bd:	data_out=16'h896b;
17'h95be:	data_out=16'h9f1;
17'h95bf:	data_out=16'h8a00;
17'h95c0:	data_out=16'h89c2;
17'h95c1:	data_out=16'h8a00;
17'h95c2:	data_out=16'h89cb;
17'h95c3:	data_out=16'h8a00;
17'h95c4:	data_out=16'h86e1;
17'h95c5:	data_out=16'h8a00;
17'h95c6:	data_out=16'ha00;
17'h95c7:	data_out=16'h81a7;
17'h95c8:	data_out=16'ha00;
17'h95c9:	data_out=16'h89c1;
17'h95ca:	data_out=16'h43;
17'h95cb:	data_out=16'h882e;
17'h95cc:	data_out=16'h89fc;
17'h95cd:	data_out=16'ha00;
17'h95ce:	data_out=16'h9ab;
17'h95cf:	data_out=16'h8729;
17'h95d0:	data_out=16'h89fe;
17'h95d1:	data_out=16'h8a00;
17'h95d2:	data_out=16'h89fe;
17'h95d3:	data_out=16'h9fd;
17'h95d4:	data_out=16'h8112;
17'h95d5:	data_out=16'h89fa;
17'h95d6:	data_out=16'h89fd;
17'h95d7:	data_out=16'h89f7;
17'h95d8:	data_out=16'h8a00;
17'h95d9:	data_out=16'h899c;
17'h95da:	data_out=16'h7ed;
17'h95db:	data_out=16'h82f1;
17'h95dc:	data_out=16'h5f2;
17'h95dd:	data_out=16'h888d;
17'h95de:	data_out=16'h8071;
17'h95df:	data_out=16'h8731;
17'h95e0:	data_out=16'h9d7;
17'h95e1:	data_out=16'h89ad;
17'h95e2:	data_out=16'h9dd;
17'h95e3:	data_out=16'h9fc;
17'h95e4:	data_out=16'ha00;
17'h95e5:	data_out=16'ha00;
17'h95e6:	data_out=16'h8971;
17'h95e7:	data_out=16'h896f;
17'h95e8:	data_out=16'h913;
17'h95e9:	data_out=16'h8a00;
17'h95ea:	data_out=16'h7ef;
17'h95eb:	data_out=16'h899e;
17'h95ec:	data_out=16'h89ff;
17'h95ed:	data_out=16'h9fc;
17'h95ee:	data_out=16'h7eb;
17'h95ef:	data_out=16'h89fd;
17'h95f0:	data_out=16'h7f0;
17'h95f1:	data_out=16'h89e1;
17'h95f2:	data_out=16'h890a;
17'h95f3:	data_out=16'h8971;
17'h95f4:	data_out=16'h89c8;
17'h95f5:	data_out=16'h89fe;
17'h95f6:	data_out=16'h9fc;
17'h95f7:	data_out=16'h89fe;
17'h95f8:	data_out=16'h8a00;
17'h95f9:	data_out=16'h8a00;
17'h95fa:	data_out=16'h9f5;
17'h95fb:	data_out=16'h9f3;
17'h95fc:	data_out=16'h8a00;
17'h95fd:	data_out=16'h83b7;
17'h95fe:	data_out=16'ha00;
17'h95ff:	data_out=16'h8a00;
17'h9600:	data_out=16'h89e3;
17'h9601:	data_out=16'ha00;
17'h9602:	data_out=16'h89ff;
17'h9603:	data_out=16'h89fa;
17'h9604:	data_out=16'h89d2;
17'h9605:	data_out=16'h89f1;
17'h9606:	data_out=16'ha00;
17'h9607:	data_out=16'h89f5;
17'h9608:	data_out=16'h898b;
17'h9609:	data_out=16'h8725;
17'h960a:	data_out=16'h8731;
17'h960b:	data_out=16'h9fb;
17'h960c:	data_out=16'h88e9;
17'h960d:	data_out=16'h8a00;
17'h960e:	data_out=16'h421;
17'h960f:	data_out=16'h89ec;
17'h9610:	data_out=16'h8859;
17'h9611:	data_out=16'ha00;
17'h9612:	data_out=16'h821c;
17'h9613:	data_out=16'h9cc;
17'h9614:	data_out=16'h85a3;
17'h9615:	data_out=16'h8a00;
17'h9616:	data_out=16'h8a00;
17'h9617:	data_out=16'h9fc;
17'h9618:	data_out=16'h8a00;
17'h9619:	data_out=16'h9fd;
17'h961a:	data_out=16'h89d0;
17'h961b:	data_out=16'h8913;
17'h961c:	data_out=16'h89fe;
17'h961d:	data_out=16'ha00;
17'h961e:	data_out=16'h8941;
17'h961f:	data_out=16'h475;
17'h9620:	data_out=16'h8925;
17'h9621:	data_out=16'h396;
17'h9622:	data_out=16'h9e2;
17'h9623:	data_out=16'ha00;
17'h9624:	data_out=16'ha00;
17'h9625:	data_out=16'h8a00;
17'h9626:	data_out=16'h8642;
17'h9627:	data_out=16'h813a;
17'h9628:	data_out=16'h4d7;
17'h9629:	data_out=16'h89fe;
17'h962a:	data_out=16'h883a;
17'h962b:	data_out=16'ha00;
17'h962c:	data_out=16'h8a00;
17'h962d:	data_out=16'ha00;
17'h962e:	data_out=16'ha00;
17'h962f:	data_out=16'h8652;
17'h9630:	data_out=16'h89c6;
17'h9631:	data_out=16'h891f;
17'h9632:	data_out=16'h8970;
17'h9633:	data_out=16'h873c;
17'h9634:	data_out=16'ha00;
17'h9635:	data_out=16'h8973;
17'h9636:	data_out=16'h87e5;
17'h9637:	data_out=16'h881;
17'h9638:	data_out=16'ha00;
17'h9639:	data_out=16'h8934;
17'h963a:	data_out=16'h89ff;
17'h963b:	data_out=16'h8973;
17'h963c:	data_out=16'h9eb;
17'h963d:	data_out=16'h89ef;
17'h963e:	data_out=16'h4ec;
17'h963f:	data_out=16'h89f5;
17'h9640:	data_out=16'h899e;
17'h9641:	data_out=16'h8a00;
17'h9642:	data_out=16'h88a2;
17'h9643:	data_out=16'h8a00;
17'h9644:	data_out=16'h8984;
17'h9645:	data_out=16'h8a00;
17'h9646:	data_out=16'ha00;
17'h9647:	data_out=16'h899a;
17'h9648:	data_out=16'ha00;
17'h9649:	data_out=16'h8a00;
17'h964a:	data_out=16'h4cc;
17'h964b:	data_out=16'h82cf;
17'h964c:	data_out=16'h89ff;
17'h964d:	data_out=16'h9ff;
17'h964e:	data_out=16'h9f3;
17'h964f:	data_out=16'h8906;
17'h9650:	data_out=16'h8a00;
17'h9651:	data_out=16'h8a00;
17'h9652:	data_out=16'h89fa;
17'h9653:	data_out=16'ha00;
17'h9654:	data_out=16'h85ac;
17'h9655:	data_out=16'h89fd;
17'h9656:	data_out=16'h89ff;
17'h9657:	data_out=16'h8a00;
17'h9658:	data_out=16'h8a00;
17'h9659:	data_out=16'h89b6;
17'h965a:	data_out=16'h9de;
17'h965b:	data_out=16'h86f8;
17'h965c:	data_out=16'h60;
17'h965d:	data_out=16'h8942;
17'h965e:	data_out=16'h852d;
17'h965f:	data_out=16'h88e2;
17'h9660:	data_out=16'h9ea;
17'h9661:	data_out=16'h898d;
17'h9662:	data_out=16'ha00;
17'h9663:	data_out=16'h8d;
17'h9664:	data_out=16'ha00;
17'h9665:	data_out=16'h9ff;
17'h9666:	data_out=16'h897a;
17'h9667:	data_out=16'h8941;
17'h9668:	data_out=16'h3cf;
17'h9669:	data_out=16'h89f5;
17'h966a:	data_out=16'h490;
17'h966b:	data_out=16'h89b8;
17'h966c:	data_out=16'h89e3;
17'h966d:	data_out=16'h811c;
17'h966e:	data_out=16'h48b;
17'h966f:	data_out=16'h89b1;
17'h9670:	data_out=16'h449;
17'h9671:	data_out=16'h89b8;
17'h9672:	data_out=16'h89c1;
17'h9673:	data_out=16'h89b0;
17'h9674:	data_out=16'h89b5;
17'h9675:	data_out=16'h89fe;
17'h9676:	data_out=16'h9fc;
17'h9677:	data_out=16'h89ff;
17'h9678:	data_out=16'h8a00;
17'h9679:	data_out=16'h8a00;
17'h967a:	data_out=16'h85da;
17'h967b:	data_out=16'h4f1;
17'h967c:	data_out=16'h8a00;
17'h967d:	data_out=16'h8a00;
17'h967e:	data_out=16'ha00;
17'h967f:	data_out=16'h8a00;
17'h9680:	data_out=16'h89c1;
17'h9681:	data_out=16'h9e4;
17'h9682:	data_out=16'h89fd;
17'h9683:	data_out=16'h89fc;
17'h9684:	data_out=16'h89e3;
17'h9685:	data_out=16'h8a00;
17'h9686:	data_out=16'h9fe;
17'h9687:	data_out=16'h89a9;
17'h9688:	data_out=16'h89a7;
17'h9689:	data_out=16'h8914;
17'h968a:	data_out=16'h88e8;
17'h968b:	data_out=16'ha00;
17'h968c:	data_out=16'h849c;
17'h968d:	data_out=16'h8a00;
17'h968e:	data_out=16'h631;
17'h968f:	data_out=16'h89df;
17'h9690:	data_out=16'h89f4;
17'h9691:	data_out=16'h8493;
17'h9692:	data_out=16'h8261;
17'h9693:	data_out=16'h9a8;
17'h9694:	data_out=16'h89bf;
17'h9695:	data_out=16'h8a00;
17'h9696:	data_out=16'h8a00;
17'h9697:	data_out=16'h891e;
17'h9698:	data_out=16'h8a00;
17'h9699:	data_out=16'h4d6;
17'h969a:	data_out=16'h89fd;
17'h969b:	data_out=16'h89c6;
17'h969c:	data_out=16'h8a00;
17'h969d:	data_out=16'ha00;
17'h969e:	data_out=16'h89f8;
17'h969f:	data_out=16'h8987;
17'h96a0:	data_out=16'h89d8;
17'h96a1:	data_out=16'h545;
17'h96a2:	data_out=16'h9d7;
17'h96a3:	data_out=16'ha00;
17'h96a4:	data_out=16'ha00;
17'h96a5:	data_out=16'h85c9;
17'h96a6:	data_out=16'h9f9;
17'h96a7:	data_out=16'h883e;
17'h96a8:	data_out=16'h474;
17'h96a9:	data_out=16'h8a00;
17'h96aa:	data_out=16'h8814;
17'h96ab:	data_out=16'ha00;
17'h96ac:	data_out=16'h8a00;
17'h96ad:	data_out=16'ha00;
17'h96ae:	data_out=16'ha00;
17'h96af:	data_out=16'h8979;
17'h96b0:	data_out=16'h8996;
17'h96b1:	data_out=16'h898e;
17'h96b2:	data_out=16'h8671;
17'h96b3:	data_out=16'h89f9;
17'h96b4:	data_out=16'ha00;
17'h96b5:	data_out=16'h8987;
17'h96b6:	data_out=16'h8970;
17'h96b7:	data_out=16'h65;
17'h96b8:	data_out=16'ha00;
17'h96b9:	data_out=16'h89fb;
17'h96ba:	data_out=16'h89f8;
17'h96bb:	data_out=16'h897d;
17'h96bc:	data_out=16'h9e2;
17'h96bd:	data_out=16'h89fb;
17'h96be:	data_out=16'h472;
17'h96bf:	data_out=16'h8a00;
17'h96c0:	data_out=16'h89d3;
17'h96c1:	data_out=16'h89ea;
17'h96c2:	data_out=16'h9ff;
17'h96c3:	data_out=16'h8a00;
17'h96c4:	data_out=16'h89a5;
17'h96c5:	data_out=16'h8a00;
17'h96c6:	data_out=16'ha00;
17'h96c7:	data_out=16'h89d0;
17'h96c8:	data_out=16'ha00;
17'h96c9:	data_out=16'h89e7;
17'h96ca:	data_out=16'h852d;
17'h96cb:	data_out=16'ha00;
17'h96cc:	data_out=16'h5c9;
17'h96cd:	data_out=16'h9db;
17'h96ce:	data_out=16'h9fa;
17'h96cf:	data_out=16'h88d5;
17'h96d0:	data_out=16'h8a00;
17'h96d1:	data_out=16'h8a00;
17'h96d2:	data_out=16'h198;
17'h96d3:	data_out=16'h43e;
17'h96d4:	data_out=16'h8988;
17'h96d5:	data_out=16'h89fe;
17'h96d6:	data_out=16'h89f0;
17'h96d7:	data_out=16'h8a00;
17'h96d8:	data_out=16'h8a00;
17'h96d9:	data_out=16'h89ea;
17'h96da:	data_out=16'h82f;
17'h96db:	data_out=16'h8979;
17'h96dc:	data_out=16'h89a1;
17'h96dd:	data_out=16'h89b9;
17'h96de:	data_out=16'h88f0;
17'h96df:	data_out=16'h89cd;
17'h96e0:	data_out=16'h9fb;
17'h96e1:	data_out=16'h89b0;
17'h96e2:	data_out=16'h817c;
17'h96e3:	data_out=16'h89af;
17'h96e4:	data_out=16'ha00;
17'h96e5:	data_out=16'h84a4;
17'h96e6:	data_out=16'h89c2;
17'h96e7:	data_out=16'h89bb;
17'h96e8:	data_out=16'h4d9;
17'h96e9:	data_out=16'h89dc;
17'h96ea:	data_out=16'h6cf;
17'h96eb:	data_out=16'h8a00;
17'h96ec:	data_out=16'h89bd;
17'h96ed:	data_out=16'h89ba;
17'h96ee:	data_out=16'h6cd;
17'h96ef:	data_out=16'h89ec;
17'h96f0:	data_out=16'h677;
17'h96f1:	data_out=16'h899e;
17'h96f2:	data_out=16'h89f2;
17'h96f3:	data_out=16'h89c4;
17'h96f4:	data_out=16'h8913;
17'h96f5:	data_out=16'h8a00;
17'h96f6:	data_out=16'h9ff;
17'h96f7:	data_out=16'h89fe;
17'h96f8:	data_out=16'h8a00;
17'h96f9:	data_out=16'h8a00;
17'h96fa:	data_out=16'h8995;
17'h96fb:	data_out=16'h472;
17'h96fc:	data_out=16'h8a00;
17'h96fd:	data_out=16'h8a00;
17'h96fe:	data_out=16'ha00;
17'h96ff:	data_out=16'h8a00;
17'h9700:	data_out=16'h89c5;
17'h9701:	data_out=16'ha00;
17'h9702:	data_out=16'h89fe;
17'h9703:	data_out=16'h8a00;
17'h9704:	data_out=16'h89f9;
17'h9705:	data_out=16'h8a00;
17'h9706:	data_out=16'ha00;
17'h9707:	data_out=16'h8904;
17'h9708:	data_out=16'h89bc;
17'h9709:	data_out=16'h898e;
17'h970a:	data_out=16'h9fd;
17'h970b:	data_out=16'h36e;
17'h970c:	data_out=16'h38e;
17'h970d:	data_out=16'h8a00;
17'h970e:	data_out=16'h8226;
17'h970f:	data_out=16'h89e2;
17'h9710:	data_out=16'h8a00;
17'h9711:	data_out=16'h8986;
17'h9712:	data_out=16'h8377;
17'h9713:	data_out=16'h52c;
17'h9714:	data_out=16'h89ff;
17'h9715:	data_out=16'h8a00;
17'h9716:	data_out=16'h8a00;
17'h9717:	data_out=16'h89cb;
17'h9718:	data_out=16'h8a00;
17'h9719:	data_out=16'h89ee;
17'h971a:	data_out=16'h8a00;
17'h971b:	data_out=16'h89f0;
17'h971c:	data_out=16'h8a00;
17'h971d:	data_out=16'h92a;
17'h971e:	data_out=16'h8a00;
17'h971f:	data_out=16'h89fe;
17'h9720:	data_out=16'h8a00;
17'h9721:	data_out=16'h8397;
17'h9722:	data_out=16'h820e;
17'h9723:	data_out=16'ha00;
17'h9724:	data_out=16'ha00;
17'h9725:	data_out=16'h8266;
17'h9726:	data_out=16'ha00;
17'h9727:	data_out=16'h89b9;
17'h9728:	data_out=16'h8654;
17'h9729:	data_out=16'h89f8;
17'h972a:	data_out=16'h8871;
17'h972b:	data_out=16'h89b3;
17'h972c:	data_out=16'h8a00;
17'h972d:	data_out=16'ha00;
17'h972e:	data_out=16'h595;
17'h972f:	data_out=16'h89e1;
17'h9730:	data_out=16'h8513;
17'h9731:	data_out=16'h89d7;
17'h9732:	data_out=16'h8538;
17'h9733:	data_out=16'h8a00;
17'h9734:	data_out=16'ha00;
17'h9735:	data_out=16'h89dd;
17'h9736:	data_out=16'h89c3;
17'h9737:	data_out=16'h89ec;
17'h9738:	data_out=16'h9af;
17'h9739:	data_out=16'h8a00;
17'h973a:	data_out=16'h89fe;
17'h973b:	data_out=16'h89bf;
17'h973c:	data_out=16'h84c1;
17'h973d:	data_out=16'h8a00;
17'h973e:	data_out=16'h866a;
17'h973f:	data_out=16'h8a00;
17'h9740:	data_out=16'h89fe;
17'h9741:	data_out=16'h89ed;
17'h9742:	data_out=16'ha00;
17'h9743:	data_out=16'h8a00;
17'h9744:	data_out=16'h89fb;
17'h9745:	data_out=16'h8a00;
17'h9746:	data_out=16'ha00;
17'h9747:	data_out=16'h89dd;
17'h9748:	data_out=16'h57f;
17'h9749:	data_out=16'h8541;
17'h974a:	data_out=16'h898e;
17'h974b:	data_out=16'ha00;
17'h974c:	data_out=16'h986;
17'h974d:	data_out=16'h82e2;
17'h974e:	data_out=16'h266;
17'h974f:	data_out=16'h9fd;
17'h9750:	data_out=16'h8a00;
17'h9751:	data_out=16'h8a00;
17'h9752:	data_out=16'h9fa;
17'h9753:	data_out=16'h89b6;
17'h9754:	data_out=16'h89e4;
17'h9755:	data_out=16'h8a00;
17'h9756:	data_out=16'h89de;
17'h9757:	data_out=16'h8a00;
17'h9758:	data_out=16'h8a00;
17'h9759:	data_out=16'h89ff;
17'h975a:	data_out=16'h89ef;
17'h975b:	data_out=16'h89e9;
17'h975c:	data_out=16'h8a00;
17'h975d:	data_out=16'h89ed;
17'h975e:	data_out=16'h89d0;
17'h975f:	data_out=16'h89f5;
17'h9760:	data_out=16'ha00;
17'h9761:	data_out=16'h89eb;
17'h9762:	data_out=16'h8967;
17'h9763:	data_out=16'h89ff;
17'h9764:	data_out=16'ha00;
17'h9765:	data_out=16'h89d5;
17'h9766:	data_out=16'h8a00;
17'h9767:	data_out=16'h89fd;
17'h9768:	data_out=16'h84af;
17'h9769:	data_out=16'h89d2;
17'h976a:	data_out=16'h8180;
17'h976b:	data_out=16'h8a00;
17'h976c:	data_out=16'h895a;
17'h976d:	data_out=16'h8a00;
17'h976e:	data_out=16'h817f;
17'h976f:	data_out=16'h8a00;
17'h9770:	data_out=16'h81cc;
17'h9771:	data_out=16'h89d3;
17'h9772:	data_out=16'h8a00;
17'h9773:	data_out=16'h89ef;
17'h9774:	data_out=16'h821c;
17'h9775:	data_out=16'h8a00;
17'h9776:	data_out=16'h12;
17'h9777:	data_out=16'h8a00;
17'h9778:	data_out=16'h8a00;
17'h9779:	data_out=16'h8a00;
17'h977a:	data_out=16'h89ff;
17'h977b:	data_out=16'h866f;
17'h977c:	data_out=16'h8a00;
17'h977d:	data_out=16'h8a00;
17'h977e:	data_out=16'ha00;
17'h977f:	data_out=16'h8a00;
17'h9780:	data_out=16'ha00;
17'h9781:	data_out=16'ha00;
17'h9782:	data_out=16'h89f1;
17'h9783:	data_out=16'h8a00;
17'h9784:	data_out=16'h6cc;
17'h9785:	data_out=16'h8a00;
17'h9786:	data_out=16'ha00;
17'h9787:	data_out=16'h89f3;
17'h9788:	data_out=16'h85fd;
17'h9789:	data_out=16'h89ff;
17'h978a:	data_out=16'ha00;
17'h978b:	data_out=16'h89e6;
17'h978c:	data_out=16'h888a;
17'h978d:	data_out=16'h8a00;
17'h978e:	data_out=16'ha00;
17'h978f:	data_out=16'h89f5;
17'h9790:	data_out=16'h8a00;
17'h9791:	data_out=16'h851e;
17'h9792:	data_out=16'h8a00;
17'h9793:	data_out=16'h89ff;
17'h9794:	data_out=16'h8a00;
17'h9795:	data_out=16'h8a00;
17'h9796:	data_out=16'h8a00;
17'h9797:	data_out=16'h8a00;
17'h9798:	data_out=16'h8a00;
17'h9799:	data_out=16'h8a00;
17'h979a:	data_out=16'h89ff;
17'h979b:	data_out=16'h8a00;
17'h979c:	data_out=16'h8a00;
17'h979d:	data_out=16'h5ba;
17'h979e:	data_out=16'h8a00;
17'h979f:	data_out=16'h8a00;
17'h97a0:	data_out=16'h8a00;
17'h97a1:	data_out=16'ha00;
17'h97a2:	data_out=16'h89f9;
17'h97a3:	data_out=16'ha00;
17'h97a4:	data_out=16'ha00;
17'h97a5:	data_out=16'h80b9;
17'h97a6:	data_out=16'ha00;
17'h97a7:	data_out=16'h89f6;
17'h97a8:	data_out=16'h9f7;
17'h97a9:	data_out=16'h8a00;
17'h97aa:	data_out=16'h892c;
17'h97ab:	data_out=16'h8a00;
17'h97ac:	data_out=16'h8a00;
17'h97ad:	data_out=16'ha00;
17'h97ae:	data_out=16'h89d9;
17'h97af:	data_out=16'h8a00;
17'h97b0:	data_out=16'ha00;
17'h97b1:	data_out=16'h82af;
17'h97b2:	data_out=16'ha00;
17'h97b3:	data_out=16'h8a00;
17'h97b4:	data_out=16'ha00;
17'h97b5:	data_out=16'h8902;
17'h97b6:	data_out=16'h89e7;
17'h97b7:	data_out=16'h89f5;
17'h97b8:	data_out=16'h9d1;
17'h97b9:	data_out=16'h8a00;
17'h97ba:	data_out=16'h8a00;
17'h97bb:	data_out=16'h9f6;
17'h97bc:	data_out=16'h8917;
17'h97bd:	data_out=16'h89fe;
17'h97be:	data_out=16'h9f7;
17'h97bf:	data_out=16'h8a00;
17'h97c0:	data_out=16'h89d8;
17'h97c1:	data_out=16'h89e7;
17'h97c2:	data_out=16'ha00;
17'h97c3:	data_out=16'h8a00;
17'h97c4:	data_out=16'h89fc;
17'h97c5:	data_out=16'h8a00;
17'h97c6:	data_out=16'ha00;
17'h97c7:	data_out=16'h8a00;
17'h97c8:	data_out=16'h8985;
17'h97c9:	data_out=16'h809f;
17'h97ca:	data_out=16'h89f4;
17'h97cb:	data_out=16'ha00;
17'h97cc:	data_out=16'ha00;
17'h97cd:	data_out=16'h89fe;
17'h97ce:	data_out=16'h872d;
17'h97cf:	data_out=16'ha00;
17'h97d0:	data_out=16'h8a00;
17'h97d1:	data_out=16'h8a00;
17'h97d2:	data_out=16'ha00;
17'h97d3:	data_out=16'h8a00;
17'h97d4:	data_out=16'h89ff;
17'h97d5:	data_out=16'h8a00;
17'h97d6:	data_out=16'ha00;
17'h97d7:	data_out=16'h89fb;
17'h97d8:	data_out=16'h8a00;
17'h97d9:	data_out=16'h82d5;
17'h97da:	data_out=16'h8a00;
17'h97db:	data_out=16'h7a4;
17'h97dc:	data_out=16'h8a00;
17'h97dd:	data_out=16'h89f1;
17'h97de:	data_out=16'h89ff;
17'h97df:	data_out=16'h89fd;
17'h97e0:	data_out=16'ha00;
17'h97e1:	data_out=16'h29b;
17'h97e2:	data_out=16'h8a00;
17'h97e3:	data_out=16'h8a00;
17'h97e4:	data_out=16'ha00;
17'h97e5:	data_out=16'h8a00;
17'h97e6:	data_out=16'h8a00;
17'h97e7:	data_out=16'h8a00;
17'h97e8:	data_out=16'h9fe;
17'h97e9:	data_out=16'h80e8;
17'h97ea:	data_out=16'ha00;
17'h97eb:	data_out=16'h8a00;
17'h97ec:	data_out=16'ha00;
17'h97ed:	data_out=16'h8a00;
17'h97ee:	data_out=16'ha00;
17'h97ef:	data_out=16'h8a00;
17'h97f0:	data_out=16'ha00;
17'h97f1:	data_out=16'h89f3;
17'h97f2:	data_out=16'h8377;
17'h97f3:	data_out=16'h67c;
17'h97f4:	data_out=16'ha00;
17'h97f5:	data_out=16'h8298;
17'h97f6:	data_out=16'h8a00;
17'h97f7:	data_out=16'h8a00;
17'h97f8:	data_out=16'h8a00;
17'h97f9:	data_out=16'h89ee;
17'h97fa:	data_out=16'h8a00;
17'h97fb:	data_out=16'h9f6;
17'h97fc:	data_out=16'h8a00;
17'h97fd:	data_out=16'h8a00;
17'h97fe:	data_out=16'h844b;
17'h97ff:	data_out=16'h8a00;
17'h9800:	data_out=16'ha00;
17'h9801:	data_out=16'ha00;
17'h9802:	data_out=16'ha00;
17'h9803:	data_out=16'h8a00;
17'h9804:	data_out=16'ha00;
17'h9805:	data_out=16'h156;
17'h9806:	data_out=16'h89f8;
17'h9807:	data_out=16'h8a00;
17'h9808:	data_out=16'ha00;
17'h9809:	data_out=16'h8a00;
17'h980a:	data_out=16'ha00;
17'h980b:	data_out=16'h8a00;
17'h980c:	data_out=16'h89c9;
17'h980d:	data_out=16'h89f2;
17'h980e:	data_out=16'ha00;
17'h980f:	data_out=16'h16c;
17'h9810:	data_out=16'h8a00;
17'h9811:	data_out=16'h479;
17'h9812:	data_out=16'h89f2;
17'h9813:	data_out=16'h89fc;
17'h9814:	data_out=16'h8a00;
17'h9815:	data_out=16'ha00;
17'h9816:	data_out=16'h6c5;
17'h9817:	data_out=16'h8a00;
17'h9818:	data_out=16'h9fb;
17'h9819:	data_out=16'h8a00;
17'h981a:	data_out=16'ha00;
17'h981b:	data_out=16'h8a00;
17'h981c:	data_out=16'h433;
17'h981d:	data_out=16'ha00;
17'h981e:	data_out=16'h8a00;
17'h981f:	data_out=16'h8a00;
17'h9820:	data_out=16'h89ed;
17'h9821:	data_out=16'ha00;
17'h9822:	data_out=16'h8a00;
17'h9823:	data_out=16'ha00;
17'h9824:	data_out=16'ha00;
17'h9825:	data_out=16'h83c5;
17'h9826:	data_out=16'ha00;
17'h9827:	data_out=16'h89de;
17'h9828:	data_out=16'ha00;
17'h9829:	data_out=16'h8a00;
17'h982a:	data_out=16'h8942;
17'h982b:	data_out=16'h8a00;
17'h982c:	data_out=16'h6d7;
17'h982d:	data_out=16'h8025;
17'h982e:	data_out=16'h8a00;
17'h982f:	data_out=16'h8a00;
17'h9830:	data_out=16'ha00;
17'h9831:	data_out=16'h76d;
17'h9832:	data_out=16'ha00;
17'h9833:	data_out=16'h8a00;
17'h9834:	data_out=16'ha00;
17'h9835:	data_out=16'ha00;
17'h9836:	data_out=16'h8b4;
17'h9837:	data_out=16'ha00;
17'h9838:	data_out=16'h87d;
17'h9839:	data_out=16'h8a00;
17'h983a:	data_out=16'h8a00;
17'h983b:	data_out=16'ha00;
17'h983c:	data_out=16'h618;
17'h983d:	data_out=16'h85b5;
17'h983e:	data_out=16'ha00;
17'h983f:	data_out=16'h20a;
17'h9840:	data_out=16'ha00;
17'h9841:	data_out=16'h82c6;
17'h9842:	data_out=16'ha00;
17'h9843:	data_out=16'h8a00;
17'h9844:	data_out=16'h9cf;
17'h9845:	data_out=16'ha00;
17'h9846:	data_out=16'ha00;
17'h9847:	data_out=16'h8a00;
17'h9848:	data_out=16'h89f6;
17'h9849:	data_out=16'h8086;
17'h984a:	data_out=16'h8a00;
17'h984b:	data_out=16'h85ae;
17'h984c:	data_out=16'h927;
17'h984d:	data_out=16'h8a00;
17'h984e:	data_out=16'h83ea;
17'h984f:	data_out=16'ha00;
17'h9850:	data_out=16'h8a00;
17'h9851:	data_out=16'h89f7;
17'h9852:	data_out=16'ha00;
17'h9853:	data_out=16'h89ff;
17'h9854:	data_out=16'h89ec;
17'h9855:	data_out=16'h89ff;
17'h9856:	data_out=16'ha00;
17'h9857:	data_out=16'ha00;
17'h9858:	data_out=16'h9dd;
17'h9859:	data_out=16'ha00;
17'h985a:	data_out=16'h8a00;
17'h985b:	data_out=16'ha00;
17'h985c:	data_out=16'h89f0;
17'h985d:	data_out=16'h9ae;
17'h985e:	data_out=16'h89ff;
17'h985f:	data_out=16'hb1;
17'h9860:	data_out=16'h9f7;
17'h9861:	data_out=16'ha00;
17'h9862:	data_out=16'h8a00;
17'h9863:	data_out=16'h8a00;
17'h9864:	data_out=16'h8785;
17'h9865:	data_out=16'h8a00;
17'h9866:	data_out=16'h8a00;
17'h9867:	data_out=16'h8a00;
17'h9868:	data_out=16'ha00;
17'h9869:	data_out=16'h9f0;
17'h986a:	data_out=16'ha00;
17'h986b:	data_out=16'h89ff;
17'h986c:	data_out=16'ha00;
17'h986d:	data_out=16'h8a00;
17'h986e:	data_out=16'ha00;
17'h986f:	data_out=16'h89f1;
17'h9870:	data_out=16'ha00;
17'h9871:	data_out=16'h89ee;
17'h9872:	data_out=16'ha00;
17'h9873:	data_out=16'ha00;
17'h9874:	data_out=16'ha00;
17'h9875:	data_out=16'ha00;
17'h9876:	data_out=16'h8a00;
17'h9877:	data_out=16'h8a00;
17'h9878:	data_out=16'h8a00;
17'h9879:	data_out=16'h81e5;
17'h987a:	data_out=16'h8a00;
17'h987b:	data_out=16'ha00;
17'h987c:	data_out=16'h9fd;
17'h987d:	data_out=16'h8a00;
17'h987e:	data_out=16'h8a00;
17'h987f:	data_out=16'h9ef;
17'h9880:	data_out=16'ha00;
17'h9881:	data_out=16'ha00;
17'h9882:	data_out=16'ha00;
17'h9883:	data_out=16'h8a00;
17'h9884:	data_out=16'ha00;
17'h9885:	data_out=16'ha00;
17'h9886:	data_out=16'h8a00;
17'h9887:	data_out=16'h8a00;
17'h9888:	data_out=16'ha00;
17'h9889:	data_out=16'h8a00;
17'h988a:	data_out=16'ha00;
17'h988b:	data_out=16'h8a00;
17'h988c:	data_out=16'h81ac;
17'h988d:	data_out=16'ha00;
17'h988e:	data_out=16'ha00;
17'h988f:	data_out=16'ha00;
17'h9890:	data_out=16'h8a00;
17'h9891:	data_out=16'h9f7;
17'h9892:	data_out=16'h874e;
17'h9893:	data_out=16'h89ef;
17'h9894:	data_out=16'h8a00;
17'h9895:	data_out=16'ha00;
17'h9896:	data_out=16'ha00;
17'h9897:	data_out=16'h8a00;
17'h9898:	data_out=16'ha00;
17'h9899:	data_out=16'h8a00;
17'h989a:	data_out=16'ha00;
17'h989b:	data_out=16'h87bf;
17'h989c:	data_out=16'ha00;
17'h989d:	data_out=16'h9a5;
17'h989e:	data_out=16'h870c;
17'h989f:	data_out=16'h8a00;
17'h98a0:	data_out=16'ha00;
17'h98a1:	data_out=16'ha00;
17'h98a2:	data_out=16'h8a00;
17'h98a3:	data_out=16'ha00;
17'h98a4:	data_out=16'ha00;
17'h98a5:	data_out=16'h89b0;
17'h98a6:	data_out=16'ha00;
17'h98a7:	data_out=16'ha00;
17'h98a8:	data_out=16'ha00;
17'h98a9:	data_out=16'h8a00;
17'h98aa:	data_out=16'h96;
17'h98ab:	data_out=16'h8a00;
17'h98ac:	data_out=16'ha00;
17'h98ad:	data_out=16'h8a00;
17'h98ae:	data_out=16'h844c;
17'h98af:	data_out=16'h87c6;
17'h98b0:	data_out=16'ha00;
17'h98b1:	data_out=16'h81f2;
17'h98b2:	data_out=16'ha00;
17'h98b3:	data_out=16'h89ff;
17'h98b4:	data_out=16'h8095;
17'h98b5:	data_out=16'ha00;
17'h98b6:	data_out=16'ha00;
17'h98b7:	data_out=16'ha00;
17'h98b8:	data_out=16'h962;
17'h98b9:	data_out=16'h8550;
17'h98ba:	data_out=16'h8a00;
17'h98bb:	data_out=16'ha00;
17'h98bc:	data_out=16'h973;
17'h98bd:	data_out=16'ha00;
17'h98be:	data_out=16'ha00;
17'h98bf:	data_out=16'ha00;
17'h98c0:	data_out=16'ha00;
17'h98c1:	data_out=16'ha00;
17'h98c2:	data_out=16'h89f7;
17'h98c3:	data_out=16'h8a00;
17'h98c4:	data_out=16'ha00;
17'h98c5:	data_out=16'ha00;
17'h98c6:	data_out=16'ha00;
17'h98c7:	data_out=16'h8a00;
17'h98c8:	data_out=16'h89ff;
17'h98c9:	data_out=16'h8749;
17'h98ca:	data_out=16'h8037;
17'h98cb:	data_out=16'h89f9;
17'h98cc:	data_out=16'h8904;
17'h98cd:	data_out=16'h8a00;
17'h98ce:	data_out=16'ha00;
17'h98cf:	data_out=16'h8984;
17'h98d0:	data_out=16'h132;
17'h98d1:	data_out=16'ha00;
17'h98d2:	data_out=16'ha00;
17'h98d3:	data_out=16'h89bf;
17'h98d4:	data_out=16'ha00;
17'h98d5:	data_out=16'h3e;
17'h98d6:	data_out=16'ha00;
17'h98d7:	data_out=16'ha00;
17'h98d8:	data_out=16'ha00;
17'h98d9:	data_out=16'ha00;
17'h98da:	data_out=16'h89ff;
17'h98db:	data_out=16'ha00;
17'h98dc:	data_out=16'h3b5;
17'h98dd:	data_out=16'ha00;
17'h98de:	data_out=16'h89eb;
17'h98df:	data_out=16'ha00;
17'h98e0:	data_out=16'h8681;
17'h98e1:	data_out=16'ha00;
17'h98e2:	data_out=16'h8a00;
17'h98e3:	data_out=16'h8a00;
17'h98e4:	data_out=16'h8847;
17'h98e5:	data_out=16'h8a00;
17'h98e6:	data_out=16'h8a00;
17'h98e7:	data_out=16'h8a00;
17'h98e8:	data_out=16'ha00;
17'h98e9:	data_out=16'ha00;
17'h98ea:	data_out=16'ha00;
17'h98eb:	data_out=16'ha00;
17'h98ec:	data_out=16'ha00;
17'h98ed:	data_out=16'h8a00;
17'h98ee:	data_out=16'ha00;
17'h98ef:	data_out=16'h8a00;
17'h98f0:	data_out=16'ha00;
17'h98f1:	data_out=16'ha00;
17'h98f2:	data_out=16'ha00;
17'h98f3:	data_out=16'ha00;
17'h98f4:	data_out=16'ha00;
17'h98f5:	data_out=16'ha00;
17'h98f6:	data_out=16'h8a00;
17'h98f7:	data_out=16'h13c;
17'h98f8:	data_out=16'h8a00;
17'h98f9:	data_out=16'ha00;
17'h98fa:	data_out=16'h8a00;
17'h98fb:	data_out=16'ha00;
17'h98fc:	data_out=16'ha00;
17'h98fd:	data_out=16'h89fb;
17'h98fe:	data_out=16'h8a00;
17'h98ff:	data_out=16'ha00;
17'h9900:	data_out=16'ha00;
17'h9901:	data_out=16'ha00;
17'h9902:	data_out=16'ha00;
17'h9903:	data_out=16'h8404;
17'h9904:	data_out=16'h6bb;
17'h9905:	data_out=16'ha00;
17'h9906:	data_out=16'h88bb;
17'h9907:	data_out=16'h8a00;
17'h9908:	data_out=16'ha00;
17'h9909:	data_out=16'h8a00;
17'h990a:	data_out=16'ha00;
17'h990b:	data_out=16'h8a00;
17'h990c:	data_out=16'h8595;
17'h990d:	data_out=16'h8743;
17'h990e:	data_out=16'h7f4;
17'h990f:	data_out=16'ha00;
17'h9910:	data_out=16'h8998;
17'h9911:	data_out=16'h3e1;
17'h9912:	data_out=16'h8904;
17'h9913:	data_out=16'h86e2;
17'h9914:	data_out=16'h8113;
17'h9915:	data_out=16'ha00;
17'h9916:	data_out=16'ha00;
17'h9917:	data_out=16'h8729;
17'h9918:	data_out=16'h875;
17'h9919:	data_out=16'h8a00;
17'h991a:	data_out=16'h4be;
17'h991b:	data_out=16'h88d4;
17'h991c:	data_out=16'ha00;
17'h991d:	data_out=16'h963;
17'h991e:	data_out=16'h87;
17'h991f:	data_out=16'h35d;
17'h9920:	data_out=16'h972;
17'h9921:	data_out=16'h7b9;
17'h9922:	data_out=16'h8a00;
17'h9923:	data_out=16'h6d9;
17'h9924:	data_out=16'h6de;
17'h9925:	data_out=16'h89ee;
17'h9926:	data_out=16'h8663;
17'h9927:	data_out=16'h6d6;
17'h9928:	data_out=16'h6eb;
17'h9929:	data_out=16'h86a7;
17'h992a:	data_out=16'h8468;
17'h992b:	data_out=16'h8a00;
17'h992c:	data_out=16'h961;
17'h992d:	data_out=16'h89df;
17'h992e:	data_out=16'h3ab;
17'h992f:	data_out=16'h8341;
17'h9930:	data_out=16'ha00;
17'h9931:	data_out=16'h8041;
17'h9932:	data_out=16'h985;
17'h9933:	data_out=16'hba;
17'h9934:	data_out=16'h8028;
17'h9935:	data_out=16'ha00;
17'h9936:	data_out=16'ha00;
17'h9937:	data_out=16'ha00;
17'h9938:	data_out=16'ha00;
17'h9939:	data_out=16'h256;
17'h993a:	data_out=16'h8a00;
17'h993b:	data_out=16'ha00;
17'h993c:	data_out=16'h9fe;
17'h993d:	data_out=16'ha00;
17'h993e:	data_out=16'h6d5;
17'h993f:	data_out=16'ha00;
17'h9940:	data_out=16'h831a;
17'h9941:	data_out=16'ha00;
17'h9942:	data_out=16'h87a3;
17'h9943:	data_out=16'h8a00;
17'h9944:	data_out=16'ha00;
17'h9945:	data_out=16'ha00;
17'h9946:	data_out=16'h8093;
17'h9947:	data_out=16'h8a00;
17'h9948:	data_out=16'h89fe;
17'h9949:	data_out=16'h89bc;
17'h994a:	data_out=16'h8566;
17'h994b:	data_out=16'h8a00;
17'h994c:	data_out=16'h89e2;
17'h994d:	data_out=16'h8a00;
17'h994e:	data_out=16'h23b;
17'h994f:	data_out=16'h8a00;
17'h9950:	data_out=16'h80d1;
17'h9951:	data_out=16'ha00;
17'h9952:	data_out=16'h78b;
17'h9953:	data_out=16'h8525;
17'h9954:	data_out=16'ha00;
17'h9955:	data_out=16'h87c;
17'h9956:	data_out=16'ha00;
17'h9957:	data_out=16'h6c7;
17'h9958:	data_out=16'ha00;
17'h9959:	data_out=16'h4d2;
17'h995a:	data_out=16'h85b1;
17'h995b:	data_out=16'ha00;
17'h995c:	data_out=16'h5c4;
17'h995d:	data_out=16'ha00;
17'h995e:	data_out=16'h84ec;
17'h995f:	data_out=16'h4e7;
17'h9960:	data_out=16'h82a6;
17'h9961:	data_out=16'ha00;
17'h9962:	data_out=16'h8a00;
17'h9963:	data_out=16'h21;
17'h9964:	data_out=16'h87dd;
17'h9965:	data_out=16'h8a00;
17'h9966:	data_out=16'h8a00;
17'h9967:	data_out=16'h8a00;
17'h9968:	data_out=16'h78c;
17'h9969:	data_out=16'ha00;
17'h996a:	data_out=16'h818;
17'h996b:	data_out=16'h861;
17'h996c:	data_out=16'ha00;
17'h996d:	data_out=16'h69;
17'h996e:	data_out=16'h817;
17'h996f:	data_out=16'h87b4;
17'h9970:	data_out=16'h805;
17'h9971:	data_out=16'h90b;
17'h9972:	data_out=16'ha00;
17'h9973:	data_out=16'ha00;
17'h9974:	data_out=16'h9ff;
17'h9975:	data_out=16'ha00;
17'h9976:	data_out=16'h8a00;
17'h9977:	data_out=16'h85d2;
17'h9978:	data_out=16'h8a00;
17'h9979:	data_out=16'ha00;
17'h997a:	data_out=16'h80ac;
17'h997b:	data_out=16'h6b8;
17'h997c:	data_out=16'h72b;
17'h997d:	data_out=16'h89f8;
17'h997e:	data_out=16'h8a00;
17'h997f:	data_out=16'ha00;
17'h9980:	data_out=16'h802e;
17'h9981:	data_out=16'h99;
17'h9982:	data_out=16'h8073;
17'h9983:	data_out=16'h82cf;
17'h9984:	data_out=16'h81e5;
17'h9985:	data_out=16'h8204;
17'h9986:	data_out=16'h80ec;
17'h9987:	data_out=16'h855e;
17'h9988:	data_out=16'h81cc;
17'h9989:	data_out=16'h8602;
17'h998a:	data_out=16'h66;
17'h998b:	data_out=16'h84ad;
17'h998c:	data_out=16'h847c;
17'h998d:	data_out=16'h82ee;
17'h998e:	data_out=16'hb8;
17'h998f:	data_out=16'h80b5;
17'h9990:	data_out=16'h8430;
17'h9991:	data_out=16'h821e;
17'h9992:	data_out=16'h8213;
17'h9993:	data_out=16'h82ec;
17'h9994:	data_out=16'h8118;
17'h9995:	data_out=16'h80a4;
17'h9996:	data_out=16'h82b2;
17'h9997:	data_out=16'h80f7;
17'h9998:	data_out=16'h815e;
17'h9999:	data_out=16'h80db;
17'h999a:	data_out=16'h8203;
17'h999b:	data_out=16'h82f1;
17'h999c:	data_out=16'h8064;
17'h999d:	data_out=16'h81ee;
17'h999e:	data_out=16'h8181;
17'h999f:	data_out=16'h8420;
17'h99a0:	data_out=16'h8343;
17'h99a1:	data_out=16'ha7;
17'h99a2:	data_out=16'h82c8;
17'h99a3:	data_out=16'hd9;
17'h99a4:	data_out=16'hd8;
17'h99a5:	data_out=16'h8333;
17'h99a6:	data_out=16'h83d0;
17'h99a7:	data_out=16'h82fc;
17'h99a8:	data_out=16'h72;
17'h99a9:	data_out=16'h8108;
17'h99aa:	data_out=16'h824f;
17'h99ab:	data_out=16'h82c8;
17'h99ac:	data_out=16'h8286;
17'h99ad:	data_out=16'h75;
17'h99ae:	data_out=16'h82ca;
17'h99af:	data_out=16'h82cd;
17'h99b0:	data_out=16'h7;
17'h99b1:	data_out=16'h809a;
17'h99b2:	data_out=16'h16;
17'h99b3:	data_out=16'h8197;
17'h99b4:	data_out=16'h8023;
17'h99b5:	data_out=16'h848d;
17'h99b6:	data_out=16'h821d;
17'h99b7:	data_out=16'h807e;
17'h99b8:	data_out=16'h493;
17'h99b9:	data_out=16'h81d8;
17'h99ba:	data_out=16'h8426;
17'h99bb:	data_out=16'h82f8;
17'h99bc:	data_out=16'h4;
17'h99bd:	data_out=16'h82f4;
17'h99be:	data_out=16'h6c;
17'h99bf:	data_out=16'h8246;
17'h99c0:	data_out=16'h8267;
17'h99c1:	data_out=16'h823a;
17'h99c2:	data_out=16'h81ba;
17'h99c3:	data_out=16'h829a;
17'h99c4:	data_out=16'h82f6;
17'h99c5:	data_out=16'h81cd;
17'h99c6:	data_out=16'h20b;
17'h99c7:	data_out=16'h83d8;
17'h99c8:	data_out=16'h82fc;
17'h99c9:	data_out=16'h834b;
17'h99ca:	data_out=16'h84a2;
17'h99cb:	data_out=16'h835f;
17'h99cc:	data_out=16'h82d2;
17'h99cd:	data_out=16'h8282;
17'h99ce:	data_out=16'h8241;
17'h99cf:	data_out=16'h8335;
17'h99d0:	data_out=16'h8300;
17'h99d1:	data_out=16'h8152;
17'h99d2:	data_out=16'he6;
17'h99d3:	data_out=16'h82d4;
17'h99d4:	data_out=16'h81ce;
17'h99d5:	data_out=16'h820e;
17'h99d6:	data_out=16'h80cc;
17'h99d7:	data_out=16'h80ad;
17'h99d8:	data_out=16'h80fb;
17'h99d9:	data_out=16'h8142;
17'h99da:	data_out=16'h8098;
17'h99db:	data_out=16'h2d6;
17'h99dc:	data_out=16'h823d;
17'h99dd:	data_out=16'h8073;
17'h99de:	data_out=16'h830c;
17'h99df:	data_out=16'h8103;
17'h99e0:	data_out=16'h8150;
17'h99e1:	data_out=16'h80eb;
17'h99e2:	data_out=16'h819a;
17'h99e3:	data_out=16'h819d;
17'h99e4:	data_out=16'h82d0;
17'h99e5:	data_out=16'h84cf;
17'h99e6:	data_out=16'h82ea;
17'h99e7:	data_out=16'h8193;
17'h99e8:	data_out=16'h8a;
17'h99e9:	data_out=16'h8182;
17'h99ea:	data_out=16'hd8;
17'h99eb:	data_out=16'h82c8;
17'h99ec:	data_out=16'h180;
17'h99ed:	data_out=16'h8195;
17'h99ee:	data_out=16'hcb;
17'h99ef:	data_out=16'h8163;
17'h99f0:	data_out=16'hc6;
17'h99f1:	data_out=16'h8303;
17'h99f2:	data_out=16'hd7;
17'h99f3:	data_out=16'h80dc;
17'h99f4:	data_out=16'hd;
17'h99f5:	data_out=16'h23c;
17'h99f6:	data_out=16'h83c1;
17'h99f7:	data_out=16'h841e;
17'h99f8:	data_out=16'h823d;
17'h99f9:	data_out=16'h8335;
17'h99fa:	data_out=16'h8160;
17'h99fb:	data_out=16'h71;
17'h99fc:	data_out=16'h8084;
17'h99fd:	data_out=16'h8212;
17'h99fe:	data_out=16'h852a;
17'h99ff:	data_out=16'h835b;
17'h9a00:	data_out=16'h54;
17'h9a01:	data_out=16'h5f;
17'h9a02:	data_out=16'h22;
17'h9a03:	data_out=16'h45;
17'h9a04:	data_out=16'h6e;
17'h9a05:	data_out=16'h61;
17'h9a06:	data_out=16'h26;
17'h9a07:	data_out=16'h58;
17'h9a08:	data_out=16'h30;
17'h9a09:	data_out=16'h16;
17'h9a0a:	data_out=16'h5b;
17'h9a0b:	data_out=16'h28;
17'h9a0c:	data_out=16'h6f;
17'h9a0d:	data_out=16'h49;
17'h9a0e:	data_out=16'h19;
17'h9a0f:	data_out=16'h49;
17'h9a10:	data_out=16'h15;
17'h9a11:	data_out=16'h64;
17'h9a12:	data_out=16'h46;
17'h9a13:	data_out=16'h47;
17'h9a14:	data_out=16'h4f;
17'h9a15:	data_out=16'h42;
17'h9a16:	data_out=16'h5d;
17'h9a17:	data_out=16'h52;
17'h9a18:	data_out=16'h28;
17'h9a19:	data_out=16'h34;
17'h9a1a:	data_out=16'h6c;
17'h9a1b:	data_out=16'h3d;
17'h9a1c:	data_out=16'h5e;
17'h9a1d:	data_out=16'h5b;
17'h9a1e:	data_out=16'h2e;
17'h9a1f:	data_out=16'h30;
17'h9a20:	data_out=16'h5c;
17'h9a21:	data_out=16'hf;
17'h9a22:	data_out=16'h21;
17'h9a23:	data_out=16'h35;
17'h9a24:	data_out=16'h35;
17'h9a25:	data_out=16'h39;
17'h9a26:	data_out=16'h16;
17'h9a27:	data_out=16'h5d;
17'h9a28:	data_out=16'hf;
17'h9a29:	data_out=16'h46;
17'h9a2a:	data_out=16'h36;
17'h9a2b:	data_out=16'h3e;
17'h9a2c:	data_out=16'h4d;
17'h9a2d:	data_out=16'h30;
17'h9a2e:	data_out=16'h1e;
17'h9a2f:	data_out=16'h64;
17'h9a30:	data_out=16'h82;
17'h9a31:	data_out=16'h68;
17'h9a32:	data_out=16'h90;
17'h9a33:	data_out=16'h54;
17'h9a34:	data_out=16'h5e;
17'h9a35:	data_out=16'h7d;
17'h9a36:	data_out=16'h33;
17'h9a37:	data_out=16'h3b;
17'h9a38:	data_out=16'h5b;
17'h9a39:	data_out=16'h38;
17'h9a3a:	data_out=16'h41;
17'h9a3b:	data_out=16'h5c;
17'h9a3c:	data_out=16'h27;
17'h9a3d:	data_out=16'h50;
17'h9a3e:	data_out=16'h1e;
17'h9a3f:	data_out=16'h61;
17'h9a40:	data_out=16'h51;
17'h9a41:	data_out=16'h35;
17'h9a42:	data_out=16'h4b;
17'h9a43:	data_out=16'h21;
17'h9a44:	data_out=16'h59;
17'h9a45:	data_out=16'h34;
17'h9a46:	data_out=16'h25;
17'h9a47:	data_out=16'h3b;
17'h9a48:	data_out=16'h16;
17'h9a49:	data_out=16'h37;
17'h9a4a:	data_out=16'h74;
17'h9a4b:	data_out=16'h73;
17'h9a4c:	data_out=16'h53;
17'h9a4d:	data_out=16'h31;
17'h9a4e:	data_out=16'h5a;
17'h9a4f:	data_out=16'h5e;
17'h9a50:	data_out=16'h41;
17'h9a51:	data_out=16'h4c;
17'h9a52:	data_out=16'h34;
17'h9a53:	data_out=16'h52;
17'h9a54:	data_out=16'h65;
17'h9a55:	data_out=16'h22;
17'h9a56:	data_out=16'h52;
17'h9a57:	data_out=16'h18;
17'h9a58:	data_out=16'h22;
17'h9a59:	data_out=16'h40;
17'h9a5a:	data_out=16'h14;
17'h9a5b:	data_out=16'h4f;
17'h9a5c:	data_out=16'h49;
17'h9a5d:	data_out=16'h4d;
17'h9a5e:	data_out=16'h62;
17'h9a5f:	data_out=16'h32;
17'h9a60:	data_out=16'h36;
17'h9a61:	data_out=16'h73;
17'h9a62:	data_out=16'h27;
17'h9a63:	data_out=16'h47;
17'h9a64:	data_out=16'h51;
17'h9a65:	data_out=16'h5d;
17'h9a66:	data_out=16'h3a;
17'h9a67:	data_out=16'h25;
17'h9a68:	data_out=16'h1a;
17'h9a69:	data_out=16'h2d;
17'h9a6a:	data_out=16'h14;
17'h9a6b:	data_out=16'h6e;
17'h9a6c:	data_out=16'h5c;
17'h9a6d:	data_out=16'h46;
17'h9a6e:	data_out=16'h11;
17'h9a6f:	data_out=16'h65;
17'h9a70:	data_out=16'h19;
17'h9a71:	data_out=16'h2c;
17'h9a72:	data_out=16'h4d;
17'h9a73:	data_out=16'h63;
17'h9a74:	data_out=16'h86;
17'h9a75:	data_out=16'h48;
17'h9a76:	data_out=16'h2e;
17'h9a77:	data_out=16'h42;
17'h9a78:	data_out=16'h39;
17'h9a79:	data_out=16'h2e;
17'h9a7a:	data_out=16'h47;
17'h9a7b:	data_out=16'h1e;
17'h9a7c:	data_out=16'h1c;
17'h9a7d:	data_out=16'h3a;
17'h9a7e:	data_out=16'h12;
17'h9a7f:	data_out=16'h51;
17'h9a80:	data_out=16'h5eb;
17'h9a81:	data_out=16'h77c;
17'h9a82:	data_out=16'h164;
17'h9a83:	data_out=16'h27a;
17'h9a84:	data_out=16'h8573;
17'h9a85:	data_out=16'h8424;
17'h9a86:	data_out=16'h8678;
17'h9a87:	data_out=16'h80a4;
17'h9a88:	data_out=16'h21a;
17'h9a89:	data_out=16'h80b1;
17'h9a8a:	data_out=16'h14e;
17'h9a8b:	data_out=16'h72;
17'h9a8c:	data_out=16'h82ba;
17'h9a8d:	data_out=16'h2fa;
17'h9a8e:	data_out=16'h80f4;
17'h9a8f:	data_out=16'h25b;
17'h9a90:	data_out=16'h3cc;
17'h9a91:	data_out=16'h84f3;
17'h9a92:	data_out=16'h67f;
17'h9a93:	data_out=16'h14a;
17'h9a94:	data_out=16'h29c;
17'h9a95:	data_out=16'h80c4;
17'h9a96:	data_out=16'h800b;
17'h9a97:	data_out=16'h483;
17'h9a98:	data_out=16'h8084;
17'h9a99:	data_out=16'h8178;
17'h9a9a:	data_out=16'h8594;
17'h9a9b:	data_out=16'h78f;
17'h9a9c:	data_out=16'h843d;
17'h9a9d:	data_out=16'h570;
17'h9a9e:	data_out=16'h509;
17'h9a9f:	data_out=16'h873f;
17'h9aa0:	data_out=16'h945;
17'h9aa1:	data_out=16'h80fb;
17'h9aa2:	data_out=16'h616;
17'h9aa3:	data_out=16'h8271;
17'h9aa4:	data_out=16'h8276;
17'h9aa5:	data_out=16'h15a;
17'h9aa6:	data_out=16'h82fa;
17'h9aa7:	data_out=16'h5c1;
17'h9aa8:	data_out=16'h80ee;
17'h9aa9:	data_out=16'h486;
17'h9aaa:	data_out=16'h7d8;
17'h9aab:	data_out=16'h103;
17'h9aac:	data_out=16'h80bd;
17'h9aad:	data_out=16'h941;
17'h9aae:	data_out=16'h54b;
17'h9aaf:	data_out=16'ha00;
17'h9ab0:	data_out=16'h84c9;
17'h9ab1:	data_out=16'h1e0;
17'h9ab2:	data_out=16'h8492;
17'h9ab3:	data_out=16'h2e6;
17'h9ab4:	data_out=16'h20a;
17'h9ab5:	data_out=16'h85bb;
17'h9ab6:	data_out=16'h655;
17'h9ab7:	data_out=16'h166;
17'h9ab8:	data_out=16'h82a5;
17'h9ab9:	data_out=16'h39c;
17'h9aba:	data_out=16'h7cc;
17'h9abb:	data_out=16'h84b0;
17'h9abc:	data_out=16'h45d;
17'h9abd:	data_out=16'h8132;
17'h9abe:	data_out=16'h80ee;
17'h9abf:	data_out=16'h855b;
17'h9ac0:	data_out=16'h84a9;
17'h9ac1:	data_out=16'h1a9;
17'h9ac2:	data_out=16'h919;
17'h9ac3:	data_out=16'h8818;
17'h9ac4:	data_out=16'h843b;
17'h9ac5:	data_out=16'h8262;
17'h9ac6:	data_out=16'h345;
17'h9ac7:	data_out=16'h230;
17'h9ac8:	data_out=16'h59f;
17'h9ac9:	data_out=16'h6d;
17'h9aca:	data_out=16'h159;
17'h9acb:	data_out=16'h881;
17'h9acc:	data_out=16'h552;
17'h9acd:	data_out=16'h6b6;
17'h9ace:	data_out=16'h5ac;
17'h9acf:	data_out=16'h35c;
17'h9ad0:	data_out=16'h84df;
17'h9ad1:	data_out=16'h8514;
17'h9ad2:	data_out=16'h831e;
17'h9ad3:	data_out=16'h9e0;
17'h9ad4:	data_out=16'ha00;
17'h9ad5:	data_out=16'h80fe;
17'h9ad6:	data_out=16'h8317;
17'h9ad7:	data_out=16'h8275;
17'h9ad8:	data_out=16'h8065;
17'h9ad9:	data_out=16'h8375;
17'h9ada:	data_out=16'h695;
17'h9adb:	data_out=16'h8879;
17'h9adc:	data_out=16'h2ac;
17'h9add:	data_out=16'h81d;
17'h9ade:	data_out=16'ha00;
17'h9adf:	data_out=16'h4d6;
17'h9ae0:	data_out=16'h80ad;
17'h9ae1:	data_out=16'h8645;
17'h9ae2:	data_out=16'h1be;
17'h9ae3:	data_out=16'h2fe;
17'h9ae4:	data_out=16'h806b;
17'h9ae5:	data_out=16'h80bb;
17'h9ae6:	data_out=16'h81cc;
17'h9ae7:	data_out=16'h2e0;
17'h9ae8:	data_out=16'h80e9;
17'h9ae9:	data_out=16'h2df;
17'h9aea:	data_out=16'h80f4;
17'h9aeb:	data_out=16'h854c;
17'h9aec:	data_out=16'ha00;
17'h9aed:	data_out=16'h319;
17'h9aee:	data_out=16'h8106;
17'h9aef:	data_out=16'h80d6;
17'h9af0:	data_out=16'h80f1;
17'h9af1:	data_out=16'hee;
17'h9af2:	data_out=16'h85a9;
17'h9af3:	data_out=16'h8483;
17'h9af4:	data_out=16'h84cd;
17'h9af5:	data_out=16'h86fe;
17'h9af6:	data_out=16'h8081;
17'h9af7:	data_out=16'h84f5;
17'h9af8:	data_out=16'h87f6;
17'h9af9:	data_out=16'h56e;
17'h9afa:	data_out=16'h2f6;
17'h9afb:	data_out=16'h80ec;
17'h9afc:	data_out=16'hc6;
17'h9afd:	data_out=16'h887c;
17'h9afe:	data_out=16'h833e;
17'h9aff:	data_out=16'h84e8;
17'h9b00:	data_out=16'ha00;
17'h9b01:	data_out=16'ha00;
17'h9b02:	data_out=16'h80a;
17'h9b03:	data_out=16'h9fd;
17'h9b04:	data_out=16'h8a00;
17'h9b05:	data_out=16'h8784;
17'h9b06:	data_out=16'h89ff;
17'h9b07:	data_out=16'h803d;
17'h9b08:	data_out=16'ha00;
17'h9b09:	data_out=16'haf;
17'h9b0a:	data_out=16'h5c7;
17'h9b0b:	data_out=16'h5ea;
17'h9b0c:	data_out=16'h877b;
17'h9b0d:	data_out=16'h9ee;
17'h9b0e:	data_out=16'h81fa;
17'h9b0f:	data_out=16'ha00;
17'h9b10:	data_out=16'ha00;
17'h9b11:	data_out=16'h8a00;
17'h9b12:	data_out=16'ha00;
17'h9b13:	data_out=16'ha00;
17'h9b14:	data_out=16'h9f5;
17'h9b15:	data_out=16'h8198;
17'h9b16:	data_out=16'h217;
17'h9b17:	data_out=16'ha00;
17'h9b18:	data_out=16'hff;
17'h9b19:	data_out=16'h846e;
17'h9b1a:	data_out=16'h8a00;
17'h9b1b:	data_out=16'ha00;
17'h9b1c:	data_out=16'h86fa;
17'h9b1d:	data_out=16'ha00;
17'h9b1e:	data_out=16'ha00;
17'h9b1f:	data_out=16'h89ff;
17'h9b20:	data_out=16'ha00;
17'h9b21:	data_out=16'h81f9;
17'h9b22:	data_out=16'ha00;
17'h9b23:	data_out=16'h86da;
17'h9b24:	data_out=16'h86dd;
17'h9b25:	data_out=16'h4cf;
17'h9b26:	data_out=16'h85ff;
17'h9b27:	data_out=16'ha00;
17'h9b28:	data_out=16'h820d;
17'h9b29:	data_out=16'ha00;
17'h9b2a:	data_out=16'ha00;
17'h9b2b:	data_out=16'h6d8;
17'h9b2c:	data_out=16'h8087;
17'h9b2d:	data_out=16'ha00;
17'h9b2e:	data_out=16'ha00;
17'h9b2f:	data_out=16'ha00;
17'h9b30:	data_out=16'h8a00;
17'h9b31:	data_out=16'h696;
17'h9b32:	data_out=16'h8a00;
17'h9b33:	data_out=16'ha00;
17'h9b34:	data_out=16'h8fd;
17'h9b35:	data_out=16'h8a00;
17'h9b36:	data_out=16'ha00;
17'h9b37:	data_out=16'h7e1;
17'h9b38:	data_out=16'h80f2;
17'h9b39:	data_out=16'ha00;
17'h9b3a:	data_out=16'h9ff;
17'h9b3b:	data_out=16'h8a00;
17'h9b3c:	data_out=16'h9f0;
17'h9b3d:	data_out=16'h57f;
17'h9b3e:	data_out=16'h820e;
17'h9b3f:	data_out=16'h8791;
17'h9b40:	data_out=16'h8a00;
17'h9b41:	data_out=16'h854;
17'h9b42:	data_out=16'ha00;
17'h9b43:	data_out=16'h8a00;
17'h9b44:	data_out=16'h898f;
17'h9b45:	data_out=16'h8197;
17'h9b46:	data_out=16'ha00;
17'h9b47:	data_out=16'h8dd;
17'h9b48:	data_out=16'ha00;
17'h9b49:	data_out=16'h1f0;
17'h9b4a:	data_out=16'h706;
17'h9b4b:	data_out=16'ha00;
17'h9b4c:	data_out=16'ha00;
17'h9b4d:	data_out=16'ha00;
17'h9b4e:	data_out=16'ha00;
17'h9b4f:	data_out=16'ha00;
17'h9b50:	data_out=16'h89fe;
17'h9b51:	data_out=16'h8a00;
17'h9b52:	data_out=16'h8a00;
17'h9b53:	data_out=16'ha00;
17'h9b54:	data_out=16'ha00;
17'h9b55:	data_out=16'h817d;
17'h9b56:	data_out=16'h88e7;
17'h9b57:	data_out=16'h8727;
17'h9b58:	data_out=16'h161;
17'h9b59:	data_out=16'h8756;
17'h9b5a:	data_out=16'ha00;
17'h9b5b:	data_out=16'h8a00;
17'h9b5c:	data_out=16'h9f5;
17'h9b5d:	data_out=16'ha00;
17'h9b5e:	data_out=16'ha00;
17'h9b5f:	data_out=16'ha00;
17'h9b60:	data_out=16'h80b2;
17'h9b61:	data_out=16'h8a00;
17'h9b62:	data_out=16'h7b8;
17'h9b63:	data_out=16'ha00;
17'h9b64:	data_out=16'h8122;
17'h9b65:	data_out=16'h46b;
17'h9b66:	data_out=16'h88be;
17'h9b67:	data_out=16'h9c3;
17'h9b68:	data_out=16'h8202;
17'h9b69:	data_out=16'ha00;
17'h9b6a:	data_out=16'h8204;
17'h9b6b:	data_out=16'h89ff;
17'h9b6c:	data_out=16'ha00;
17'h9b6d:	data_out=16'ha00;
17'h9b6e:	data_out=16'h8203;
17'h9b6f:	data_out=16'h376;
17'h9b70:	data_out=16'h81ff;
17'h9b71:	data_out=16'h4e4;
17'h9b72:	data_out=16'h88ef;
17'h9b73:	data_out=16'h86db;
17'h9b74:	data_out=16'h89fe;
17'h9b75:	data_out=16'h8a00;
17'h9b76:	data_out=16'h81e2;
17'h9b77:	data_out=16'h8760;
17'h9b78:	data_out=16'h8a00;
17'h9b79:	data_out=16'ha00;
17'h9b7a:	data_out=16'ha00;
17'h9b7b:	data_out=16'h820e;
17'h9b7c:	data_out=16'h538;
17'h9b7d:	data_out=16'h8a00;
17'h9b7e:	data_out=16'h873f;
17'h9b7f:	data_out=16'h89b6;
17'h9b80:	data_out=16'h9ff;
17'h9b81:	data_out=16'ha00;
17'h9b82:	data_out=16'h9fa;
17'h9b83:	data_out=16'h8f3;
17'h9b84:	data_out=16'h8a00;
17'h9b85:	data_out=16'h856d;
17'h9b86:	data_out=16'h89e9;
17'h9b87:	data_out=16'h84c8;
17'h9b88:	data_out=16'ha00;
17'h9b89:	data_out=16'h89fb;
17'h9b8a:	data_out=16'h823f;
17'h9b8b:	data_out=16'ha00;
17'h9b8c:	data_out=16'h84cd;
17'h9b8d:	data_out=16'h8fe;
17'h9b8e:	data_out=16'h83a2;
17'h9b8f:	data_out=16'ha00;
17'h9b90:	data_out=16'h8fb;
17'h9b91:	data_out=16'h89f7;
17'h9b92:	data_out=16'ha00;
17'h9b93:	data_out=16'h910;
17'h9b94:	data_out=16'h9f8;
17'h9b95:	data_out=16'h8a00;
17'h9b96:	data_out=16'h8762;
17'h9b97:	data_out=16'ha00;
17'h9b98:	data_out=16'h13b;
17'h9b99:	data_out=16'h8323;
17'h9b9a:	data_out=16'h89fb;
17'h9b9b:	data_out=16'h9fc;
17'h9b9c:	data_out=16'h85ef;
17'h9b9d:	data_out=16'ha00;
17'h9b9e:	data_out=16'h9fd;
17'h9b9f:	data_out=16'h89ef;
17'h9ba0:	data_out=16'ha00;
17'h9ba1:	data_out=16'h8388;
17'h9ba2:	data_out=16'h9a1;
17'h9ba3:	data_out=16'h8a00;
17'h9ba4:	data_out=16'h8a00;
17'h9ba5:	data_out=16'h83d1;
17'h9ba6:	data_out=16'h8a00;
17'h9ba7:	data_out=16'ha00;
17'h9ba8:	data_out=16'h835f;
17'h9ba9:	data_out=16'h9fe;
17'h9baa:	data_out=16'ha00;
17'h9bab:	data_out=16'ha00;
17'h9bac:	data_out=16'h89ff;
17'h9bad:	data_out=16'ha00;
17'h9bae:	data_out=16'h9fc;
17'h9baf:	data_out=16'ha00;
17'h9bb0:	data_out=16'h89fe;
17'h9bb1:	data_out=16'h709;
17'h9bb2:	data_out=16'h89fd;
17'h9bb3:	data_out=16'ha00;
17'h9bb4:	data_out=16'ha00;
17'h9bb5:	data_out=16'h89fd;
17'h9bb6:	data_out=16'ha00;
17'h9bb7:	data_out=16'h9f8;
17'h9bb8:	data_out=16'ha00;
17'h9bb9:	data_out=16'ha00;
17'h9bba:	data_out=16'h8e7;
17'h9bbb:	data_out=16'h89f6;
17'h9bbc:	data_out=16'h9fd;
17'h9bbd:	data_out=16'h844d;
17'h9bbe:	data_out=16'h835e;
17'h9bbf:	data_out=16'h868b;
17'h9bc0:	data_out=16'h89fd;
17'h9bc1:	data_out=16'h9fa;
17'h9bc2:	data_out=16'h97a;
17'h9bc3:	data_out=16'h8a00;
17'h9bc4:	data_out=16'h89ef;
17'h9bc5:	data_out=16'h8a00;
17'h9bc6:	data_out=16'h9fd;
17'h9bc7:	data_out=16'h171;
17'h9bc8:	data_out=16'ha00;
17'h9bc9:	data_out=16'h8834;
17'h9bca:	data_out=16'ha00;
17'h9bcb:	data_out=16'ha00;
17'h9bcc:	data_out=16'h91d;
17'h9bcd:	data_out=16'h9fe;
17'h9bce:	data_out=16'ha00;
17'h9bcf:	data_out=16'h618;
17'h9bd0:	data_out=16'h89fc;
17'h9bd1:	data_out=16'h89fe;
17'h9bd2:	data_out=16'h8a00;
17'h9bd3:	data_out=16'ha00;
17'h9bd4:	data_out=16'ha00;
17'h9bd5:	data_out=16'h3e7;
17'h9bd6:	data_out=16'h8a00;
17'h9bd7:	data_out=16'h8a00;
17'h9bd8:	data_out=16'h84d;
17'h9bd9:	data_out=16'h89ff;
17'h9bda:	data_out=16'ha00;
17'h9bdb:	data_out=16'h89f4;
17'h9bdc:	data_out=16'ha00;
17'h9bdd:	data_out=16'ha00;
17'h9bde:	data_out=16'ha00;
17'h9bdf:	data_out=16'ha00;
17'h9be0:	data_out=16'h89ff;
17'h9be1:	data_out=16'h89fc;
17'h9be2:	data_out=16'h9f3;
17'h9be3:	data_out=16'ha00;
17'h9be4:	data_out=16'h1a8;
17'h9be5:	data_out=16'h91c;
17'h9be6:	data_out=16'h891e;
17'h9be7:	data_out=16'ha00;
17'h9be8:	data_out=16'h8384;
17'h9be9:	data_out=16'h968;
17'h9bea:	data_out=16'h83c2;
17'h9beb:	data_out=16'h89f9;
17'h9bec:	data_out=16'h9ff;
17'h9bed:	data_out=16'ha00;
17'h9bee:	data_out=16'h83c1;
17'h9bef:	data_out=16'h80aa;
17'h9bf0:	data_out=16'h83b1;
17'h9bf1:	data_out=16'ha00;
17'h9bf2:	data_out=16'h89fe;
17'h9bf3:	data_out=16'h89fd;
17'h9bf4:	data_out=16'h89f8;
17'h9bf5:	data_out=16'hac;
17'h9bf6:	data_out=16'h514;
17'h9bf7:	data_out=16'h890e;
17'h9bf8:	data_out=16'h8a00;
17'h9bf9:	data_out=16'ha00;
17'h9bfa:	data_out=16'ha00;
17'h9bfb:	data_out=16'h835c;
17'h9bfc:	data_out=16'h9c8;
17'h9bfd:	data_out=16'h89fb;
17'h9bfe:	data_out=16'h8a00;
17'h9bff:	data_out=16'h8a00;
17'h9c00:	data_out=16'h12;
17'h9c01:	data_out=16'h9fd;
17'h9c02:	data_out=16'h763;
17'h9c03:	data_out=16'h8724;
17'h9c04:	data_out=16'h89f7;
17'h9c05:	data_out=16'h89ff;
17'h9c06:	data_out=16'h89f5;
17'h9c07:	data_out=16'h89f6;
17'h9c08:	data_out=16'h84ad;
17'h9c09:	data_out=16'h89ec;
17'h9c0a:	data_out=16'h8a00;
17'h9c0b:	data_out=16'h21f;
17'h9c0c:	data_out=16'h89fd;
17'h9c0d:	data_out=16'h559;
17'h9c0e:	data_out=16'h815a;
17'h9c0f:	data_out=16'h9e6;
17'h9c10:	data_out=16'h8094;
17'h9c11:	data_out=16'h89f2;
17'h9c12:	data_out=16'ha00;
17'h9c13:	data_out=16'h84b9;
17'h9c14:	data_out=16'h77c;
17'h9c15:	data_out=16'h8a00;
17'h9c16:	data_out=16'h8a00;
17'h9c17:	data_out=16'h8b3;
17'h9c18:	data_out=16'h3e;
17'h9c19:	data_out=16'h818b;
17'h9c1a:	data_out=16'h89e1;
17'h9c1b:	data_out=16'h89e;
17'h9c1c:	data_out=16'h8767;
17'h9c1d:	data_out=16'h86fe;
17'h9c1e:	data_out=16'h915;
17'h9c1f:	data_out=16'h89fa;
17'h9c20:	data_out=16'h9fb;
17'h9c21:	data_out=16'h8112;
17'h9c22:	data_out=16'h9f9;
17'h9c23:	data_out=16'h8a00;
17'h9c24:	data_out=16'h8a00;
17'h9c25:	data_out=16'h8a00;
17'h9c26:	data_out=16'h8a00;
17'h9c27:	data_out=16'h80d5;
17'h9c28:	data_out=16'h80c2;
17'h9c29:	data_out=16'h9d0;
17'h9c2a:	data_out=16'h9e2;
17'h9c2b:	data_out=16'ha00;
17'h9c2c:	data_out=16'h8a00;
17'h9c2d:	data_out=16'ha00;
17'h9c2e:	data_out=16'h9e4;
17'h9c2f:	data_out=16'ha00;
17'h9c30:	data_out=16'h88b1;
17'h9c31:	data_out=16'h89fb;
17'h9c32:	data_out=16'h89f5;
17'h9c33:	data_out=16'h9ef;
17'h9c34:	data_out=16'h81f5;
17'h9c35:	data_out=16'h89fd;
17'h9c36:	data_out=16'h9f5;
17'h9c37:	data_out=16'h734;
17'h9c38:	data_out=16'ha00;
17'h9c39:	data_out=16'h9f2;
17'h9c3a:	data_out=16'h5f8;
17'h9c3b:	data_out=16'h8a00;
17'h9c3c:	data_out=16'h9ec;
17'h9c3d:	data_out=16'h8990;
17'h9c3e:	data_out=16'h80c1;
17'h9c3f:	data_out=16'h89ff;
17'h9c40:	data_out=16'h89fa;
17'h9c41:	data_out=16'h552;
17'h9c42:	data_out=16'h8a00;
17'h9c43:	data_out=16'h8a00;
17'h9c44:	data_out=16'h89f6;
17'h9c45:	data_out=16'h8a00;
17'h9c46:	data_out=16'h9f4;
17'h9c47:	data_out=16'h8774;
17'h9c48:	data_out=16'ha00;
17'h9c49:	data_out=16'h8a00;
17'h9c4a:	data_out=16'h711;
17'h9c4b:	data_out=16'h85;
17'h9c4c:	data_out=16'h80a8;
17'h9c4d:	data_out=16'ha00;
17'h9c4e:	data_out=16'ha00;
17'h9c4f:	data_out=16'h888a;
17'h9c50:	data_out=16'h89fc;
17'h9c51:	data_out=16'h89ff;
17'h9c52:	data_out=16'h89f9;
17'h9c53:	data_out=16'ha00;
17'h9c54:	data_out=16'ha00;
17'h9c55:	data_out=16'h49c;
17'h9c56:	data_out=16'h8a00;
17'h9c57:	data_out=16'h89ff;
17'h9c58:	data_out=16'h8aa;
17'h9c59:	data_out=16'h89f9;
17'h9c5a:	data_out=16'h9ee;
17'h9c5b:	data_out=16'h89f3;
17'h9c5c:	data_out=16'h9cd;
17'h9c5d:	data_out=16'h9fe;
17'h9c5e:	data_out=16'h9fe;
17'h9c5f:	data_out=16'ha00;
17'h9c60:	data_out=16'h8a00;
17'h9c61:	data_out=16'h8a00;
17'h9c62:	data_out=16'h86e;
17'h9c63:	data_out=16'h9f8;
17'h9c64:	data_out=16'h83f4;
17'h9c65:	data_out=16'h89f2;
17'h9c66:	data_out=16'h89f2;
17'h9c67:	data_out=16'ha00;
17'h9c68:	data_out=16'h80f5;
17'h9c69:	data_out=16'h89d7;
17'h9c6a:	data_out=16'h81a1;
17'h9c6b:	data_out=16'h89f5;
17'h9c6c:	data_out=16'h9f2;
17'h9c6d:	data_out=16'h9f6;
17'h9c6e:	data_out=16'h819f;
17'h9c6f:	data_out=16'h89fe;
17'h9c70:	data_out=16'h8177;
17'h9c71:	data_out=16'h9f4;
17'h9c72:	data_out=16'h89fb;
17'h9c73:	data_out=16'h89fa;
17'h9c74:	data_out=16'h88a8;
17'h9c75:	data_out=16'h83ff;
17'h9c76:	data_out=16'h8518;
17'h9c77:	data_out=16'h898d;
17'h9c78:	data_out=16'h89f9;
17'h9c79:	data_out=16'h939;
17'h9c7a:	data_out=16'h9a5;
17'h9c7b:	data_out=16'h80c0;
17'h9c7c:	data_out=16'h9b5;
17'h9c7d:	data_out=16'h89ef;
17'h9c7e:	data_out=16'h89fe;
17'h9c7f:	data_out=16'h89a8;
17'h9c80:	data_out=16'h86ee;
17'h9c81:	data_out=16'h89c9;
17'h9c82:	data_out=16'h89ff;
17'h9c83:	data_out=16'h8a00;
17'h9c84:	data_out=16'h8985;
17'h9c85:	data_out=16'h8a00;
17'h9c86:	data_out=16'h89f8;
17'h9c87:	data_out=16'h89fa;
17'h9c88:	data_out=16'h826a;
17'h9c89:	data_out=16'h89d7;
17'h9c8a:	data_out=16'h89db;
17'h9c8b:	data_out=16'h88b9;
17'h9c8c:	data_out=16'h857b;
17'h9c8d:	data_out=16'h89fe;
17'h9c8e:	data_out=16'h78a;
17'h9c8f:	data_out=16'h89fc;
17'h9c90:	data_out=16'h595;
17'h9c91:	data_out=16'h89f5;
17'h9c92:	data_out=16'h82bf;
17'h9c93:	data_out=16'h89fe;
17'h9c94:	data_out=16'h8a00;
17'h9c95:	data_out=16'h8a00;
17'h9c96:	data_out=16'h89ff;
17'h9c97:	data_out=16'h8a00;
17'h9c98:	data_out=16'h88e2;
17'h9c99:	data_out=16'ha00;
17'h9c9a:	data_out=16'h89fe;
17'h9c9b:	data_out=16'h8a00;
17'h9c9c:	data_out=16'h8a00;
17'h9c9d:	data_out=16'h89fd;
17'h9c9e:	data_out=16'h89ff;
17'h9c9f:	data_out=16'h89ff;
17'h9ca0:	data_out=16'h89fb;
17'h9ca1:	data_out=16'h7c7;
17'h9ca2:	data_out=16'h9ff;
17'h9ca3:	data_out=16'ha00;
17'h9ca4:	data_out=16'ha00;
17'h9ca5:	data_out=16'h89f7;
17'h9ca6:	data_out=16'h8652;
17'h9ca7:	data_out=16'h89fe;
17'h9ca8:	data_out=16'h7cb;
17'h9ca9:	data_out=16'h39;
17'h9caa:	data_out=16'h89fd;
17'h9cab:	data_out=16'ha00;
17'h9cac:	data_out=16'h8a00;
17'h9cad:	data_out=16'h9fc;
17'h9cae:	data_out=16'h8377;
17'h9caf:	data_out=16'h89fe;
17'h9cb0:	data_out=16'h85d3;
17'h9cb1:	data_out=16'h8a00;
17'h9cb2:	data_out=16'h89fd;
17'h9cb3:	data_out=16'h89ff;
17'h9cb4:	data_out=16'h889c;
17'h9cb5:	data_out=16'h89ff;
17'h9cb6:	data_out=16'h8892;
17'h9cb7:	data_out=16'h8a00;
17'h9cb8:	data_out=16'h723;
17'h9cb9:	data_out=16'h89ff;
17'h9cba:	data_out=16'hb5;
17'h9cbb:	data_out=16'h8a00;
17'h9cbc:	data_out=16'h837e;
17'h9cbd:	data_out=16'h89fb;
17'h9cbe:	data_out=16'h7c9;
17'h9cbf:	data_out=16'h8a00;
17'h9cc0:	data_out=16'h89fb;
17'h9cc1:	data_out=16'h8a00;
17'h9cc2:	data_out=16'h9e8;
17'h9cc3:	data_out=16'h8a00;
17'h9cc4:	data_out=16'h89ff;
17'h9cc5:	data_out=16'h8a00;
17'h9cc6:	data_out=16'h9f1;
17'h9cc7:	data_out=16'h84e0;
17'h9cc8:	data_out=16'h309;
17'h9cc9:	data_out=16'h89fc;
17'h9cca:	data_out=16'h85f0;
17'h9ccb:	data_out=16'h9c7;
17'h9ccc:	data_out=16'ha00;
17'h9ccd:	data_out=16'ha00;
17'h9cce:	data_out=16'h837e;
17'h9ccf:	data_out=16'h8274;
17'h9cd0:	data_out=16'h8a00;
17'h9cd1:	data_out=16'h8a00;
17'h9cd2:	data_out=16'h9f6;
17'h9cd3:	data_out=16'h89fd;
17'h9cd4:	data_out=16'h863f;
17'h9cd5:	data_out=16'h8366;
17'h9cd6:	data_out=16'h8a00;
17'h9cd7:	data_out=16'h891f;
17'h9cd8:	data_out=16'h3e1;
17'h9cd9:	data_out=16'h89e8;
17'h9cda:	data_out=16'h878c;
17'h9cdb:	data_out=16'h89ff;
17'h9cdc:	data_out=16'h8a00;
17'h9cdd:	data_out=16'h88aa;
17'h9cde:	data_out=16'h8a00;
17'h9cdf:	data_out=16'h559;
17'h9ce0:	data_out=16'h7e3;
17'h9ce1:	data_out=16'h8a00;
17'h9ce2:	data_out=16'h8a00;
17'h9ce3:	data_out=16'h89ff;
17'h9ce4:	data_out=16'h8347;
17'h9ce5:	data_out=16'h8a00;
17'h9ce6:	data_out=16'h8717;
17'h9ce7:	data_out=16'ha00;
17'h9ce8:	data_out=16'h7dc;
17'h9ce9:	data_out=16'hdf;
17'h9cea:	data_out=16'h756;
17'h9ceb:	data_out=16'h8a00;
17'h9cec:	data_out=16'h84ce;
17'h9ced:	data_out=16'h89ff;
17'h9cee:	data_out=16'h759;
17'h9cef:	data_out=16'h8a00;
17'h9cf0:	data_out=16'h77a;
17'h9cf1:	data_out=16'h89fb;
17'h9cf2:	data_out=16'h8a00;
17'h9cf3:	data_out=16'h89fa;
17'h9cf4:	data_out=16'h85c7;
17'h9cf5:	data_out=16'h8a00;
17'h9cf6:	data_out=16'h586;
17'h9cf7:	data_out=16'h873b;
17'h9cf8:	data_out=16'h8029;
17'h9cf9:	data_out=16'h8841;
17'h9cfa:	data_out=16'h8a00;
17'h9cfb:	data_out=16'h7ca;
17'h9cfc:	data_out=16'h87c8;
17'h9cfd:	data_out=16'h89fd;
17'h9cfe:	data_out=16'h89f9;
17'h9cff:	data_out=16'h89fe;
17'h9d00:	data_out=16'h869d;
17'h9d01:	data_out=16'h89f7;
17'h9d02:	data_out=16'h539;
17'h9d03:	data_out=16'h89f8;
17'h9d04:	data_out=16'h87ea;
17'h9d05:	data_out=16'h89ff;
17'h9d06:	data_out=16'h89ff;
17'h9d07:	data_out=16'h8f6;
17'h9d08:	data_out=16'h861f;
17'h9d09:	data_out=16'h875e;
17'h9d0a:	data_out=16'h869e;
17'h9d0b:	data_out=16'h877a;
17'h9d0c:	data_out=16'h9cd;
17'h9d0d:	data_out=16'h89f5;
17'h9d0e:	data_out=16'h9f8;
17'h9d0f:	data_out=16'h85c2;
17'h9d10:	data_out=16'h89fa;
17'h9d11:	data_out=16'h89f8;
17'h9d12:	data_out=16'h89a7;
17'h9d13:	data_out=16'h8223;
17'h9d14:	data_out=16'h89ff;
17'h9d15:	data_out=16'h89f9;
17'h9d16:	data_out=16'h89f7;
17'h9d17:	data_out=16'h89fe;
17'h9d18:	data_out=16'h874e;
17'h9d19:	data_out=16'ha00;
17'h9d1a:	data_out=16'h89ef;
17'h9d1b:	data_out=16'h89fb;
17'h9d1c:	data_out=16'h8a00;
17'h9d1d:	data_out=16'h8a00;
17'h9d1e:	data_out=16'h89fe;
17'h9d1f:	data_out=16'h8a00;
17'h9d20:	data_out=16'h89f2;
17'h9d21:	data_out=16'h9f6;
17'h9d22:	data_out=16'h9fc;
17'h9d23:	data_out=16'ha00;
17'h9d24:	data_out=16'ha00;
17'h9d25:	data_out=16'h33f;
17'h9d26:	data_out=16'h9ff;
17'h9d27:	data_out=16'h89f6;
17'h9d28:	data_out=16'h9e2;
17'h9d29:	data_out=16'h921;
17'h9d2a:	data_out=16'h8417;
17'h9d2b:	data_out=16'ha00;
17'h9d2c:	data_out=16'h89fa;
17'h9d2d:	data_out=16'h9f9;
17'h9d2e:	data_out=16'h89fe;
17'h9d2f:	data_out=16'h89fc;
17'h9d30:	data_out=16'h386;
17'h9d31:	data_out=16'h8a00;
17'h9d32:	data_out=16'h86ec;
17'h9d33:	data_out=16'h8a00;
17'h9d34:	data_out=16'h89e7;
17'h9d35:	data_out=16'h89f2;
17'h9d36:	data_out=16'h89cc;
17'h9d37:	data_out=16'h353;
17'h9d38:	data_out=16'h8a00;
17'h9d39:	data_out=16'h89ff;
17'h9d3a:	data_out=16'h876b;
17'h9d3b:	data_out=16'h89e9;
17'h9d3c:	data_out=16'h8266;
17'h9d3d:	data_out=16'h89df;
17'h9d3e:	data_out=16'h9e1;
17'h9d3f:	data_out=16'h89ff;
17'h9d40:	data_out=16'h8936;
17'h9d41:	data_out=16'h89fb;
17'h9d42:	data_out=16'h9f4;
17'h9d43:	data_out=16'h8a00;
17'h9d44:	data_out=16'h89fe;
17'h9d45:	data_out=16'h89f9;
17'h9d46:	data_out=16'h9fd;
17'h9d47:	data_out=16'ha00;
17'h9d48:	data_out=16'h89f1;
17'h9d49:	data_out=16'h80b7;
17'h9d4a:	data_out=16'h889e;
17'h9d4b:	data_out=16'h9d0;
17'h9d4c:	data_out=16'ha00;
17'h9d4d:	data_out=16'h9fe;
17'h9d4e:	data_out=16'h4cd;
17'h9d4f:	data_out=16'ha00;
17'h9d50:	data_out=16'h89ff;
17'h9d51:	data_out=16'h8627;
17'h9d52:	data_out=16'ha00;
17'h9d53:	data_out=16'h89fd;
17'h9d54:	data_out=16'h89f1;
17'h9d55:	data_out=16'h33;
17'h9d56:	data_out=16'h5a2;
17'h9d57:	data_out=16'h44a;
17'h9d58:	data_out=16'h370;
17'h9d59:	data_out=16'h89b9;
17'h9d5a:	data_out=16'h89fe;
17'h9d5b:	data_out=16'h89f9;
17'h9d5c:	data_out=16'h8a00;
17'h9d5d:	data_out=16'h89dd;
17'h9d5e:	data_out=16'h89fe;
17'h9d5f:	data_out=16'h894c;
17'h9d60:	data_out=16'ha00;
17'h9d61:	data_out=16'h89e2;
17'h9d62:	data_out=16'h89ff;
17'h9d63:	data_out=16'h89ff;
17'h9d64:	data_out=16'h87eb;
17'h9d65:	data_out=16'h89fb;
17'h9d66:	data_out=16'h254;
17'h9d67:	data_out=16'h613;
17'h9d68:	data_out=16'h9f3;
17'h9d69:	data_out=16'h74c;
17'h9d6a:	data_out=16'h9f2;
17'h9d6b:	data_out=16'h89ff;
17'h9d6c:	data_out=16'h8330;
17'h9d6d:	data_out=16'h89ff;
17'h9d6e:	data_out=16'h9f2;
17'h9d6f:	data_out=16'h89ef;
17'h9d70:	data_out=16'h9f6;
17'h9d71:	data_out=16'h892c;
17'h9d72:	data_out=16'h89ef;
17'h9d73:	data_out=16'h89de;
17'h9d74:	data_out=16'h5eb;
17'h9d75:	data_out=16'h8a00;
17'h9d76:	data_out=16'ha00;
17'h9d77:	data_out=16'h8146;
17'h9d78:	data_out=16'h852f;
17'h9d79:	data_out=16'h3b4;
17'h9d7a:	data_out=16'h89ff;
17'h9d7b:	data_out=16'h9e1;
17'h9d7c:	data_out=16'h89f8;
17'h9d7d:	data_out=16'h8a00;
17'h9d7e:	data_out=16'h89fa;
17'h9d7f:	data_out=16'h8a00;
17'h9d80:	data_out=16'h88b1;
17'h9d81:	data_out=16'h89fd;
17'h9d82:	data_out=16'h9f0;
17'h9d83:	data_out=16'h84dc;
17'h9d84:	data_out=16'h89f5;
17'h9d85:	data_out=16'h8a00;
17'h9d86:	data_out=16'h8a00;
17'h9d87:	data_out=16'h9fe;
17'h9d88:	data_out=16'h890d;
17'h9d89:	data_out=16'h854c;
17'h9d8a:	data_out=16'h84f4;
17'h9d8b:	data_out=16'h85f6;
17'h9d8c:	data_out=16'ha00;
17'h9d8d:	data_out=16'h85ae;
17'h9d8e:	data_out=16'h9fe;
17'h9d8f:	data_out=16'h9fd;
17'h9d90:	data_out=16'h89eb;
17'h9d91:	data_out=16'h8a00;
17'h9d92:	data_out=16'h896b;
17'h9d93:	data_out=16'ha00;
17'h9d94:	data_out=16'h89ef;
17'h9d95:	data_out=16'h89fe;
17'h9d96:	data_out=16'h89ee;
17'h9d97:	data_out=16'h89d9;
17'h9d98:	data_out=16'h89fe;
17'h9d99:	data_out=16'ha00;
17'h9d9a:	data_out=16'h8a00;
17'h9d9b:	data_out=16'h8916;
17'h9d9c:	data_out=16'h89f4;
17'h9d9d:	data_out=16'h8a00;
17'h9d9e:	data_out=16'h89de;
17'h9d9f:	data_out=16'h8a00;
17'h9da0:	data_out=16'h89ff;
17'h9da1:	data_out=16'h9fe;
17'h9da2:	data_out=16'ha00;
17'h9da3:	data_out=16'h9ff;
17'h9da4:	data_out=16'h9ff;
17'h9da5:	data_out=16'h9ff;
17'h9da6:	data_out=16'ha00;
17'h9da7:	data_out=16'h89fc;
17'h9da8:	data_out=16'h9f5;
17'h9da9:	data_out=16'h9f9;
17'h9daa:	data_out=16'ha00;
17'h9dab:	data_out=16'h84fb;
17'h9dac:	data_out=16'h89f9;
17'h9dad:	data_out=16'ha00;
17'h9dae:	data_out=16'h866d;
17'h9daf:	data_out=16'h89f4;
17'h9db0:	data_out=16'ha00;
17'h9db1:	data_out=16'h8a00;
17'h9db2:	data_out=16'h81e6;
17'h9db3:	data_out=16'h89fc;
17'h9db4:	data_out=16'h89fc;
17'h9db5:	data_out=16'h89f5;
17'h9db6:	data_out=16'h8923;
17'h9db7:	data_out=16'h9d0;
17'h9db8:	data_out=16'h8a00;
17'h9db9:	data_out=16'h89fc;
17'h9dba:	data_out=16'h86a1;
17'h9dbb:	data_out=16'h89fe;
17'h9dbc:	data_out=16'h9f6;
17'h9dbd:	data_out=16'h89f8;
17'h9dbe:	data_out=16'h9f4;
17'h9dbf:	data_out=16'h8a00;
17'h9dc0:	data_out=16'h89d0;
17'h9dc1:	data_out=16'h89bb;
17'h9dc2:	data_out=16'ha00;
17'h9dc3:	data_out=16'h89ff;
17'h9dc4:	data_out=16'h8a00;
17'h9dc5:	data_out=16'h89fe;
17'h9dc6:	data_out=16'ha00;
17'h9dc7:	data_out=16'ha00;
17'h9dc8:	data_out=16'h89fa;
17'h9dc9:	data_out=16'ha00;
17'h9dca:	data_out=16'h89f8;
17'h9dcb:	data_out=16'h9fa;
17'h9dcc:	data_out=16'ha00;
17'h9dcd:	data_out=16'h9f8;
17'h9dce:	data_out=16'ha00;
17'h9dcf:	data_out=16'ha00;
17'h9dd0:	data_out=16'h89fb;
17'h9dd1:	data_out=16'h82f6;
17'h9dd2:	data_out=16'ha00;
17'h9dd3:	data_out=16'h89fc;
17'h9dd4:	data_out=16'h89f3;
17'h9dd5:	data_out=16'h5e4;
17'h9dd6:	data_out=16'h9b9;
17'h9dd7:	data_out=16'h2d8;
17'h9dd8:	data_out=16'h2d4;
17'h9dd9:	data_out=16'h89cb;
17'h9dda:	data_out=16'h89f5;
17'h9ddb:	data_out=16'h8a00;
17'h9ddc:	data_out=16'h8a00;
17'h9ddd:	data_out=16'h8971;
17'h9dde:	data_out=16'h89f6;
17'h9ddf:	data_out=16'h89d2;
17'h9de0:	data_out=16'ha00;
17'h9de1:	data_out=16'h89fd;
17'h9de2:	data_out=16'h85f1;
17'h9de3:	data_out=16'h89fc;
17'h9de4:	data_out=16'h8966;
17'h9de5:	data_out=16'h8a00;
17'h9de6:	data_out=16'h38f;
17'h9de7:	data_out=16'ha00;
17'h9de8:	data_out=16'h9fc;
17'h9de9:	data_out=16'h784;
17'h9dea:	data_out=16'h9fe;
17'h9deb:	data_out=16'h8a00;
17'h9dec:	data_out=16'h8181;
17'h9ded:	data_out=16'h89fc;
17'h9dee:	data_out=16'h9fe;
17'h9def:	data_out=16'h89f8;
17'h9df0:	data_out=16'h9fe;
17'h9df1:	data_out=16'h8816;
17'h9df2:	data_out=16'h89ff;
17'h9df3:	data_out=16'h89f1;
17'h9df4:	data_out=16'ha00;
17'h9df5:	data_out=16'h8a00;
17'h9df6:	data_out=16'h9f6;
17'h9df7:	data_out=16'h47e;
17'h9df8:	data_out=16'h45a;
17'h9df9:	data_out=16'h9f0;
17'h9dfa:	data_out=16'h89f9;
17'h9dfb:	data_out=16'h9f4;
17'h9dfc:	data_out=16'h8a00;
17'h9dfd:	data_out=16'h8a00;
17'h9dfe:	data_out=16'h89ce;
17'h9dff:	data_out=16'h8a00;
17'h9e00:	data_out=16'h8808;
17'h9e01:	data_out=16'h89fc;
17'h9e02:	data_out=16'ha00;
17'h9e03:	data_out=16'h49f;
17'h9e04:	data_out=16'h89ff;
17'h9e05:	data_out=16'h8a00;
17'h9e06:	data_out=16'h8a00;
17'h9e07:	data_out=16'h9f4;
17'h9e08:	data_out=16'h881a;
17'h9e09:	data_out=16'h7c1;
17'h9e0a:	data_out=16'h840c;
17'h9e0b:	data_out=16'h8806;
17'h9e0c:	data_out=16'ha00;
17'h9e0d:	data_out=16'h9f2;
17'h9e0e:	data_out=16'ha00;
17'h9e0f:	data_out=16'ha00;
17'h9e10:	data_out=16'h89cd;
17'h9e11:	data_out=16'h8a00;
17'h9e12:	data_out=16'h86a1;
17'h9e13:	data_out=16'ha00;
17'h9e14:	data_out=16'h89ed;
17'h9e15:	data_out=16'h89f1;
17'h9e16:	data_out=16'h8955;
17'h9e17:	data_out=16'h8943;
17'h9e18:	data_out=16'h89fa;
17'h9e19:	data_out=16'h9f9;
17'h9e1a:	data_out=16'h8a00;
17'h9e1b:	data_out=16'h850b;
17'h9e1c:	data_out=16'h89a6;
17'h9e1d:	data_out=16'h8a00;
17'h9e1e:	data_out=16'h8786;
17'h9e1f:	data_out=16'h8a00;
17'h9e20:	data_out=16'h8a00;
17'h9e21:	data_out=16'ha00;
17'h9e22:	data_out=16'ha00;
17'h9e23:	data_out=16'ha00;
17'h9e24:	data_out=16'ha00;
17'h9e25:	data_out=16'ha00;
17'h9e26:	data_out=16'ha00;
17'h9e27:	data_out=16'h8a00;
17'h9e28:	data_out=16'ha00;
17'h9e29:	data_out=16'ha00;
17'h9e2a:	data_out=16'ha00;
17'h9e2b:	data_out=16'h89d6;
17'h9e2c:	data_out=16'h89d2;
17'h9e2d:	data_out=16'ha00;
17'h9e2e:	data_out=16'h895e;
17'h9e2f:	data_out=16'h89f3;
17'h9e30:	data_out=16'ha00;
17'h9e31:	data_out=16'h8a00;
17'h9e32:	data_out=16'h82e1;
17'h9e33:	data_out=16'h89f9;
17'h9e34:	data_out=16'h89db;
17'h9e35:	data_out=16'h89ec;
17'h9e36:	data_out=16'h8724;
17'h9e37:	data_out=16'ha00;
17'h9e38:	data_out=16'h8a00;
17'h9e39:	data_out=16'h89f8;
17'h9e3a:	data_out=16'h8332;
17'h9e3b:	data_out=16'h8a00;
17'h9e3c:	data_out=16'ha00;
17'h9e3d:	data_out=16'h89cc;
17'h9e3e:	data_out=16'ha00;
17'h9e3f:	data_out=16'h8a00;
17'h9e40:	data_out=16'h89bc;
17'h9e41:	data_out=16'h881a;
17'h9e42:	data_out=16'ha00;
17'h9e43:	data_out=16'h89f8;
17'h9e44:	data_out=16'h8a00;
17'h9e45:	data_out=16'h89ef;
17'h9e46:	data_out=16'ha00;
17'h9e47:	data_out=16'ha00;
17'h9e48:	data_out=16'h89e9;
17'h9e49:	data_out=16'ha00;
17'h9e4a:	data_out=16'h8a00;
17'h9e4b:	data_out=16'ha00;
17'h9e4c:	data_out=16'ha00;
17'h9e4d:	data_out=16'ha00;
17'h9e4e:	data_out=16'ha00;
17'h9e4f:	data_out=16'ha00;
17'h9e50:	data_out=16'h89f8;
17'h9e51:	data_out=16'h9e3;
17'h9e52:	data_out=16'ha00;
17'h9e53:	data_out=16'h8a00;
17'h9e54:	data_out=16'h89f2;
17'h9e55:	data_out=16'ha00;
17'h9e56:	data_out=16'ha00;
17'h9e57:	data_out=16'h9ee;
17'h9e58:	data_out=16'h9d4;
17'h9e59:	data_out=16'h899d;
17'h9e5a:	data_out=16'h89f5;
17'h9e5b:	data_out=16'h8a00;
17'h9e5c:	data_out=16'h8a00;
17'h9e5d:	data_out=16'h8880;
17'h9e5e:	data_out=16'h89eb;
17'h9e5f:	data_out=16'h89d3;
17'h9e60:	data_out=16'ha00;
17'h9e61:	data_out=16'h89fc;
17'h9e62:	data_out=16'h867c;
17'h9e63:	data_out=16'h89fb;
17'h9e64:	data_out=16'h89ed;
17'h9e65:	data_out=16'h8a00;
17'h9e66:	data_out=16'h812c;
17'h9e67:	data_out=16'ha00;
17'h9e68:	data_out=16'ha00;
17'h9e69:	data_out=16'ha00;
17'h9e6a:	data_out=16'ha00;
17'h9e6b:	data_out=16'h8a00;
17'h9e6c:	data_out=16'h8380;
17'h9e6d:	data_out=16'h89fa;
17'h9e6e:	data_out=16'ha00;
17'h9e6f:	data_out=16'h89fe;
17'h9e70:	data_out=16'ha00;
17'h9e71:	data_out=16'h8499;
17'h9e72:	data_out=16'h89d4;
17'h9e73:	data_out=16'h89e4;
17'h9e74:	data_out=16'ha00;
17'h9e75:	data_out=16'h8a00;
17'h9e76:	data_out=16'h9f6;
17'h9e77:	data_out=16'ha00;
17'h9e78:	data_out=16'h868c;
17'h9e79:	data_out=16'h9f3;
17'h9e7a:	data_out=16'h89f4;
17'h9e7b:	data_out=16'ha00;
17'h9e7c:	data_out=16'h8a00;
17'h9e7d:	data_out=16'h8a00;
17'h9e7e:	data_out=16'h89ae;
17'h9e7f:	data_out=16'h8a00;
17'h9e80:	data_out=16'h8887;
17'h9e81:	data_out=16'h89f9;
17'h9e82:	data_out=16'ha00;
17'h9e83:	data_out=16'ha00;
17'h9e84:	data_out=16'h8a00;
17'h9e85:	data_out=16'h8a00;
17'h9e86:	data_out=16'h8a00;
17'h9e87:	data_out=16'h9ff;
17'h9e88:	data_out=16'h2c8;
17'h9e89:	data_out=16'ha00;
17'h9e8a:	data_out=16'h9ea;
17'h9e8b:	data_out=16'h89bf;
17'h9e8c:	data_out=16'h9ff;
17'h9e8d:	data_out=16'ha00;
17'h9e8e:	data_out=16'ha00;
17'h9e8f:	data_out=16'ha00;
17'h9e90:	data_out=16'h89ad;
17'h9e91:	data_out=16'h8a00;
17'h9e92:	data_out=16'h849b;
17'h9e93:	data_out=16'h303;
17'h9e94:	data_out=16'h89d7;
17'h9e95:	data_out=16'h89e9;
17'h9e96:	data_out=16'h87f7;
17'h9e97:	data_out=16'h89c1;
17'h9e98:	data_out=16'h95c;
17'h9e99:	data_out=16'h8973;
17'h9e9a:	data_out=16'h8a00;
17'h9e9b:	data_out=16'h85;
17'h9e9c:	data_out=16'h899c;
17'h9e9d:	data_out=16'h8a00;
17'h9e9e:	data_out=16'h8481;
17'h9e9f:	data_out=16'h8a00;
17'h9ea0:	data_out=16'h8a00;
17'h9ea1:	data_out=16'ha00;
17'h9ea2:	data_out=16'ha00;
17'h9ea3:	data_out=16'ha00;
17'h9ea4:	data_out=16'ha00;
17'h9ea5:	data_out=16'ha00;
17'h9ea6:	data_out=16'ha00;
17'h9ea7:	data_out=16'h8a00;
17'h9ea8:	data_out=16'ha00;
17'h9ea9:	data_out=16'ha00;
17'h9eaa:	data_out=16'ha00;
17'h9eab:	data_out=16'h89ff;
17'h9eac:	data_out=16'h89ac;
17'h9ead:	data_out=16'ha00;
17'h9eae:	data_out=16'h8483;
17'h9eaf:	data_out=16'h89ea;
17'h9eb0:	data_out=16'ha00;
17'h9eb1:	data_out=16'h8a00;
17'h9eb2:	data_out=16'h820a;
17'h9eb3:	data_out=16'h89f9;
17'h9eb4:	data_out=16'h89d6;
17'h9eb5:	data_out=16'h89df;
17'h9eb6:	data_out=16'h83f7;
17'h9eb7:	data_out=16'ha00;
17'h9eb8:	data_out=16'h8a00;
17'h9eb9:	data_out=16'h89f6;
17'h9eba:	data_out=16'ha00;
17'h9ebb:	data_out=16'h8a00;
17'h9ebc:	data_out=16'h4f6;
17'h9ebd:	data_out=16'h89b3;
17'h9ebe:	data_out=16'ha00;
17'h9ebf:	data_out=16'h8a00;
17'h9ec0:	data_out=16'h89b7;
17'h9ec1:	data_out=16'h853;
17'h9ec2:	data_out=16'ha00;
17'h9ec3:	data_out=16'h8a00;
17'h9ec4:	data_out=16'h8a00;
17'h9ec5:	data_out=16'h89e7;
17'h9ec6:	data_out=16'ha00;
17'h9ec7:	data_out=16'h9fe;
17'h9ec8:	data_out=16'h89b3;
17'h9ec9:	data_out=16'ha00;
17'h9eca:	data_out=16'h89ff;
17'h9ecb:	data_out=16'ha00;
17'h9ecc:	data_out=16'ha00;
17'h9ecd:	data_out=16'h9ff;
17'h9ece:	data_out=16'h9ff;
17'h9ecf:	data_out=16'ha00;
17'h9ed0:	data_out=16'h89f8;
17'h9ed1:	data_out=16'h9ff;
17'h9ed2:	data_out=16'ha00;
17'h9ed3:	data_out=16'h89ff;
17'h9ed4:	data_out=16'h89da;
17'h9ed5:	data_out=16'ha00;
17'h9ed6:	data_out=16'ha00;
17'h9ed7:	data_out=16'h9ff;
17'h9ed8:	data_out=16'h9da;
17'h9ed9:	data_out=16'h86b3;
17'h9eda:	data_out=16'h89e2;
17'h9edb:	data_out=16'h8a00;
17'h9edc:	data_out=16'h8a00;
17'h9edd:	data_out=16'h85ab;
17'h9ede:	data_out=16'h89ad;
17'h9edf:	data_out=16'h89dc;
17'h9ee0:	data_out=16'ha00;
17'h9ee1:	data_out=16'h89f1;
17'h9ee2:	data_out=16'h8754;
17'h9ee3:	data_out=16'h89ff;
17'h9ee4:	data_out=16'h89ff;
17'h9ee5:	data_out=16'h8a00;
17'h9ee6:	data_out=16'h89de;
17'h9ee7:	data_out=16'ha00;
17'h9ee8:	data_out=16'ha00;
17'h9ee9:	data_out=16'ha00;
17'h9eea:	data_out=16'ha00;
17'h9eeb:	data_out=16'h8a00;
17'h9eec:	data_out=16'h9ef;
17'h9eed:	data_out=16'h89fe;
17'h9eee:	data_out=16'ha00;
17'h9eef:	data_out=16'h89fe;
17'h9ef0:	data_out=16'ha00;
17'h9ef1:	data_out=16'h327;
17'h9ef2:	data_out=16'h89d1;
17'h9ef3:	data_out=16'h89af;
17'h9ef4:	data_out=16'ha00;
17'h9ef5:	data_out=16'h8a00;
17'h9ef6:	data_out=16'h9e9;
17'h9ef7:	data_out=16'ha00;
17'h9ef8:	data_out=16'h8a00;
17'h9ef9:	data_out=16'ha00;
17'h9efa:	data_out=16'h89e8;
17'h9efb:	data_out=16'ha00;
17'h9efc:	data_out=16'h8a00;
17'h9efd:	data_out=16'h8a00;
17'h9efe:	data_out=16'h89df;
17'h9eff:	data_out=16'h8a00;
17'h9f00:	data_out=16'h97f;
17'h9f01:	data_out=16'h89cd;
17'h9f02:	data_out=16'ha00;
17'h9f03:	data_out=16'ha00;
17'h9f04:	data_out=16'h8a00;
17'h9f05:	data_out=16'h8a00;
17'h9f06:	data_out=16'h8a00;
17'h9f07:	data_out=16'ha00;
17'h9f08:	data_out=16'h95c;
17'h9f09:	data_out=16'ha00;
17'h9f0a:	data_out=16'h9ee;
17'h9f0b:	data_out=16'h89fd;
17'h9f0c:	data_out=16'h9c5;
17'h9f0d:	data_out=16'ha00;
17'h9f0e:	data_out=16'ha00;
17'h9f0f:	data_out=16'ha00;
17'h9f10:	data_out=16'h89e8;
17'h9f11:	data_out=16'h8a00;
17'h9f12:	data_out=16'hf9;
17'h9f13:	data_out=16'h47a;
17'h9f14:	data_out=16'h89e5;
17'h9f15:	data_out=16'h9cb;
17'h9f16:	data_out=16'h9f6;
17'h9f17:	data_out=16'h88e8;
17'h9f18:	data_out=16'h999;
17'h9f19:	data_out=16'h8a00;
17'h9f1a:	data_out=16'h8a00;
17'h9f1b:	data_out=16'ha00;
17'h9f1c:	data_out=16'h8884;
17'h9f1d:	data_out=16'h8a00;
17'h9f1e:	data_out=16'h4c6;
17'h9f1f:	data_out=16'h8a00;
17'h9f20:	data_out=16'h8a00;
17'h9f21:	data_out=16'ha00;
17'h9f22:	data_out=16'h9fb;
17'h9f23:	data_out=16'ha00;
17'h9f24:	data_out=16'ha00;
17'h9f25:	data_out=16'ha00;
17'h9f26:	data_out=16'ha00;
17'h9f27:	data_out=16'h8a00;
17'h9f28:	data_out=16'ha00;
17'h9f29:	data_out=16'ha00;
17'h9f2a:	data_out=16'h9f5;
17'h9f2b:	data_out=16'h8a00;
17'h9f2c:	data_out=16'h9cd;
17'h9f2d:	data_out=16'h89ca;
17'h9f2e:	data_out=16'h97e;
17'h9f2f:	data_out=16'h89d7;
17'h9f30:	data_out=16'ha00;
17'h9f31:	data_out=16'h8a00;
17'h9f32:	data_out=16'h211;
17'h9f33:	data_out=16'h8a00;
17'h9f34:	data_out=16'h89ce;
17'h9f35:	data_out=16'h88f5;
17'h9f36:	data_out=16'h9c1;
17'h9f37:	data_out=16'ha00;
17'h9f38:	data_out=16'h8a00;
17'h9f39:	data_out=16'h8a00;
17'h9f3a:	data_out=16'h9e5;
17'h9f3b:	data_out=16'h89f3;
17'h9f3c:	data_out=16'h9d2;
17'h9f3d:	data_out=16'h89b4;
17'h9f3e:	data_out=16'ha00;
17'h9f3f:	data_out=16'h8a00;
17'h9f40:	data_out=16'h89b8;
17'h9f41:	data_out=16'ha00;
17'h9f42:	data_out=16'ha00;
17'h9f43:	data_out=16'h8a00;
17'h9f44:	data_out=16'h8a00;
17'h9f45:	data_out=16'h9cc;
17'h9f46:	data_out=16'h9d3;
17'h9f47:	data_out=16'h976;
17'h9f48:	data_out=16'h89c1;
17'h9f49:	data_out=16'ha00;
17'h9f4a:	data_out=16'h89ff;
17'h9f4b:	data_out=16'ha00;
17'h9f4c:	data_out=16'ha00;
17'h9f4d:	data_out=16'h89a3;
17'h9f4e:	data_out=16'h9ff;
17'h9f4f:	data_out=16'ha00;
17'h9f50:	data_out=16'h89f0;
17'h9f51:	data_out=16'ha00;
17'h9f52:	data_out=16'ha00;
17'h9f53:	data_out=16'h8a00;
17'h9f54:	data_out=16'h8a00;
17'h9f55:	data_out=16'ha00;
17'h9f56:	data_out=16'ha00;
17'h9f57:	data_out=16'h9fe;
17'h9f58:	data_out=16'h9ed;
17'h9f59:	data_out=16'h8511;
17'h9f5a:	data_out=16'h89e9;
17'h9f5b:	data_out=16'h8a00;
17'h9f5c:	data_out=16'h8a00;
17'h9f5d:	data_out=16'ha00;
17'h9f5e:	data_out=16'h8859;
17'h9f5f:	data_out=16'h8874;
17'h9f60:	data_out=16'ha00;
17'h9f61:	data_out=16'h89c3;
17'h9f62:	data_out=16'h6e4;
17'h9f63:	data_out=16'h8a00;
17'h9f64:	data_out=16'h8a00;
17'h9f65:	data_out=16'h8a00;
17'h9f66:	data_out=16'h89ff;
17'h9f67:	data_out=16'ha00;
17'h9f68:	data_out=16'ha00;
17'h9f69:	data_out=16'ha00;
17'h9f6a:	data_out=16'ha00;
17'h9f6b:	data_out=16'h8a00;
17'h9f6c:	data_out=16'h9f2;
17'h9f6d:	data_out=16'h8a00;
17'h9f6e:	data_out=16'ha00;
17'h9f6f:	data_out=16'h89b8;
17'h9f70:	data_out=16'ha00;
17'h9f71:	data_out=16'h9f1;
17'h9f72:	data_out=16'h89a4;
17'h9f73:	data_out=16'h89c0;
17'h9f74:	data_out=16'ha00;
17'h9f75:	data_out=16'h8a00;
17'h9f76:	data_out=16'h93b;
17'h9f77:	data_out=16'ha00;
17'h9f78:	data_out=16'h8a00;
17'h9f79:	data_out=16'ha00;
17'h9f7a:	data_out=16'h89f5;
17'h9f7b:	data_out=16'ha00;
17'h9f7c:	data_out=16'h85ad;
17'h9f7d:	data_out=16'h8a00;
17'h9f7e:	data_out=16'h8a00;
17'h9f7f:	data_out=16'h8a00;
17'h9f80:	data_out=16'h9d9;
17'h9f81:	data_out=16'h8987;
17'h9f82:	data_out=16'ha00;
17'h9f83:	data_out=16'h9f9;
17'h9f84:	data_out=16'h89ff;
17'h9f85:	data_out=16'h8a00;
17'h9f86:	data_out=16'h8a00;
17'h9f87:	data_out=16'ha00;
17'h9f88:	data_out=16'h9ad;
17'h9f89:	data_out=16'h83d1;
17'h9f8a:	data_out=16'h9e5;
17'h9f8b:	data_out=16'h8a00;
17'h9f8c:	data_out=16'h919;
17'h9f8d:	data_out=16'ha00;
17'h9f8e:	data_out=16'ha00;
17'h9f8f:	data_out=16'h9ff;
17'h9f90:	data_out=16'h8a00;
17'h9f91:	data_out=16'h8a00;
17'h9f92:	data_out=16'h448;
17'h9f93:	data_out=16'h9ca;
17'h9f94:	data_out=16'h8a00;
17'h9f95:	data_out=16'h654;
17'h9f96:	data_out=16'h9ee;
17'h9f97:	data_out=16'h89b7;
17'h9f98:	data_out=16'h9db;
17'h9f99:	data_out=16'h8a00;
17'h9f9a:	data_out=16'h8a00;
17'h9f9b:	data_out=16'h9fe;
17'h9f9c:	data_out=16'h8529;
17'h9f9d:	data_out=16'h8a00;
17'h9f9e:	data_out=16'h8028;
17'h9f9f:	data_out=16'h8a00;
17'h9fa0:	data_out=16'h8a00;
17'h9fa1:	data_out=16'ha00;
17'h9fa2:	data_out=16'h89f3;
17'h9fa3:	data_out=16'ha00;
17'h9fa4:	data_out=16'ha00;
17'h9fa5:	data_out=16'ha00;
17'h9fa6:	data_out=16'ha00;
17'h9fa7:	data_out=16'h8a00;
17'h9fa8:	data_out=16'ha00;
17'h9fa9:	data_out=16'ha00;
17'h9faa:	data_out=16'h9f0;
17'h9fab:	data_out=16'h8a00;
17'h9fac:	data_out=16'h9e8;
17'h9fad:	data_out=16'h8a00;
17'h9fae:	data_out=16'h989;
17'h9faf:	data_out=16'h89dd;
17'h9fb0:	data_out=16'h8180;
17'h9fb1:	data_out=16'h89fa;
17'h9fb2:	data_out=16'h89db;
17'h9fb3:	data_out=16'h8a00;
17'h9fb4:	data_out=16'h88fb;
17'h9fb5:	data_out=16'h870f;
17'h9fb6:	data_out=16'h9e9;
17'h9fb7:	data_out=16'ha00;
17'h9fb8:	data_out=16'h8a00;
17'h9fb9:	data_out=16'h8a00;
17'h9fba:	data_out=16'h52;
17'h9fbb:	data_out=16'h3e7;
17'h9fbc:	data_out=16'h9ee;
17'h9fbd:	data_out=16'h89e8;
17'h9fbe:	data_out=16'ha00;
17'h9fbf:	data_out=16'h8a00;
17'h9fc0:	data_out=16'h8a00;
17'h9fc1:	data_out=16'ha00;
17'h9fc2:	data_out=16'ha00;
17'h9fc3:	data_out=16'h8a00;
17'h9fc4:	data_out=16'h8a00;
17'h9fc5:	data_out=16'h9c6;
17'h9fc6:	data_out=16'h9f2;
17'h9fc7:	data_out=16'h837;
17'h9fc8:	data_out=16'h89d4;
17'h9fc9:	data_out=16'ha00;
17'h9fca:	data_out=16'h8a00;
17'h9fcb:	data_out=16'h273;
17'h9fcc:	data_out=16'ha00;
17'h9fcd:	data_out=16'h8a00;
17'h9fce:	data_out=16'h9ff;
17'h9fcf:	data_out=16'ha00;
17'h9fd0:	data_out=16'h8a00;
17'h9fd1:	data_out=16'h9ff;
17'h9fd2:	data_out=16'ha00;
17'h9fd3:	data_out=16'h8a00;
17'h9fd4:	data_out=16'h8a00;
17'h9fd5:	data_out=16'h9ff;
17'h9fd6:	data_out=16'ha00;
17'h9fd7:	data_out=16'h9fd;
17'h9fd8:	data_out=16'h9fe;
17'h9fd9:	data_out=16'h89e7;
17'h9fda:	data_out=16'h89d9;
17'h9fdb:	data_out=16'h8a00;
17'h9fdc:	data_out=16'h501;
17'h9fdd:	data_out=16'h9fc;
17'h9fde:	data_out=16'h8370;
17'h9fdf:	data_out=16'h89b3;
17'h9fe0:	data_out=16'ha00;
17'h9fe1:	data_out=16'h89f3;
17'h9fe2:	data_out=16'h8519;
17'h9fe3:	data_out=16'h8a00;
17'h9fe4:	data_out=16'h8a00;
17'h9fe5:	data_out=16'h8a00;
17'h9fe6:	data_out=16'h8a00;
17'h9fe7:	data_out=16'h8f2;
17'h9fe8:	data_out=16'ha00;
17'h9fe9:	data_out=16'ha00;
17'h9fea:	data_out=16'ha00;
17'h9feb:	data_out=16'h8a00;
17'h9fec:	data_out=16'h9f8;
17'h9fed:	data_out=16'h8a00;
17'h9fee:	data_out=16'ha00;
17'h9fef:	data_out=16'h89e6;
17'h9ff0:	data_out=16'ha00;
17'h9ff1:	data_out=16'h9fa;
17'h9ff2:	data_out=16'h89da;
17'h9ff3:	data_out=16'h89f0;
17'h9ff4:	data_out=16'h4f5;
17'h9ff5:	data_out=16'h9e2;
17'h9ff6:	data_out=16'h8a00;
17'h9ff7:	data_out=16'h9ed;
17'h9ff8:	data_out=16'h8a00;
17'h9ff9:	data_out=16'ha00;
17'h9ffa:	data_out=16'h8a00;
17'h9ffb:	data_out=16'ha00;
17'h9ffc:	data_out=16'h851;
17'h9ffd:	data_out=16'h8a00;
17'h9ffe:	data_out=16'h8a00;
17'h9fff:	data_out=16'h8a00;
17'ha000:	data_out=16'h9b1;
17'ha001:	data_out=16'h8211;
17'ha002:	data_out=16'ha00;
17'ha003:	data_out=16'h894d;
17'ha004:	data_out=16'h89fe;
17'ha005:	data_out=16'h89eb;
17'ha006:	data_out=16'h89f8;
17'ha007:	data_out=16'ha00;
17'ha008:	data_out=16'h96a;
17'ha009:	data_out=16'h89e2;
17'ha00a:	data_out=16'h880e;
17'ha00b:	data_out=16'h8a00;
17'ha00c:	data_out=16'h9c4;
17'ha00d:	data_out=16'ha00;
17'ha00e:	data_out=16'ha00;
17'ha00f:	data_out=16'h9fe;
17'ha010:	data_out=16'h8a00;
17'ha011:	data_out=16'h8a00;
17'ha012:	data_out=16'h89f3;
17'ha013:	data_out=16'h871e;
17'ha014:	data_out=16'h8a00;
17'ha015:	data_out=16'h8783;
17'ha016:	data_out=16'h693;
17'ha017:	data_out=16'h89ea;
17'ha018:	data_out=16'h9ac;
17'ha019:	data_out=16'h8a00;
17'ha01a:	data_out=16'h8a00;
17'ha01b:	data_out=16'h3cc;
17'ha01c:	data_out=16'h8995;
17'ha01d:	data_out=16'h89f0;
17'ha01e:	data_out=16'h89ff;
17'ha01f:	data_out=16'h8a00;
17'ha020:	data_out=16'h8a00;
17'ha021:	data_out=16'ha00;
17'ha022:	data_out=16'h89f9;
17'ha023:	data_out=16'ha00;
17'ha024:	data_out=16'ha00;
17'ha025:	data_out=16'h891d;
17'ha026:	data_out=16'ha00;
17'ha027:	data_out=16'h8a00;
17'ha028:	data_out=16'ha00;
17'ha029:	data_out=16'h7bf;
17'ha02a:	data_out=16'h9d8;
17'ha02b:	data_out=16'h8a00;
17'ha02c:	data_out=16'h83a1;
17'ha02d:	data_out=16'h8a00;
17'ha02e:	data_out=16'h89f3;
17'ha02f:	data_out=16'h89b3;
17'ha030:	data_out=16'h8900;
17'ha031:	data_out=16'h89be;
17'ha032:	data_out=16'h8a00;
17'ha033:	data_out=16'h8a00;
17'ha034:	data_out=16'h56b;
17'ha035:	data_out=16'h8a00;
17'ha036:	data_out=16'h969;
17'ha037:	data_out=16'h9ff;
17'ha038:	data_out=16'h899e;
17'ha039:	data_out=16'h8a00;
17'ha03a:	data_out=16'h89fe;
17'ha03b:	data_out=16'h82f;
17'ha03c:	data_out=16'h87c;
17'ha03d:	data_out=16'h8a00;
17'ha03e:	data_out=16'ha00;
17'ha03f:	data_out=16'h89ea;
17'ha040:	data_out=16'h8a00;
17'ha041:	data_out=16'ha00;
17'ha042:	data_out=16'h9ff;
17'ha043:	data_out=16'h8a00;
17'ha044:	data_out=16'h8a00;
17'ha045:	data_out=16'h8716;
17'ha046:	data_out=16'h91d;
17'ha047:	data_out=16'h89fe;
17'ha048:	data_out=16'h8996;
17'ha049:	data_out=16'h89ac;
17'ha04a:	data_out=16'h89fd;
17'ha04b:	data_out=16'h8680;
17'ha04c:	data_out=16'ha00;
17'ha04d:	data_out=16'h8a00;
17'ha04e:	data_out=16'h9fe;
17'ha04f:	data_out=16'h9fc;
17'ha050:	data_out=16'h8a00;
17'ha051:	data_out=16'h9f4;
17'ha052:	data_out=16'ha00;
17'ha053:	data_out=16'h89ff;
17'ha054:	data_out=16'h8a00;
17'ha055:	data_out=16'h84a;
17'ha056:	data_out=16'ha00;
17'ha057:	data_out=16'h89e6;
17'ha058:	data_out=16'h9fa;
17'ha059:	data_out=16'h8a00;
17'ha05a:	data_out=16'h9d0;
17'ha05b:	data_out=16'h8a00;
17'ha05c:	data_out=16'ha00;
17'ha05d:	data_out=16'h9fc;
17'ha05e:	data_out=16'h85c4;
17'ha05f:	data_out=16'h8a00;
17'ha060:	data_out=16'h9e4;
17'ha061:	data_out=16'h8a00;
17'ha062:	data_out=16'h89c5;
17'ha063:	data_out=16'h8a00;
17'ha064:	data_out=16'h8a00;
17'ha065:	data_out=16'h89ff;
17'ha066:	data_out=16'h8a00;
17'ha067:	data_out=16'h8a00;
17'ha068:	data_out=16'ha00;
17'ha069:	data_out=16'h9ea;
17'ha06a:	data_out=16'ha00;
17'ha06b:	data_out=16'h8a00;
17'ha06c:	data_out=16'h9f9;
17'ha06d:	data_out=16'h8a00;
17'ha06e:	data_out=16'ha00;
17'ha06f:	data_out=16'h8932;
17'ha070:	data_out=16'ha00;
17'ha071:	data_out=16'h9aa;
17'ha072:	data_out=16'h89c6;
17'ha073:	data_out=16'h89e2;
17'ha074:	data_out=16'h8605;
17'ha075:	data_out=16'h9ff;
17'ha076:	data_out=16'h8a00;
17'ha077:	data_out=16'h89c1;
17'ha078:	data_out=16'h8a00;
17'ha079:	data_out=16'ha00;
17'ha07a:	data_out=16'h8a00;
17'ha07b:	data_out=16'ha00;
17'ha07c:	data_out=16'h671;
17'ha07d:	data_out=16'h8a00;
17'ha07e:	data_out=16'h8a00;
17'ha07f:	data_out=16'h8a00;
17'ha080:	data_out=16'h9fd;
17'ha081:	data_out=16'h9ed;
17'ha082:	data_out=16'h3a9;
17'ha083:	data_out=16'h8998;
17'ha084:	data_out=16'h8a00;
17'ha085:	data_out=16'h9f1;
17'ha086:	data_out=16'h89fb;
17'ha087:	data_out=16'h975;
17'ha088:	data_out=16'h9a6;
17'ha089:	data_out=16'h8a00;
17'ha08a:	data_out=16'h7c3;
17'ha08b:	data_out=16'h8a00;
17'ha08c:	data_out=16'h975;
17'ha08d:	data_out=16'ha00;
17'ha08e:	data_out=16'h9fd;
17'ha08f:	data_out=16'h89fe;
17'ha090:	data_out=16'h8a00;
17'ha091:	data_out=16'h8a00;
17'ha092:	data_out=16'h8a00;
17'ha093:	data_out=16'h898b;
17'ha094:	data_out=16'h8a00;
17'ha095:	data_out=16'h89f2;
17'ha096:	data_out=16'h8f0;
17'ha097:	data_out=16'h89cd;
17'ha098:	data_out=16'h8a00;
17'ha099:	data_out=16'h8a00;
17'ha09a:	data_out=16'h8a00;
17'ha09b:	data_out=16'h8896;
17'ha09c:	data_out=16'h8370;
17'ha09d:	data_out=16'h89da;
17'ha09e:	data_out=16'h8a00;
17'ha09f:	data_out=16'h8a00;
17'ha0a0:	data_out=16'h8a00;
17'ha0a1:	data_out=16'h9fd;
17'ha0a2:	data_out=16'h8a00;
17'ha0a3:	data_out=16'h590;
17'ha0a4:	data_out=16'h600;
17'ha0a5:	data_out=16'h8a00;
17'ha0a6:	data_out=16'h897d;
17'ha0a7:	data_out=16'h8a00;
17'ha0a8:	data_out=16'h9fb;
17'ha0a9:	data_out=16'h89d4;
17'ha0aa:	data_out=16'h89fc;
17'ha0ab:	data_out=16'h8a00;
17'ha0ac:	data_out=16'h41c;
17'ha0ad:	data_out=16'h8a00;
17'ha0ae:	data_out=16'h8a00;
17'ha0af:	data_out=16'h89b3;
17'ha0b0:	data_out=16'h99f;
17'ha0b1:	data_out=16'h9d3;
17'ha0b2:	data_out=16'h8a00;
17'ha0b3:	data_out=16'h8a00;
17'ha0b4:	data_out=16'ha00;
17'ha0b5:	data_out=16'h8a00;
17'ha0b6:	data_out=16'h893d;
17'ha0b7:	data_out=16'h89d9;
17'ha0b8:	data_out=16'ha00;
17'ha0b9:	data_out=16'h8a00;
17'ha0ba:	data_out=16'h8a00;
17'ha0bb:	data_out=16'h8da;
17'ha0bc:	data_out=16'h8e8;
17'ha0bd:	data_out=16'h8a00;
17'ha0be:	data_out=16'h9fb;
17'ha0bf:	data_out=16'h9f7;
17'ha0c0:	data_out=16'h8a00;
17'ha0c1:	data_out=16'ha00;
17'ha0c2:	data_out=16'h9ff;
17'ha0c3:	data_out=16'h8a00;
17'ha0c4:	data_out=16'h8a00;
17'ha0c5:	data_out=16'h89f0;
17'ha0c6:	data_out=16'h95f;
17'ha0c7:	data_out=16'h8a00;
17'ha0c8:	data_out=16'h89f0;
17'ha0c9:	data_out=16'h8a00;
17'ha0ca:	data_out=16'h86ca;
17'ha0cb:	data_out=16'h81c1;
17'ha0cc:	data_out=16'h89e0;
17'ha0cd:	data_out=16'h8a00;
17'ha0ce:	data_out=16'h8607;
17'ha0cf:	data_out=16'h8a00;
17'ha0d0:	data_out=16'h8a00;
17'ha0d1:	data_out=16'h583;
17'ha0d2:	data_out=16'h9ea;
17'ha0d3:	data_out=16'h89ef;
17'ha0d4:	data_out=16'h8a00;
17'ha0d5:	data_out=16'h89d7;
17'ha0d6:	data_out=16'h3fa;
17'ha0d7:	data_out=16'h8a00;
17'ha0d8:	data_out=16'h9f9;
17'ha0d9:	data_out=16'h8a00;
17'ha0da:	data_out=16'h9f4;
17'ha0db:	data_out=16'h8a00;
17'ha0dc:	data_out=16'ha00;
17'ha0dd:	data_out=16'h8277;
17'ha0de:	data_out=16'h8858;
17'ha0df:	data_out=16'h8a00;
17'ha0e0:	data_out=16'h89e4;
17'ha0e1:	data_out=16'h8a00;
17'ha0e2:	data_out=16'h89c9;
17'ha0e3:	data_out=16'h8a00;
17'ha0e4:	data_out=16'h89f7;
17'ha0e5:	data_out=16'h8a00;
17'ha0e6:	data_out=16'h8a00;
17'ha0e7:	data_out=16'h8a00;
17'ha0e8:	data_out=16'h9fd;
17'ha0e9:	data_out=16'h8172;
17'ha0ea:	data_out=16'h9fd;
17'ha0eb:	data_out=16'h89f9;
17'ha0ec:	data_out=16'h9ff;
17'ha0ed:	data_out=16'h8a00;
17'ha0ee:	data_out=16'h9fd;
17'ha0ef:	data_out=16'h86dd;
17'ha0f0:	data_out=16'h9fd;
17'ha0f1:	data_out=16'h89ff;
17'ha0f2:	data_out=16'h8a00;
17'ha0f3:	data_out=16'h89f6;
17'ha0f4:	data_out=16'h9fe;
17'ha0f5:	data_out=16'ha00;
17'ha0f6:	data_out=16'h8a00;
17'ha0f7:	data_out=16'h8a00;
17'ha0f8:	data_out=16'h8a00;
17'ha0f9:	data_out=16'ha00;
17'ha0fa:	data_out=16'h8a00;
17'ha0fb:	data_out=16'h9fb;
17'ha0fc:	data_out=16'h8a00;
17'ha0fd:	data_out=16'h8a00;
17'ha0fe:	data_out=16'h8a00;
17'ha0ff:	data_out=16'h89d5;
17'ha100:	data_out=16'ha00;
17'ha101:	data_out=16'h9fd;
17'ha102:	data_out=16'h8a00;
17'ha103:	data_out=16'h191;
17'ha104:	data_out=16'h8a00;
17'ha105:	data_out=16'ha00;
17'ha106:	data_out=16'h89e1;
17'ha107:	data_out=16'h8a00;
17'ha108:	data_out=16'h597;
17'ha109:	data_out=16'h8a00;
17'ha10a:	data_out=16'h8a00;
17'ha10b:	data_out=16'h8a00;
17'ha10c:	data_out=16'h89fd;
17'ha10d:	data_out=16'h9fc;
17'ha10e:	data_out=16'h89fb;
17'ha10f:	data_out=16'h8a00;
17'ha110:	data_out=16'h8a00;
17'ha111:	data_out=16'h8a00;
17'ha112:	data_out=16'h89ef;
17'ha113:	data_out=16'h293;
17'ha114:	data_out=16'h89bf;
17'ha115:	data_out=16'h8732;
17'ha116:	data_out=16'h9c8;
17'ha117:	data_out=16'h9df;
17'ha118:	data_out=16'h8a00;
17'ha119:	data_out=16'h8a00;
17'ha11a:	data_out=16'h8804;
17'ha11b:	data_out=16'h29d;
17'ha11c:	data_out=16'ha00;
17'ha11d:	data_out=16'h805e;
17'ha11e:	data_out=16'h89ff;
17'ha11f:	data_out=16'h8a00;
17'ha120:	data_out=16'h89f5;
17'ha121:	data_out=16'h89fa;
17'ha122:	data_out=16'h8a00;
17'ha123:	data_out=16'h8a00;
17'ha124:	data_out=16'h8a00;
17'ha125:	data_out=16'h8a00;
17'ha126:	data_out=16'h8a00;
17'ha127:	data_out=16'h8a00;
17'ha128:	data_out=16'h89f9;
17'ha129:	data_out=16'h8a00;
17'ha12a:	data_out=16'h89ff;
17'ha12b:	data_out=16'h8a00;
17'ha12c:	data_out=16'h97e;
17'ha12d:	data_out=16'h8a00;
17'ha12e:	data_out=16'h89ff;
17'ha12f:	data_out=16'h9fe;
17'ha130:	data_out=16'h89ef;
17'ha131:	data_out=16'h99f;
17'ha132:	data_out=16'h8a00;
17'ha133:	data_out=16'h89da;
17'ha134:	data_out=16'ha00;
17'ha135:	data_out=16'h8a00;
17'ha136:	data_out=16'h89ef;
17'ha137:	data_out=16'h8a00;
17'ha138:	data_out=16'ha00;
17'ha139:	data_out=16'h89f0;
17'ha13a:	data_out=16'h8a00;
17'ha13b:	data_out=16'h8a00;
17'ha13c:	data_out=16'h9d4;
17'ha13d:	data_out=16'h8a00;
17'ha13e:	data_out=16'h89ef;
17'ha13f:	data_out=16'ha00;
17'ha140:	data_out=16'h8a00;
17'ha141:	data_out=16'ha00;
17'ha142:	data_out=16'h89e5;
17'ha143:	data_out=16'h8a00;
17'ha144:	data_out=16'h812a;
17'ha145:	data_out=16'h84f0;
17'ha146:	data_out=16'h8558;
17'ha147:	data_out=16'h8a00;
17'ha148:	data_out=16'h89b7;
17'ha149:	data_out=16'h8a00;
17'ha14a:	data_out=16'h89f5;
17'ha14b:	data_out=16'h89f6;
17'ha14c:	data_out=16'h8a00;
17'ha14d:	data_out=16'h8a00;
17'ha14e:	data_out=16'h806f;
17'ha14f:	data_out=16'h8a00;
17'ha150:	data_out=16'h86ed;
17'ha151:	data_out=16'h7f2;
17'ha152:	data_out=16'h8a00;
17'ha153:	data_out=16'h5e1;
17'ha154:	data_out=16'h89ec;
17'ha155:	data_out=16'h89f9;
17'ha156:	data_out=16'h8a00;
17'ha157:	data_out=16'h8a00;
17'ha158:	data_out=16'ha00;
17'ha159:	data_out=16'h8a00;
17'ha15a:	data_out=16'ha00;
17'ha15b:	data_out=16'h8a00;
17'ha15c:	data_out=16'ha00;
17'ha15d:	data_out=16'h693;
17'ha15e:	data_out=16'ha00;
17'ha15f:	data_out=16'h8a00;
17'ha160:	data_out=16'h8a00;
17'ha161:	data_out=16'h87af;
17'ha162:	data_out=16'h873c;
17'ha163:	data_out=16'h89b2;
17'ha164:	data_out=16'h8666;
17'ha165:	data_out=16'h8a00;
17'ha166:	data_out=16'h8a00;
17'ha167:	data_out=16'h8a00;
17'ha168:	data_out=16'h89fa;
17'ha169:	data_out=16'h8a00;
17'ha16a:	data_out=16'h89fb;
17'ha16b:	data_out=16'h89f4;
17'ha16c:	data_out=16'ha00;
17'ha16d:	data_out=16'h89bc;
17'ha16e:	data_out=16'h89fb;
17'ha16f:	data_out=16'h9da;
17'ha170:	data_out=16'h89fb;
17'ha171:	data_out=16'h89ff;
17'ha172:	data_out=16'h8a00;
17'ha173:	data_out=16'h8305;
17'ha174:	data_out=16'h892c;
17'ha175:	data_out=16'ha00;
17'ha176:	data_out=16'h8a00;
17'ha177:	data_out=16'h8a00;
17'ha178:	data_out=16'h8a00;
17'ha179:	data_out=16'h850a;
17'ha17a:	data_out=16'h8619;
17'ha17b:	data_out=16'h89de;
17'ha17c:	data_out=16'h8a00;
17'ha17d:	data_out=16'h8a00;
17'ha17e:	data_out=16'h8a00;
17'ha17f:	data_out=16'hd3;
17'ha180:	data_out=16'h949;
17'ha181:	data_out=16'h95f;
17'ha182:	data_out=16'h8a00;
17'ha183:	data_out=16'h6b5;
17'ha184:	data_out=16'h8a00;
17'ha185:	data_out=16'h818f;
17'ha186:	data_out=16'h8612;
17'ha187:	data_out=16'h8a00;
17'ha188:	data_out=16'h255;
17'ha189:	data_out=16'h8a00;
17'ha18a:	data_out=16'h8a00;
17'ha18b:	data_out=16'h8a00;
17'ha18c:	data_out=16'h8a00;
17'ha18d:	data_out=16'ha00;
17'ha18e:	data_out=16'h8a00;
17'ha18f:	data_out=16'h89ff;
17'ha190:	data_out=16'h8a00;
17'ha191:	data_out=16'h8a00;
17'ha192:	data_out=16'ha00;
17'ha193:	data_out=16'h9fb;
17'ha194:	data_out=16'h9f1;
17'ha195:	data_out=16'h8a00;
17'ha196:	data_out=16'h838;
17'ha197:	data_out=16'ha00;
17'ha198:	data_out=16'h8a00;
17'ha199:	data_out=16'h8a00;
17'ha19a:	data_out=16'h8a00;
17'ha19b:	data_out=16'h709;
17'ha19c:	data_out=16'h9cf;
17'ha19d:	data_out=16'h89f1;
17'ha19e:	data_out=16'h520;
17'ha19f:	data_out=16'h89ad;
17'ha1a0:	data_out=16'h89eb;
17'ha1a1:	data_out=16'h8a00;
17'ha1a2:	data_out=16'h8a00;
17'ha1a3:	data_out=16'h8a00;
17'ha1a4:	data_out=16'h8a00;
17'ha1a5:	data_out=16'h8a00;
17'ha1a6:	data_out=16'h8a00;
17'ha1a7:	data_out=16'h8a00;
17'ha1a8:	data_out=16'h89fd;
17'ha1a9:	data_out=16'h8a00;
17'ha1aa:	data_out=16'h89ff;
17'ha1ab:	data_out=16'h8187;
17'ha1ac:	data_out=16'h78c;
17'ha1ad:	data_out=16'h8a00;
17'ha1ae:	data_out=16'h89c2;
17'ha1af:	data_out=16'h9ee;
17'ha1b0:	data_out=16'h8a00;
17'ha1b1:	data_out=16'h8a00;
17'ha1b2:	data_out=16'h8a00;
17'ha1b3:	data_out=16'ha00;
17'ha1b4:	data_out=16'h9cb;
17'ha1b5:	data_out=16'h8a00;
17'ha1b6:	data_out=16'h89f3;
17'ha1b7:	data_out=16'h8a00;
17'ha1b8:	data_out=16'ha00;
17'ha1b9:	data_out=16'ha00;
17'ha1ba:	data_out=16'h8a00;
17'ha1bb:	data_out=16'h8a00;
17'ha1bc:	data_out=16'h65c;
17'ha1bd:	data_out=16'h8a00;
17'ha1be:	data_out=16'h89fd;
17'ha1bf:	data_out=16'h81ad;
17'ha1c0:	data_out=16'h8a00;
17'ha1c1:	data_out=16'h9ff;
17'ha1c2:	data_out=16'h8a00;
17'ha1c3:	data_out=16'h8a00;
17'ha1c4:	data_out=16'h8a00;
17'ha1c5:	data_out=16'h8a00;
17'ha1c6:	data_out=16'h8a00;
17'ha1c7:	data_out=16'h8a00;
17'ha1c8:	data_out=16'h5bd;
17'ha1c9:	data_out=16'h8a00;
17'ha1ca:	data_out=16'h88b4;
17'ha1cb:	data_out=16'h8a00;
17'ha1cc:	data_out=16'h8a00;
17'ha1cd:	data_out=16'h8a00;
17'ha1ce:	data_out=16'h77e;
17'ha1cf:	data_out=16'h8a00;
17'ha1d0:	data_out=16'h42d;
17'ha1d1:	data_out=16'h9cb;
17'ha1d2:	data_out=16'h8a00;
17'ha1d3:	data_out=16'h9bc;
17'ha1d4:	data_out=16'h8536;
17'ha1d5:	data_out=16'h8a00;
17'ha1d6:	data_out=16'h8a00;
17'ha1d7:	data_out=16'h8a00;
17'ha1d8:	data_out=16'ha00;
17'ha1d9:	data_out=16'h8a00;
17'ha1da:	data_out=16'ha00;
17'ha1db:	data_out=16'h8a00;
17'ha1dc:	data_out=16'ha00;
17'ha1dd:	data_out=16'h89ee;
17'ha1de:	data_out=16'ha00;
17'ha1df:	data_out=16'h89fc;
17'ha1e0:	data_out=16'h8a00;
17'ha1e1:	data_out=16'h8a00;
17'ha1e2:	data_out=16'h9b4;
17'ha1e3:	data_out=16'ha00;
17'ha1e4:	data_out=16'h8626;
17'ha1e5:	data_out=16'h8a00;
17'ha1e6:	data_out=16'h8a00;
17'ha1e7:	data_out=16'h8a00;
17'ha1e8:	data_out=16'h89fe;
17'ha1e9:	data_out=16'h8a00;
17'ha1ea:	data_out=16'h8a00;
17'ha1eb:	data_out=16'h8a00;
17'ha1ec:	data_out=16'h98b;
17'ha1ed:	data_out=16'ha00;
17'ha1ee:	data_out=16'h8a00;
17'ha1ef:	data_out=16'h89f8;
17'ha1f0:	data_out=16'h8a00;
17'ha1f1:	data_out=16'h4da;
17'ha1f2:	data_out=16'h8a00;
17'ha1f3:	data_out=16'h8a00;
17'ha1f4:	data_out=16'h8a00;
17'ha1f5:	data_out=16'h9bc;
17'ha1f6:	data_out=16'h8a00;
17'ha1f7:	data_out=16'h8a00;
17'ha1f8:	data_out=16'h89f9;
17'ha1f9:	data_out=16'h88d9;
17'ha1fa:	data_out=16'ha00;
17'ha1fb:	data_out=16'h89fd;
17'ha1fc:	data_out=16'h89fb;
17'ha1fd:	data_out=16'h89c4;
17'ha1fe:	data_out=16'h89ae;
17'ha1ff:	data_out=16'h1d1;
17'ha200:	data_out=16'h89fc;
17'ha201:	data_out=16'h8a00;
17'ha202:	data_out=16'h8a00;
17'ha203:	data_out=16'h4f5;
17'ha204:	data_out=16'h8a00;
17'ha205:	data_out=16'h8a00;
17'ha206:	data_out=16'h9ff;
17'ha207:	data_out=16'h8a00;
17'ha208:	data_out=16'h233;
17'ha209:	data_out=16'h8a00;
17'ha20a:	data_out=16'h8a00;
17'ha20b:	data_out=16'h8f2;
17'ha20c:	data_out=16'h8a00;
17'ha20d:	data_out=16'h8f1;
17'ha20e:	data_out=16'h89fe;
17'ha20f:	data_out=16'h89fd;
17'ha210:	data_out=16'h8a00;
17'ha211:	data_out=16'h8a00;
17'ha212:	data_out=16'ha00;
17'ha213:	data_out=16'h4aa;
17'ha214:	data_out=16'h9a3;
17'ha215:	data_out=16'h8a00;
17'ha216:	data_out=16'h8a00;
17'ha217:	data_out=16'h9ec;
17'ha218:	data_out=16'h89fd;
17'ha219:	data_out=16'h8a00;
17'ha21a:	data_out=16'h8a00;
17'ha21b:	data_out=16'h798;
17'ha21c:	data_out=16'h965;
17'ha21d:	data_out=16'h89f7;
17'ha21e:	data_out=16'h75d;
17'ha21f:	data_out=16'h515;
17'ha220:	data_out=16'h89f6;
17'ha221:	data_out=16'h89fa;
17'ha222:	data_out=16'h89ed;
17'ha223:	data_out=16'h8a00;
17'ha224:	data_out=16'h8a00;
17'ha225:	data_out=16'h8a00;
17'ha226:	data_out=16'h8a00;
17'ha227:	data_out=16'h8a00;
17'ha228:	data_out=16'h89f5;
17'ha229:	data_out=16'h8a00;
17'ha22a:	data_out=16'h8a00;
17'ha22b:	data_out=16'h9f5;
17'ha22c:	data_out=16'h8a00;
17'ha22d:	data_out=16'h475;
17'ha22e:	data_out=16'h9df;
17'ha22f:	data_out=16'h9e7;
17'ha230:	data_out=16'h8a00;
17'ha231:	data_out=16'h8a00;
17'ha232:	data_out=16'h8a00;
17'ha233:	data_out=16'ha00;
17'ha234:	data_out=16'h5a7;
17'ha235:	data_out=16'h8a00;
17'ha236:	data_out=16'h85fb;
17'ha237:	data_out=16'h8a00;
17'ha238:	data_out=16'ha00;
17'ha239:	data_out=16'ha00;
17'ha23a:	data_out=16'h8a00;
17'ha23b:	data_out=16'h8a00;
17'ha23c:	data_out=16'h89e1;
17'ha23d:	data_out=16'h8a00;
17'ha23e:	data_out=16'h89f5;
17'ha23f:	data_out=16'h8a00;
17'ha240:	data_out=16'h8a00;
17'ha241:	data_out=16'h986;
17'ha242:	data_out=16'h8a00;
17'ha243:	data_out=16'h8a00;
17'ha244:	data_out=16'h8a00;
17'ha245:	data_out=16'h8a00;
17'ha246:	data_out=16'h8a00;
17'ha247:	data_out=16'h8a00;
17'ha248:	data_out=16'h9f7;
17'ha249:	data_out=16'h8a00;
17'ha24a:	data_out=16'h2fc;
17'ha24b:	data_out=16'h8a00;
17'ha24c:	data_out=16'h8a00;
17'ha24d:	data_out=16'h89df;
17'ha24e:	data_out=16'h968;
17'ha24f:	data_out=16'h8a00;
17'ha250:	data_out=16'h8a00;
17'ha251:	data_out=16'h780;
17'ha252:	data_out=16'h8a00;
17'ha253:	data_out=16'h9c3;
17'ha254:	data_out=16'h84ba;
17'ha255:	data_out=16'h8a00;
17'ha256:	data_out=16'h8a00;
17'ha257:	data_out=16'h8a00;
17'ha258:	data_out=16'h9be;
17'ha259:	data_out=16'h8a00;
17'ha25a:	data_out=16'ha00;
17'ha25b:	data_out=16'h8a00;
17'ha25c:	data_out=16'h9e9;
17'ha25d:	data_out=16'h89f0;
17'ha25e:	data_out=16'ha00;
17'ha25f:	data_out=16'h88b7;
17'ha260:	data_out=16'h8a00;
17'ha261:	data_out=16'h8a00;
17'ha262:	data_out=16'h9c6;
17'ha263:	data_out=16'ha00;
17'ha264:	data_out=16'h89f4;
17'ha265:	data_out=16'h8a00;
17'ha266:	data_out=16'h8a00;
17'ha267:	data_out=16'h8a00;
17'ha268:	data_out=16'h89f7;
17'ha269:	data_out=16'h8a00;
17'ha26a:	data_out=16'h8a00;
17'ha26b:	data_out=16'h8a00;
17'ha26c:	data_out=16'h89f5;
17'ha26d:	data_out=16'ha00;
17'ha26e:	data_out=16'h8a00;
17'ha26f:	data_out=16'h8a00;
17'ha270:	data_out=16'h89ff;
17'ha271:	data_out=16'h8f5;
17'ha272:	data_out=16'h8a00;
17'ha273:	data_out=16'h8a00;
17'ha274:	data_out=16'h8a00;
17'ha275:	data_out=16'h8501;
17'ha276:	data_out=16'h89cf;
17'ha277:	data_out=16'h8a00;
17'ha278:	data_out=16'h8971;
17'ha279:	data_out=16'h813d;
17'ha27a:	data_out=16'h9fe;
17'ha27b:	data_out=16'h89f5;
17'ha27c:	data_out=16'h8518;
17'ha27d:	data_out=16'h89ba;
17'ha27e:	data_out=16'h389;
17'ha27f:	data_out=16'h89ed;
17'ha280:	data_out=16'h8a00;
17'ha281:	data_out=16'h89df;
17'ha282:	data_out=16'h8a00;
17'ha283:	data_out=16'h87de;
17'ha284:	data_out=16'h8a00;
17'ha285:	data_out=16'h8a00;
17'ha286:	data_out=16'h9fe;
17'ha287:	data_out=16'h8a00;
17'ha288:	data_out=16'h8176;
17'ha289:	data_out=16'h89a2;
17'ha28a:	data_out=16'h8a00;
17'ha28b:	data_out=16'ha00;
17'ha28c:	data_out=16'h89d5;
17'ha28d:	data_out=16'h8a00;
17'ha28e:	data_out=16'h1d4;
17'ha28f:	data_out=16'h897c;
17'ha290:	data_out=16'h869f;
17'ha291:	data_out=16'h88f4;
17'ha292:	data_out=16'h9af;
17'ha293:	data_out=16'h1a6;
17'ha294:	data_out=16'h9ef;
17'ha295:	data_out=16'h8a00;
17'ha296:	data_out=16'h8a00;
17'ha297:	data_out=16'h9fb;
17'ha298:	data_out=16'h8a00;
17'ha299:	data_out=16'h8974;
17'ha29a:	data_out=16'h8a00;
17'ha29b:	data_out=16'h99e;
17'ha29c:	data_out=16'h86b4;
17'ha29d:	data_out=16'h83af;
17'ha29e:	data_out=16'h975;
17'ha29f:	data_out=16'h99d;
17'ha2a0:	data_out=16'h89f1;
17'ha2a1:	data_out=16'h3b6;
17'ha2a2:	data_out=16'h888e;
17'ha2a3:	data_out=16'h8a00;
17'ha2a4:	data_out=16'h8a00;
17'ha2a5:	data_out=16'h8a00;
17'ha2a6:	data_out=16'h89ff;
17'ha2a7:	data_out=16'h89cd;
17'ha2a8:	data_out=16'h6cc;
17'ha2a9:	data_out=16'h861;
17'ha2aa:	data_out=16'h8a00;
17'ha2ab:	data_out=16'ha00;
17'ha2ac:	data_out=16'h8a00;
17'ha2ad:	data_out=16'ha00;
17'ha2ae:	data_out=16'h9d5;
17'ha2af:	data_out=16'h299;
17'ha2b0:	data_out=16'h8a00;
17'ha2b1:	data_out=16'h8a00;
17'ha2b2:	data_out=16'h8a00;
17'ha2b3:	data_out=16'h9fd;
17'ha2b4:	data_out=16'h84de;
17'ha2b5:	data_out=16'h8a00;
17'ha2b6:	data_out=16'h8457;
17'ha2b7:	data_out=16'hbb;
17'ha2b8:	data_out=16'ha00;
17'ha2b9:	data_out=16'h9fd;
17'ha2ba:	data_out=16'h8a00;
17'ha2bb:	data_out=16'h8a00;
17'ha2bc:	data_out=16'h8493;
17'ha2bd:	data_out=16'h8a00;
17'ha2be:	data_out=16'h6dc;
17'ha2bf:	data_out=16'h8a00;
17'ha2c0:	data_out=16'h8a00;
17'ha2c1:	data_out=16'h8a00;
17'ha2c2:	data_out=16'h8a00;
17'ha2c3:	data_out=16'h8a00;
17'ha2c4:	data_out=16'h8a00;
17'ha2c5:	data_out=16'h8a00;
17'ha2c6:	data_out=16'h9e8;
17'ha2c7:	data_out=16'h89d1;
17'ha2c8:	data_out=16'h9f1;
17'ha2c9:	data_out=16'h8a00;
17'ha2ca:	data_out=16'h998;
17'ha2cb:	data_out=16'h89bf;
17'ha2cc:	data_out=16'h8a00;
17'ha2cd:	data_out=16'h87fd;
17'ha2ce:	data_out=16'h9d9;
17'ha2cf:	data_out=16'h8a00;
17'ha2d0:	data_out=16'h89f7;
17'ha2d1:	data_out=16'h89fc;
17'ha2d2:	data_out=16'h8a00;
17'ha2d3:	data_out=16'h9c0;
17'ha2d4:	data_out=16'h872b;
17'ha2d5:	data_out=16'h80c4;
17'ha2d6:	data_out=16'h8a00;
17'ha2d7:	data_out=16'h8a00;
17'ha2d8:	data_out=16'h86ad;
17'ha2d9:	data_out=16'h8a00;
17'ha2da:	data_out=16'h9fc;
17'ha2db:	data_out=16'h8a00;
17'ha2dc:	data_out=16'h9d9;
17'ha2dd:	data_out=16'h89a4;
17'ha2de:	data_out=16'h2aa;
17'ha2df:	data_out=16'h88b4;
17'ha2e0:	data_out=16'h8a00;
17'ha2e1:	data_out=16'h8a00;
17'ha2e2:	data_out=16'h9e5;
17'ha2e3:	data_out=16'h9fe;
17'ha2e4:	data_out=16'h8934;
17'ha2e5:	data_out=16'h86dd;
17'ha2e6:	data_out=16'h883e;
17'ha2e7:	data_out=16'h89e8;
17'ha2e8:	data_out=16'h521;
17'ha2e9:	data_out=16'h878e;
17'ha2ea:	data_out=16'hbc;
17'ha2eb:	data_out=16'h8a00;
17'ha2ec:	data_out=16'h8a00;
17'ha2ed:	data_out=16'h9fe;
17'ha2ee:	data_out=16'hbd;
17'ha2ef:	data_out=16'h8a00;
17'ha2f0:	data_out=16'h154;
17'ha2f1:	data_out=16'h8d5;
17'ha2f2:	data_out=16'h8a00;
17'ha2f3:	data_out=16'h8a00;
17'ha2f4:	data_out=16'h8a00;
17'ha2f5:	data_out=16'h89fc;
17'ha2f6:	data_out=16'ha00;
17'ha2f7:	data_out=16'h89ef;
17'ha2f8:	data_out=16'h8990;
17'ha2f9:	data_out=16'h88bb;
17'ha2fa:	data_out=16'h9fa;
17'ha2fb:	data_out=16'h6e4;
17'ha2fc:	data_out=16'h8a00;
17'ha2fd:	data_out=16'h89ca;
17'ha2fe:	data_out=16'ha00;
17'ha2ff:	data_out=16'h8a00;
17'ha300:	data_out=16'h8a00;
17'ha301:	data_out=16'h87d4;
17'ha302:	data_out=16'h8a00;
17'ha303:	data_out=16'h8975;
17'ha304:	data_out=16'h8a00;
17'ha305:	data_out=16'h8a00;
17'ha306:	data_out=16'h9ff;
17'ha307:	data_out=16'h8a00;
17'ha308:	data_out=16'h89c5;
17'ha309:	data_out=16'h9e3;
17'ha30a:	data_out=16'h8904;
17'ha30b:	data_out=16'ha00;
17'ha30c:	data_out=16'h8911;
17'ha30d:	data_out=16'h8a00;
17'ha30e:	data_out=16'h388;
17'ha30f:	data_out=16'h8a00;
17'ha310:	data_out=16'h59a;
17'ha311:	data_out=16'ha00;
17'ha312:	data_out=16'h7bf;
17'ha313:	data_out=16'h84f6;
17'ha314:	data_out=16'h9ec;
17'ha315:	data_out=16'h8a00;
17'ha316:	data_out=16'h8a00;
17'ha317:	data_out=16'h9ef;
17'ha318:	data_out=16'h8a00;
17'ha319:	data_out=16'ha00;
17'ha31a:	data_out=16'h89e6;
17'ha31b:	data_out=16'h326;
17'ha31c:	data_out=16'h89ab;
17'ha31d:	data_out=16'ha00;
17'ha31e:	data_out=16'h877a;
17'ha31f:	data_out=16'h99d;
17'ha320:	data_out=16'h896c;
17'ha321:	data_out=16'h4d4;
17'ha322:	data_out=16'ha00;
17'ha323:	data_out=16'h8a00;
17'ha324:	data_out=16'h8a00;
17'ha325:	data_out=16'h89f9;
17'ha326:	data_out=16'h89d0;
17'ha327:	data_out=16'h8453;
17'ha328:	data_out=16'h788;
17'ha329:	data_out=16'h9de;
17'ha32a:	data_out=16'h8a00;
17'ha32b:	data_out=16'ha00;
17'ha32c:	data_out=16'h8a00;
17'ha32d:	data_out=16'ha00;
17'ha32e:	data_out=16'h9e4;
17'ha32f:	data_out=16'h83d0;
17'ha330:	data_out=16'h89d1;
17'ha331:	data_out=16'h891e;
17'ha332:	data_out=16'h89b5;
17'ha333:	data_out=16'ha00;
17'ha334:	data_out=16'h8439;
17'ha335:	data_out=16'h89b5;
17'ha336:	data_out=16'h885a;
17'ha337:	data_out=16'h897c;
17'ha338:	data_out=16'ha00;
17'ha339:	data_out=16'h9ff;
17'ha33a:	data_out=16'h886b;
17'ha33b:	data_out=16'h89ab;
17'ha33c:	data_out=16'h510;
17'ha33d:	data_out=16'h8a00;
17'ha33e:	data_out=16'h796;
17'ha33f:	data_out=16'h8a00;
17'ha340:	data_out=16'h899b;
17'ha341:	data_out=16'h8a00;
17'ha342:	data_out=16'h89d0;
17'ha343:	data_out=16'h89d8;
17'ha344:	data_out=16'h89c7;
17'ha345:	data_out=16'h8a00;
17'ha346:	data_out=16'ha00;
17'ha347:	data_out=16'h84b9;
17'ha348:	data_out=16'ha00;
17'ha349:	data_out=16'h89c8;
17'ha34a:	data_out=16'h3c9;
17'ha34b:	data_out=16'h8924;
17'ha34c:	data_out=16'h89ff;
17'ha34d:	data_out=16'ha00;
17'ha34e:	data_out=16'h98f;
17'ha34f:	data_out=16'h89e2;
17'ha350:	data_out=16'h8953;
17'ha351:	data_out=16'h89ff;
17'ha352:	data_out=16'h8a00;
17'ha353:	data_out=16'h9f5;
17'ha354:	data_out=16'h8655;
17'ha355:	data_out=16'h89fc;
17'ha356:	data_out=16'h8a00;
17'ha357:	data_out=16'h89fd;
17'ha358:	data_out=16'h89fe;
17'ha359:	data_out=16'h89b6;
17'ha35a:	data_out=16'h9b1;
17'ha35b:	data_out=16'h8964;
17'ha35c:	data_out=16'h8971;
17'ha35d:	data_out=16'h894b;
17'ha35e:	data_out=16'h8139;
17'ha35f:	data_out=16'h88ec;
17'ha360:	data_out=16'h9b7;
17'ha361:	data_out=16'h8a00;
17'ha362:	data_out=16'h9f1;
17'ha363:	data_out=16'h9ff;
17'ha364:	data_out=16'h9f9;
17'ha365:	data_out=16'ha00;
17'ha366:	data_out=16'h9f1;
17'ha367:	data_out=16'h8929;
17'ha368:	data_out=16'h617;
17'ha369:	data_out=16'h8a00;
17'ha36a:	data_out=16'h2cf;
17'ha36b:	data_out=16'h8984;
17'ha36c:	data_out=16'h8a00;
17'ha36d:	data_out=16'h9ff;
17'ha36e:	data_out=16'h2cf;
17'ha36f:	data_out=16'h89aa;
17'ha370:	data_out=16'h32c;
17'ha371:	data_out=16'h8a00;
17'ha372:	data_out=16'h89df;
17'ha373:	data_out=16'h8a00;
17'ha374:	data_out=16'h89db;
17'ha375:	data_out=16'h89f9;
17'ha376:	data_out=16'ha00;
17'ha377:	data_out=16'h89b5;
17'ha378:	data_out=16'h89cb;
17'ha379:	data_out=16'h8a00;
17'ha37a:	data_out=16'h9f7;
17'ha37b:	data_out=16'h79a;
17'ha37c:	data_out=16'h8a00;
17'ha37d:	data_out=16'h82dc;
17'ha37e:	data_out=16'ha00;
17'ha37f:	data_out=16'h8a00;
17'ha380:	data_out=16'h8a00;
17'ha381:	data_out=16'h879b;
17'ha382:	data_out=16'h8a00;
17'ha383:	data_out=16'h88a1;
17'ha384:	data_out=16'h8a00;
17'ha385:	data_out=16'h8a00;
17'ha386:	data_out=16'ha00;
17'ha387:	data_out=16'h8a00;
17'ha388:	data_out=16'h89df;
17'ha389:	data_out=16'h9fe;
17'ha38a:	data_out=16'h84ed;
17'ha38b:	data_out=16'ha00;
17'ha38c:	data_out=16'h8896;
17'ha38d:	data_out=16'h8a00;
17'ha38e:	data_out=16'h89fe;
17'ha38f:	data_out=16'h8a00;
17'ha390:	data_out=16'ha00;
17'ha391:	data_out=16'ha00;
17'ha392:	data_out=16'h8a00;
17'ha393:	data_out=16'h9a5;
17'ha394:	data_out=16'h8030;
17'ha395:	data_out=16'h8a00;
17'ha396:	data_out=16'h8a00;
17'ha397:	data_out=16'h9f2;
17'ha398:	data_out=16'h8a00;
17'ha399:	data_out=16'ha00;
17'ha39a:	data_out=16'h89ef;
17'ha39b:	data_out=16'h8948;
17'ha39c:	data_out=16'h89e6;
17'ha39d:	data_out=16'ha00;
17'ha39e:	data_out=16'h8848;
17'ha39f:	data_out=16'h97c;
17'ha3a0:	data_out=16'h89b4;
17'ha3a1:	data_out=16'h89fe;
17'ha3a2:	data_out=16'ha00;
17'ha3a3:	data_out=16'h38;
17'ha3a4:	data_out=16'h8078;
17'ha3a5:	data_out=16'h23b;
17'ha3a6:	data_out=16'h88bb;
17'ha3a7:	data_out=16'h8538;
17'ha3a8:	data_out=16'h8837;
17'ha3a9:	data_out=16'h9d8;
17'ha3aa:	data_out=16'h8a00;
17'ha3ab:	data_out=16'ha00;
17'ha3ac:	data_out=16'h8a00;
17'ha3ad:	data_out=16'ha00;
17'ha3ae:	data_out=16'ha00;
17'ha3af:	data_out=16'h86eb;
17'ha3b0:	data_out=16'h8704;
17'ha3b1:	data_out=16'h892d;
17'ha3b2:	data_out=16'h899c;
17'ha3b3:	data_out=16'h780;
17'ha3b4:	data_out=16'h9fd;
17'ha3b5:	data_out=16'h89b3;
17'ha3b6:	data_out=16'h89d9;
17'ha3b7:	data_out=16'h89fc;
17'ha3b8:	data_out=16'ha00;
17'ha3b9:	data_out=16'h8563;
17'ha3ba:	data_out=16'h84c;
17'ha3bb:	data_out=16'h8998;
17'ha3bc:	data_out=16'h9fc;
17'ha3bd:	data_out=16'h89f3;
17'ha3be:	data_out=16'h881e;
17'ha3bf:	data_out=16'h8a00;
17'ha3c0:	data_out=16'h89a2;
17'ha3c1:	data_out=16'h8a00;
17'ha3c2:	data_out=16'h8967;
17'ha3c3:	data_out=16'h89fd;
17'ha3c4:	data_out=16'h89cb;
17'ha3c5:	data_out=16'h8a00;
17'ha3c6:	data_out=16'ha00;
17'ha3c7:	data_out=16'h8381;
17'ha3c8:	data_out=16'ha00;
17'ha3c9:	data_out=16'h83e6;
17'ha3ca:	data_out=16'h87ee;
17'ha3cb:	data_out=16'h87cd;
17'ha3cc:	data_out=16'h89fe;
17'ha3cd:	data_out=16'ha00;
17'ha3ce:	data_out=16'h6c8;
17'ha3cf:	data_out=16'h86a2;
17'ha3d0:	data_out=16'h8958;
17'ha3d1:	data_out=16'h8a00;
17'ha3d2:	data_out=16'h8a00;
17'ha3d3:	data_out=16'h9fe;
17'ha3d4:	data_out=16'h8810;
17'ha3d5:	data_out=16'h8668;
17'ha3d6:	data_out=16'h8a00;
17'ha3d7:	data_out=16'h89fb;
17'ha3d8:	data_out=16'h8a00;
17'ha3d9:	data_out=16'h899b;
17'ha3da:	data_out=16'h4ec;
17'ha3db:	data_out=16'h890d;
17'ha3dc:	data_out=16'h89cb;
17'ha3dd:	data_out=16'h89ce;
17'ha3de:	data_out=16'h8517;
17'ha3df:	data_out=16'h896b;
17'ha3e0:	data_out=16'h9c5;
17'ha3e1:	data_out=16'h89fa;
17'ha3e2:	data_out=16'h9fa;
17'ha3e3:	data_out=16'h9fe;
17'ha3e4:	data_out=16'h9fe;
17'ha3e5:	data_out=16'ha00;
17'ha3e6:	data_out=16'h9fd;
17'ha3e7:	data_out=16'h9eb;
17'ha3e8:	data_out=16'h89f7;
17'ha3e9:	data_out=16'h8a00;
17'ha3ea:	data_out=16'h89fe;
17'ha3eb:	data_out=16'h899f;
17'ha3ec:	data_out=16'h8a00;
17'ha3ed:	data_out=16'h9ff;
17'ha3ee:	data_out=16'h89fe;
17'ha3ef:	data_out=16'h89c1;
17'ha3f0:	data_out=16'h89fe;
17'ha3f1:	data_out=16'h8a00;
17'ha3f2:	data_out=16'h89c5;
17'ha3f3:	data_out=16'h89e9;
17'ha3f4:	data_out=16'h87a4;
17'ha3f5:	data_out=16'h89fe;
17'ha3f6:	data_out=16'ha00;
17'ha3f7:	data_out=16'h896a;
17'ha3f8:	data_out=16'h89f4;
17'ha3f9:	data_out=16'h8a00;
17'ha3fa:	data_out=16'h81bf;
17'ha3fb:	data_out=16'h881a;
17'ha3fc:	data_out=16'h8a00;
17'ha3fd:	data_out=16'h89fc;
17'ha3fe:	data_out=16'ha00;
17'ha3ff:	data_out=16'h8a00;
17'ha400:	data_out=16'h8a00;
17'ha401:	data_out=16'h88de;
17'ha402:	data_out=16'h8a00;
17'ha403:	data_out=16'h86c6;
17'ha404:	data_out=16'h8a00;
17'ha405:	data_out=16'h8a00;
17'ha406:	data_out=16'ha00;
17'ha407:	data_out=16'h871a;
17'ha408:	data_out=16'h89d7;
17'ha409:	data_out=16'ha00;
17'ha40a:	data_out=16'h897c;
17'ha40b:	data_out=16'ha00;
17'ha40c:	data_out=16'h82bf;
17'ha40d:	data_out=16'h8a00;
17'ha40e:	data_out=16'h8a00;
17'ha40f:	data_out=16'h8a00;
17'ha410:	data_out=16'h9f8;
17'ha411:	data_out=16'h8084;
17'ha412:	data_out=16'h8a00;
17'ha413:	data_out=16'h9cf;
17'ha414:	data_out=16'h8045;
17'ha415:	data_out=16'h8a00;
17'ha416:	data_out=16'h8a00;
17'ha417:	data_out=16'ha00;
17'ha418:	data_out=16'h8a00;
17'ha419:	data_out=16'ha00;
17'ha41a:	data_out=16'h8a00;
17'ha41b:	data_out=16'h87e5;
17'ha41c:	data_out=16'h89e3;
17'ha41d:	data_out=16'ha00;
17'ha41e:	data_out=16'h897a;
17'ha41f:	data_out=16'h82fb;
17'ha420:	data_out=16'h89f7;
17'ha421:	data_out=16'h89ff;
17'ha422:	data_out=16'ha00;
17'ha423:	data_out=16'h780;
17'ha424:	data_out=16'h6f9;
17'ha425:	data_out=16'h5b4;
17'ha426:	data_out=16'h9f7;
17'ha427:	data_out=16'h8996;
17'ha428:	data_out=16'h89ff;
17'ha429:	data_out=16'h9ea;
17'ha42a:	data_out=16'h8993;
17'ha42b:	data_out=16'ha00;
17'ha42c:	data_out=16'h8a00;
17'ha42d:	data_out=16'ha00;
17'ha42e:	data_out=16'ha00;
17'ha42f:	data_out=16'h8911;
17'ha430:	data_out=16'h894f;
17'ha431:	data_out=16'h89c4;
17'ha432:	data_out=16'h8994;
17'ha433:	data_out=16'h8658;
17'ha434:	data_out=16'h9fc;
17'ha435:	data_out=16'h89ef;
17'ha436:	data_out=16'h89d5;
17'ha437:	data_out=16'h89f2;
17'ha438:	data_out=16'ha00;
17'ha439:	data_out=16'h8950;
17'ha43a:	data_out=16'h2c6;
17'ha43b:	data_out=16'h89df;
17'ha43c:	data_out=16'ha00;
17'ha43d:	data_out=16'h8a00;
17'ha43e:	data_out=16'h89ff;
17'ha43f:	data_out=16'h8a00;
17'ha440:	data_out=16'h89df;
17'ha441:	data_out=16'h8a00;
17'ha442:	data_out=16'h9ff;
17'ha443:	data_out=16'h8793;
17'ha444:	data_out=16'h8a00;
17'ha445:	data_out=16'h8a00;
17'ha446:	data_out=16'ha00;
17'ha447:	data_out=16'h86ff;
17'ha448:	data_out=16'ha00;
17'ha449:	data_out=16'h25e;
17'ha44a:	data_out=16'h8980;
17'ha44b:	data_out=16'h9ff;
17'ha44c:	data_out=16'h436;
17'ha44d:	data_out=16'ha00;
17'ha44e:	data_out=16'h9f9;
17'ha44f:	data_out=16'h8411;
17'ha450:	data_out=16'h89cf;
17'ha451:	data_out=16'h8a00;
17'ha452:	data_out=16'h89fe;
17'ha453:	data_out=16'h5dc;
17'ha454:	data_out=16'h89b0;
17'ha455:	data_out=16'h6cd;
17'ha456:	data_out=16'h8a00;
17'ha457:	data_out=16'h8a00;
17'ha458:	data_out=16'h8a00;
17'ha459:	data_out=16'h89d9;
17'ha45a:	data_out=16'h9c2;
17'ha45b:	data_out=16'h89ed;
17'ha45c:	data_out=16'h89d6;
17'ha45d:	data_out=16'h89d0;
17'ha45e:	data_out=16'h8775;
17'ha45f:	data_out=16'h89ee;
17'ha460:	data_out=16'ha00;
17'ha461:	data_out=16'h89fe;
17'ha462:	data_out=16'ha00;
17'ha463:	data_out=16'h8198;
17'ha464:	data_out=16'ha00;
17'ha465:	data_out=16'ha00;
17'ha466:	data_out=16'ha00;
17'ha467:	data_out=16'ha00;
17'ha468:	data_out=16'h89ff;
17'ha469:	data_out=16'h89f4;
17'ha46a:	data_out=16'h8a00;
17'ha46b:	data_out=16'h8a00;
17'ha46c:	data_out=16'h8a00;
17'ha46d:	data_out=16'h82d8;
17'ha46e:	data_out=16'h8a00;
17'ha46f:	data_out=16'h89ca;
17'ha470:	data_out=16'h8a00;
17'ha471:	data_out=16'h8a00;
17'ha472:	data_out=16'h89f3;
17'ha473:	data_out=16'h89e9;
17'ha474:	data_out=16'h895b;
17'ha475:	data_out=16'h8a00;
17'ha476:	data_out=16'ha00;
17'ha477:	data_out=16'h891e;
17'ha478:	data_out=16'h89ff;
17'ha479:	data_out=16'h8a00;
17'ha47a:	data_out=16'h8418;
17'ha47b:	data_out=16'h89ff;
17'ha47c:	data_out=16'h8a00;
17'ha47d:	data_out=16'h8a00;
17'ha47e:	data_out=16'ha00;
17'ha47f:	data_out=16'h8a00;
17'ha480:	data_out=16'h8a00;
17'ha481:	data_out=16'h89d8;
17'ha482:	data_out=16'h8a00;
17'ha483:	data_out=16'h88b6;
17'ha484:	data_out=16'h8a00;
17'ha485:	data_out=16'h8a00;
17'ha486:	data_out=16'ha00;
17'ha487:	data_out=16'h73f;
17'ha488:	data_out=16'h8a00;
17'ha489:	data_out=16'ha00;
17'ha48a:	data_out=16'h89af;
17'ha48b:	data_out=16'ha00;
17'ha48c:	data_out=16'ha00;
17'ha48d:	data_out=16'h8a00;
17'ha48e:	data_out=16'h8a00;
17'ha48f:	data_out=16'h89fb;
17'ha490:	data_out=16'h820e;
17'ha491:	data_out=16'h89e0;
17'ha492:	data_out=16'h8a00;
17'ha493:	data_out=16'h9ec;
17'ha494:	data_out=16'h895a;
17'ha495:	data_out=16'h8a00;
17'ha496:	data_out=16'h8a00;
17'ha497:	data_out=16'h8285;
17'ha498:	data_out=16'h8a00;
17'ha499:	data_out=16'ha00;
17'ha49a:	data_out=16'h8a00;
17'ha49b:	data_out=16'h89e7;
17'ha49c:	data_out=16'h8a00;
17'ha49d:	data_out=16'h823c;
17'ha49e:	data_out=16'h89fe;
17'ha49f:	data_out=16'h89f6;
17'ha4a0:	data_out=16'h8a00;
17'ha4a1:	data_out=16'h8a00;
17'ha4a2:	data_out=16'ha00;
17'ha4a3:	data_out=16'ha00;
17'ha4a4:	data_out=16'h9ff;
17'ha4a5:	data_out=16'h85a;
17'ha4a6:	data_out=16'ha00;
17'ha4a7:	data_out=16'h89f3;
17'ha4a8:	data_out=16'h8a00;
17'ha4a9:	data_out=16'h9d3;
17'ha4aa:	data_out=16'h892f;
17'ha4ab:	data_out=16'ha00;
17'ha4ac:	data_out=16'h8a00;
17'ha4ad:	data_out=16'ha00;
17'ha4ae:	data_out=16'ha00;
17'ha4af:	data_out=16'h89ed;
17'ha4b0:	data_out=16'h8970;
17'ha4b1:	data_out=16'h89fd;
17'ha4b2:	data_out=16'h89b3;
17'ha4b3:	data_out=16'h89fa;
17'ha4b4:	data_out=16'h9a8;
17'ha4b5:	data_out=16'h8a00;
17'ha4b6:	data_out=16'h89fa;
17'ha4b7:	data_out=16'h8a00;
17'ha4b8:	data_out=16'h96a;
17'ha4b9:	data_out=16'h89fd;
17'ha4ba:	data_out=16'h30e;
17'ha4bb:	data_out=16'h89ef;
17'ha4bc:	data_out=16'h9eb;
17'ha4bd:	data_out=16'h8a00;
17'ha4be:	data_out=16'h8a00;
17'ha4bf:	data_out=16'h8a00;
17'ha4c0:	data_out=16'h8a00;
17'ha4c1:	data_out=16'h8a00;
17'ha4c2:	data_out=16'ha00;
17'ha4c3:	data_out=16'h89fe;
17'ha4c4:	data_out=16'h8a00;
17'ha4c5:	data_out=16'h8a00;
17'ha4c6:	data_out=16'ha00;
17'ha4c7:	data_out=16'h8125;
17'ha4c8:	data_out=16'ha00;
17'ha4c9:	data_out=16'h656;
17'ha4ca:	data_out=16'h89ac;
17'ha4cb:	data_out=16'ha00;
17'ha4cc:	data_out=16'h9e1;
17'ha4cd:	data_out=16'ha00;
17'ha4ce:	data_out=16'h464;
17'ha4cf:	data_out=16'ha00;
17'ha4d0:	data_out=16'h89fd;
17'ha4d1:	data_out=16'h8a00;
17'ha4d2:	data_out=16'h35d;
17'ha4d3:	data_out=16'h89d6;
17'ha4d4:	data_out=16'h8a00;
17'ha4d5:	data_out=16'h89f6;
17'ha4d6:	data_out=16'h8a00;
17'ha4d7:	data_out=16'h8a00;
17'ha4d8:	data_out=16'h8a00;
17'ha4d9:	data_out=16'h8a00;
17'ha4da:	data_out=16'h89f0;
17'ha4db:	data_out=16'h8a00;
17'ha4dc:	data_out=16'h8a00;
17'ha4dd:	data_out=16'h89f4;
17'ha4de:	data_out=16'h899c;
17'ha4df:	data_out=16'h89fe;
17'ha4e0:	data_out=16'ha00;
17'ha4e1:	data_out=16'h8a00;
17'ha4e2:	data_out=16'ha00;
17'ha4e3:	data_out=16'h89f9;
17'ha4e4:	data_out=16'ha00;
17'ha4e5:	data_out=16'h9fc;
17'ha4e6:	data_out=16'h9ff;
17'ha4e7:	data_out=16'h9fd;
17'ha4e8:	data_out=16'h8a00;
17'ha4e9:	data_out=16'h8a00;
17'ha4ea:	data_out=16'h8a00;
17'ha4eb:	data_out=16'h8a00;
17'ha4ec:	data_out=16'h8a00;
17'ha4ed:	data_out=16'h89f9;
17'ha4ee:	data_out=16'h8a00;
17'ha4ef:	data_out=16'h89f3;
17'ha4f0:	data_out=16'h8a00;
17'ha4f1:	data_out=16'h8a00;
17'ha4f2:	data_out=16'h8a00;
17'ha4f3:	data_out=16'h8a00;
17'ha4f4:	data_out=16'h8979;
17'ha4f5:	data_out=16'h8a00;
17'ha4f6:	data_out=16'ha00;
17'ha4f7:	data_out=16'h8946;
17'ha4f8:	data_out=16'h8397;
17'ha4f9:	data_out=16'h8a00;
17'ha4fa:	data_out=16'h89bd;
17'ha4fb:	data_out=16'h8a00;
17'ha4fc:	data_out=16'h8a00;
17'ha4fd:	data_out=16'h8a00;
17'ha4fe:	data_out=16'ha00;
17'ha4ff:	data_out=16'h8a00;
17'ha500:	data_out=16'h8a00;
17'ha501:	data_out=16'h884b;
17'ha502:	data_out=16'h8a00;
17'ha503:	data_out=16'h89cf;
17'ha504:	data_out=16'h8a00;
17'ha505:	data_out=16'h8a00;
17'ha506:	data_out=16'ha00;
17'ha507:	data_out=16'h8386;
17'ha508:	data_out=16'h8a00;
17'ha509:	data_out=16'h3e8;
17'ha50a:	data_out=16'h620;
17'ha50b:	data_out=16'ha00;
17'ha50c:	data_out=16'ha00;
17'ha50d:	data_out=16'h8a00;
17'ha50e:	data_out=16'h8a00;
17'ha50f:	data_out=16'h89fa;
17'ha510:	data_out=16'h89fa;
17'ha511:	data_out=16'h89fe;
17'ha512:	data_out=16'h8a00;
17'ha513:	data_out=16'h9d0;
17'ha514:	data_out=16'h89ff;
17'ha515:	data_out=16'h8a00;
17'ha516:	data_out=16'h8a00;
17'ha517:	data_out=16'h895f;
17'ha518:	data_out=16'h8a00;
17'ha519:	data_out=16'ha00;
17'ha51a:	data_out=16'h8a00;
17'ha51b:	data_out=16'h89ff;
17'ha51c:	data_out=16'h8a00;
17'ha51d:	data_out=16'h50;
17'ha51e:	data_out=16'h8a00;
17'ha51f:	data_out=16'h8a00;
17'ha520:	data_out=16'h8a00;
17'ha521:	data_out=16'h8a00;
17'ha522:	data_out=16'h9f5;
17'ha523:	data_out=16'h9ff;
17'ha524:	data_out=16'h9ff;
17'ha525:	data_out=16'h4e2;
17'ha526:	data_out=16'ha00;
17'ha527:	data_out=16'h8a00;
17'ha528:	data_out=16'h8a00;
17'ha529:	data_out=16'h9e6;
17'ha52a:	data_out=16'h8931;
17'ha52b:	data_out=16'h886b;
17'ha52c:	data_out=16'h8a00;
17'ha52d:	data_out=16'ha00;
17'ha52e:	data_out=16'h61e;
17'ha52f:	data_out=16'h8a00;
17'ha530:	data_out=16'h94d;
17'ha531:	data_out=16'h8a00;
17'ha532:	data_out=16'h8da;
17'ha533:	data_out=16'h8a00;
17'ha534:	data_out=16'ha00;
17'ha535:	data_out=16'h8a00;
17'ha536:	data_out=16'h8a00;
17'ha537:	data_out=16'h8a00;
17'ha538:	data_out=16'h6b7;
17'ha539:	data_out=16'h8a00;
17'ha53a:	data_out=16'h89e3;
17'ha53b:	data_out=16'h8a00;
17'ha53c:	data_out=16'h9f3;
17'ha53d:	data_out=16'h8a00;
17'ha53e:	data_out=16'h8a00;
17'ha53f:	data_out=16'h8a00;
17'ha540:	data_out=16'h8a00;
17'ha541:	data_out=16'h8a00;
17'ha542:	data_out=16'ha00;
17'ha543:	data_out=16'h8a00;
17'ha544:	data_out=16'h8a00;
17'ha545:	data_out=16'h8a00;
17'ha546:	data_out=16'ha00;
17'ha547:	data_out=16'h89c6;
17'ha548:	data_out=16'h79a;
17'ha549:	data_out=16'h26b;
17'ha54a:	data_out=16'h89d7;
17'ha54b:	data_out=16'ha00;
17'ha54c:	data_out=16'ha00;
17'ha54d:	data_out=16'h9f6;
17'ha54e:	data_out=16'h8541;
17'ha54f:	data_out=16'ha00;
17'ha550:	data_out=16'h8a00;
17'ha551:	data_out=16'h8a00;
17'ha552:	data_out=16'h9fe;
17'ha553:	data_out=16'h8a00;
17'ha554:	data_out=16'h8a00;
17'ha555:	data_out=16'h8a00;
17'ha556:	data_out=16'h8a00;
17'ha557:	data_out=16'h8a00;
17'ha558:	data_out=16'h8a00;
17'ha559:	data_out=16'h8a00;
17'ha55a:	data_out=16'h8a00;
17'ha55b:	data_out=16'h8a00;
17'ha55c:	data_out=16'h8a00;
17'ha55d:	data_out=16'h8a00;
17'ha55e:	data_out=16'h89f0;
17'ha55f:	data_out=16'h8a00;
17'ha560:	data_out=16'ha00;
17'ha561:	data_out=16'h8a00;
17'ha562:	data_out=16'ha00;
17'ha563:	data_out=16'h8a00;
17'ha564:	data_out=16'ha00;
17'ha565:	data_out=16'h43a;
17'ha566:	data_out=16'h8592;
17'ha567:	data_out=16'h9e7;
17'ha568:	data_out=16'h8a00;
17'ha569:	data_out=16'h8a00;
17'ha56a:	data_out=16'h8a00;
17'ha56b:	data_out=16'h8a00;
17'ha56c:	data_out=16'h89f3;
17'ha56d:	data_out=16'h8a00;
17'ha56e:	data_out=16'h8a00;
17'ha56f:	data_out=16'h8a00;
17'ha570:	data_out=16'h8a00;
17'ha571:	data_out=16'h89f9;
17'ha572:	data_out=16'h8a00;
17'ha573:	data_out=16'h89f0;
17'ha574:	data_out=16'h984;
17'ha575:	data_out=16'h8a00;
17'ha576:	data_out=16'ha00;
17'ha577:	data_out=16'h89fc;
17'ha578:	data_out=16'h554;
17'ha579:	data_out=16'h8a00;
17'ha57a:	data_out=16'h8a00;
17'ha57b:	data_out=16'h8a00;
17'ha57c:	data_out=16'h8a00;
17'ha57d:	data_out=16'h8a00;
17'ha57e:	data_out=16'ha00;
17'ha57f:	data_out=16'h8a00;
17'ha580:	data_out=16'h89fd;
17'ha581:	data_out=16'h8188;
17'ha582:	data_out=16'h8a00;
17'ha583:	data_out=16'h8a00;
17'ha584:	data_out=16'h89ff;
17'ha585:	data_out=16'h8a00;
17'ha586:	data_out=16'ha00;
17'ha587:	data_out=16'h881a;
17'ha588:	data_out=16'h8a00;
17'ha589:	data_out=16'h877e;
17'ha58a:	data_out=16'ha00;
17'ha58b:	data_out=16'h4fe;
17'ha58c:	data_out=16'ha00;
17'ha58d:	data_out=16'h8a00;
17'ha58e:	data_out=16'h896e;
17'ha58f:	data_out=16'h89fd;
17'ha590:	data_out=16'h8a00;
17'ha591:	data_out=16'h89fd;
17'ha592:	data_out=16'h8a00;
17'ha593:	data_out=16'hcd;
17'ha594:	data_out=16'h8a00;
17'ha595:	data_out=16'h8a00;
17'ha596:	data_out=16'h8a00;
17'ha597:	data_out=16'h89fb;
17'ha598:	data_out=16'h8a00;
17'ha599:	data_out=16'h9f8;
17'ha59a:	data_out=16'h8a00;
17'ha59b:	data_out=16'h8a00;
17'ha59c:	data_out=16'h8a00;
17'ha59d:	data_out=16'h8169;
17'ha59e:	data_out=16'h8a00;
17'ha59f:	data_out=16'h8a00;
17'ha5a0:	data_out=16'h8a00;
17'ha5a1:	data_out=16'h89d4;
17'ha5a2:	data_out=16'h9eb;
17'ha5a3:	data_out=16'ha00;
17'ha5a4:	data_out=16'ha00;
17'ha5a5:	data_out=16'h89b;
17'ha5a6:	data_out=16'ha00;
17'ha5a7:	data_out=16'h8a00;
17'ha5a8:	data_out=16'h89fe;
17'ha5a9:	data_out=16'h867b;
17'ha5aa:	data_out=16'h89d2;
17'ha5ab:	data_out=16'h8a00;
17'ha5ac:	data_out=16'h8a00;
17'ha5ad:	data_out=16'ha00;
17'ha5ae:	data_out=16'h8934;
17'ha5af:	data_out=16'h8a00;
17'ha5b0:	data_out=16'ha00;
17'ha5b1:	data_out=16'h89fe;
17'ha5b2:	data_out=16'ha00;
17'ha5b3:	data_out=16'h8a00;
17'ha5b4:	data_out=16'ha00;
17'ha5b5:	data_out=16'h89ff;
17'ha5b6:	data_out=16'h8a00;
17'ha5b7:	data_out=16'h8a00;
17'ha5b8:	data_out=16'h3f3;
17'ha5b9:	data_out=16'h8a00;
17'ha5ba:	data_out=16'h89ff;
17'ha5bb:	data_out=16'h7b3;
17'ha5bc:	data_out=16'h1bb;
17'ha5bd:	data_out=16'h8a00;
17'ha5be:	data_out=16'h89fe;
17'ha5bf:	data_out=16'h8a00;
17'ha5c0:	data_out=16'h89e0;
17'ha5c1:	data_out=16'h8a00;
17'ha5c2:	data_out=16'ha00;
17'ha5c3:	data_out=16'h8a00;
17'ha5c4:	data_out=16'h8a00;
17'ha5c5:	data_out=16'h8a00;
17'ha5c6:	data_out=16'ha00;
17'ha5c7:	data_out=16'h89f3;
17'ha5c8:	data_out=16'h89b5;
17'ha5c9:	data_out=16'h7f8;
17'ha5ca:	data_out=16'h8a00;
17'ha5cb:	data_out=16'ha00;
17'ha5cc:	data_out=16'ha00;
17'ha5cd:	data_out=16'h3c2;
17'ha5ce:	data_out=16'h89f5;
17'ha5cf:	data_out=16'ha00;
17'ha5d0:	data_out=16'h8a00;
17'ha5d1:	data_out=16'h8a00;
17'ha5d2:	data_out=16'ha00;
17'ha5d3:	data_out=16'h8a00;
17'ha5d4:	data_out=16'h8a00;
17'ha5d5:	data_out=16'h8a00;
17'ha5d6:	data_out=16'h89fa;
17'ha5d7:	data_out=16'h8a00;
17'ha5d8:	data_out=16'h8a00;
17'ha5d9:	data_out=16'h89d8;
17'ha5da:	data_out=16'h8a00;
17'ha5db:	data_out=16'h89ff;
17'ha5dc:	data_out=16'h8a00;
17'ha5dd:	data_out=16'h89fb;
17'ha5de:	data_out=16'h89fd;
17'ha5df:	data_out=16'h8a00;
17'ha5e0:	data_out=16'ha00;
17'ha5e1:	data_out=16'h8932;
17'ha5e2:	data_out=16'h88ab;
17'ha5e3:	data_out=16'h8a00;
17'ha5e4:	data_out=16'h9f6;
17'ha5e5:	data_out=16'h9ff;
17'ha5e6:	data_out=16'h8a00;
17'ha5e7:	data_out=16'h89ff;
17'ha5e8:	data_out=16'h89fc;
17'ha5e9:	data_out=16'h8a00;
17'ha5ea:	data_out=16'h89a1;
17'ha5eb:	data_out=16'h8a00;
17'ha5ec:	data_out=16'h89f5;
17'ha5ed:	data_out=16'h8a00;
17'ha5ee:	data_out=16'h899a;
17'ha5ef:	data_out=16'h6d9;
17'ha5f0:	data_out=16'h8969;
17'ha5f1:	data_out=16'h89fd;
17'ha5f2:	data_out=16'h89f6;
17'ha5f3:	data_out=16'h95a;
17'ha5f4:	data_out=16'ha00;
17'ha5f5:	data_out=16'h8a00;
17'ha5f6:	data_out=16'h89ff;
17'ha5f7:	data_out=16'h89f6;
17'ha5f8:	data_out=16'h9fe;
17'ha5f9:	data_out=16'h8a00;
17'ha5fa:	data_out=16'h8a00;
17'ha5fb:	data_out=16'h89fe;
17'ha5fc:	data_out=16'h8a00;
17'ha5fd:	data_out=16'h8a00;
17'ha5fe:	data_out=16'h9e4;
17'ha5ff:	data_out=16'h8a00;
17'ha600:	data_out=16'h89f4;
17'ha601:	data_out=16'h1db;
17'ha602:	data_out=16'h89fe;
17'ha603:	data_out=16'h8a00;
17'ha604:	data_out=16'h9e9;
17'ha605:	data_out=16'h89f4;
17'ha606:	data_out=16'h8079;
17'ha607:	data_out=16'h89f9;
17'ha608:	data_out=16'h8a00;
17'ha609:	data_out=16'h89ed;
17'ha60a:	data_out=16'ha00;
17'ha60b:	data_out=16'h89fa;
17'ha60c:	data_out=16'h89f8;
17'ha60d:	data_out=16'h8a00;
17'ha60e:	data_out=16'ha00;
17'ha60f:	data_out=16'h8a00;
17'ha610:	data_out=16'h8a00;
17'ha611:	data_out=16'h386;
17'ha612:	data_out=16'h8a00;
17'ha613:	data_out=16'h89ff;
17'ha614:	data_out=16'h8a00;
17'ha615:	data_out=16'h89ff;
17'ha616:	data_out=16'h8a00;
17'ha617:	data_out=16'h8a00;
17'ha618:	data_out=16'h8a00;
17'ha619:	data_out=16'h89f7;
17'ha61a:	data_out=16'h9ff;
17'ha61b:	data_out=16'h8a00;
17'ha61c:	data_out=16'h8a00;
17'ha61d:	data_out=16'h8688;
17'ha61e:	data_out=16'h8a00;
17'ha61f:	data_out=16'h8a00;
17'ha620:	data_out=16'h8a00;
17'ha621:	data_out=16'ha00;
17'ha622:	data_out=16'h89ea;
17'ha623:	data_out=16'ha00;
17'ha624:	data_out=16'ha00;
17'ha625:	data_out=16'h85ab;
17'ha626:	data_out=16'h803c;
17'ha627:	data_out=16'h89ff;
17'ha628:	data_out=16'h9ff;
17'ha629:	data_out=16'h89f1;
17'ha62a:	data_out=16'h89fb;
17'ha62b:	data_out=16'h8a00;
17'ha62c:	data_out=16'h8a00;
17'ha62d:	data_out=16'ha00;
17'ha62e:	data_out=16'h89f8;
17'ha62f:	data_out=16'h8a00;
17'ha630:	data_out=16'ha00;
17'ha631:	data_out=16'h600;
17'ha632:	data_out=16'ha00;
17'ha633:	data_out=16'h8a00;
17'ha634:	data_out=16'h9fb;
17'ha635:	data_out=16'h89f2;
17'ha636:	data_out=16'h8a00;
17'ha637:	data_out=16'h8a00;
17'ha638:	data_out=16'h712;
17'ha639:	data_out=16'h8a00;
17'ha63a:	data_out=16'h8a00;
17'ha63b:	data_out=16'h9f5;
17'ha63c:	data_out=16'h85b6;
17'ha63d:	data_out=16'h8a00;
17'ha63e:	data_out=16'h9ff;
17'ha63f:	data_out=16'h89f2;
17'ha640:	data_out=16'h83de;
17'ha641:	data_out=16'h89fd;
17'ha642:	data_out=16'ha00;
17'ha643:	data_out=16'h8a00;
17'ha644:	data_out=16'h89fc;
17'ha645:	data_out=16'h89ff;
17'ha646:	data_out=16'h9f7;
17'ha647:	data_out=16'h8a00;
17'ha648:	data_out=16'h89f7;
17'ha649:	data_out=16'h86c9;
17'ha64a:	data_out=16'h8a00;
17'ha64b:	data_out=16'ha00;
17'ha64c:	data_out=16'ha00;
17'ha64d:	data_out=16'h89f0;
17'ha64e:	data_out=16'h89f4;
17'ha64f:	data_out=16'h55a;
17'ha650:	data_out=16'h8a00;
17'ha651:	data_out=16'h8a00;
17'ha652:	data_out=16'ha00;
17'ha653:	data_out=16'h8a00;
17'ha654:	data_out=16'h8a00;
17'ha655:	data_out=16'h8a00;
17'ha656:	data_out=16'h817c;
17'ha657:	data_out=16'h876b;
17'ha658:	data_out=16'h8a00;
17'ha659:	data_out=16'ha00;
17'ha65a:	data_out=16'h8a00;
17'ha65b:	data_out=16'h8ac;
17'ha65c:	data_out=16'h8a00;
17'ha65d:	data_out=16'h89fe;
17'ha65e:	data_out=16'h8a00;
17'ha65f:	data_out=16'h8a00;
17'ha660:	data_out=16'h9f6;
17'ha661:	data_out=16'h4c9;
17'ha662:	data_out=16'h8a00;
17'ha663:	data_out=16'h8a00;
17'ha664:	data_out=16'h838e;
17'ha665:	data_out=16'h89ae;
17'ha666:	data_out=16'h8a00;
17'ha667:	data_out=16'h8a00;
17'ha668:	data_out=16'ha00;
17'ha669:	data_out=16'h8a00;
17'ha66a:	data_out=16'ha00;
17'ha66b:	data_out=16'h8a00;
17'ha66c:	data_out=16'h8d5;
17'ha66d:	data_out=16'h8a00;
17'ha66e:	data_out=16'ha00;
17'ha66f:	data_out=16'h6ea;
17'ha670:	data_out=16'ha00;
17'ha671:	data_out=16'h8a00;
17'ha672:	data_out=16'h9fd;
17'ha673:	data_out=16'ha00;
17'ha674:	data_out=16'ha00;
17'ha675:	data_out=16'h9f0;
17'ha676:	data_out=16'h8a00;
17'ha677:	data_out=16'h8a00;
17'ha678:	data_out=16'h82c3;
17'ha679:	data_out=16'h89ff;
17'ha67a:	data_out=16'h8a00;
17'ha67b:	data_out=16'h9ff;
17'ha67c:	data_out=16'h8a00;
17'ha67d:	data_out=16'h8a00;
17'ha67e:	data_out=16'h89e2;
17'ha67f:	data_out=16'h8a00;
17'ha680:	data_out=16'ha00;
17'ha681:	data_out=16'h9fe;
17'ha682:	data_out=16'h5c5;
17'ha683:	data_out=16'h8a00;
17'ha684:	data_out=16'ha00;
17'ha685:	data_out=16'ha00;
17'ha686:	data_out=16'h8a00;
17'ha687:	data_out=16'h8a00;
17'ha688:	data_out=16'h98b;
17'ha689:	data_out=16'h8a00;
17'ha68a:	data_out=16'ha00;
17'ha68b:	data_out=16'h8a00;
17'ha68c:	data_out=16'h8a00;
17'ha68d:	data_out=16'h89f8;
17'ha68e:	data_out=16'ha00;
17'ha68f:	data_out=16'h89fd;
17'ha690:	data_out=16'h8a00;
17'ha691:	data_out=16'h98f;
17'ha692:	data_out=16'h89fb;
17'ha693:	data_out=16'h89fd;
17'ha694:	data_out=16'h8a00;
17'ha695:	data_out=16'ha00;
17'ha696:	data_out=16'h844e;
17'ha697:	data_out=16'h8a00;
17'ha698:	data_out=16'h523;
17'ha699:	data_out=16'h8a00;
17'ha69a:	data_out=16'ha00;
17'ha69b:	data_out=16'h8a00;
17'ha69c:	data_out=16'h972;
17'ha69d:	data_out=16'h87ba;
17'ha69e:	data_out=16'h8a00;
17'ha69f:	data_out=16'h8a00;
17'ha6a0:	data_out=16'h8761;
17'ha6a1:	data_out=16'ha00;
17'ha6a2:	data_out=16'h8a00;
17'ha6a3:	data_out=16'ha00;
17'ha6a4:	data_out=16'ha00;
17'ha6a5:	data_out=16'h89f1;
17'ha6a6:	data_out=16'h89f8;
17'ha6a7:	data_out=16'h89d7;
17'ha6a8:	data_out=16'ha00;
17'ha6a9:	data_out=16'h8a00;
17'ha6aa:	data_out=16'h89fe;
17'ha6ab:	data_out=16'h8a00;
17'ha6ac:	data_out=16'h8113;
17'ha6ad:	data_out=16'h89aa;
17'ha6ae:	data_out=16'h8a00;
17'ha6af:	data_out=16'h8a00;
17'ha6b0:	data_out=16'ha00;
17'ha6b1:	data_out=16'h89bb;
17'ha6b2:	data_out=16'ha00;
17'ha6b3:	data_out=16'h8a00;
17'ha6b4:	data_out=16'h8258;
17'ha6b5:	data_out=16'ha00;
17'ha6b6:	data_out=16'h89e4;
17'ha6b7:	data_out=16'h80b1;
17'ha6b8:	data_out=16'h9fb;
17'ha6b9:	data_out=16'h8a00;
17'ha6ba:	data_out=16'h8a00;
17'ha6bb:	data_out=16'ha00;
17'ha6bc:	data_out=16'h80ce;
17'ha6bd:	data_out=16'h44c;
17'ha6be:	data_out=16'ha00;
17'ha6bf:	data_out=16'ha00;
17'ha6c0:	data_out=16'h87c7;
17'ha6c1:	data_out=16'h891e;
17'ha6c2:	data_out=16'h89f9;
17'ha6c3:	data_out=16'h8a00;
17'ha6c4:	data_out=16'h806d;
17'ha6c5:	data_out=16'ha00;
17'ha6c6:	data_out=16'h225;
17'ha6c7:	data_out=16'h8a00;
17'ha6c8:	data_out=16'h8a00;
17'ha6c9:	data_out=16'h89ed;
17'ha6ca:	data_out=16'h8a00;
17'ha6cb:	data_out=16'h89f6;
17'ha6cc:	data_out=16'h896d;
17'ha6cd:	data_out=16'h8a00;
17'ha6ce:	data_out=16'h89d6;
17'ha6cf:	data_out=16'h8a00;
17'ha6d0:	data_out=16'h8549;
17'ha6d1:	data_out=16'h86;
17'ha6d2:	data_out=16'ha00;
17'ha6d3:	data_out=16'h8a00;
17'ha6d4:	data_out=16'h89c8;
17'ha6d5:	data_out=16'h881c;
17'ha6d6:	data_out=16'ha00;
17'ha6d7:	data_out=16'h20a;
17'ha6d8:	data_out=16'h9ea;
17'ha6d9:	data_out=16'ha00;
17'ha6da:	data_out=16'h8a00;
17'ha6db:	data_out=16'ha00;
17'ha6dc:	data_out=16'h8a00;
17'ha6dd:	data_out=16'h83ed;
17'ha6de:	data_out=16'h8a00;
17'ha6df:	data_out=16'h813f;
17'ha6e0:	data_out=16'h89ff;
17'ha6e1:	data_out=16'ha00;
17'ha6e2:	data_out=16'h8a00;
17'ha6e3:	data_out=16'h8a00;
17'ha6e4:	data_out=16'h880c;
17'ha6e5:	data_out=16'h8a00;
17'ha6e6:	data_out=16'h8a00;
17'ha6e7:	data_out=16'h8a00;
17'ha6e8:	data_out=16'ha00;
17'ha6e9:	data_out=16'h808;
17'ha6ea:	data_out=16'ha00;
17'ha6eb:	data_out=16'h795;
17'ha6ec:	data_out=16'ha00;
17'ha6ed:	data_out=16'h8a00;
17'ha6ee:	data_out=16'ha00;
17'ha6ef:	data_out=16'h8a00;
17'ha6f0:	data_out=16'ha00;
17'ha6f1:	data_out=16'h89fe;
17'ha6f2:	data_out=16'ha00;
17'ha6f3:	data_out=16'ha00;
17'ha6f4:	data_out=16'ha00;
17'ha6f5:	data_out=16'ha00;
17'ha6f6:	data_out=16'h8a00;
17'ha6f7:	data_out=16'h8a00;
17'ha6f8:	data_out=16'h8a00;
17'ha6f9:	data_out=16'h8865;
17'ha6fa:	data_out=16'h8a00;
17'ha6fb:	data_out=16'ha00;
17'ha6fc:	data_out=16'h4ae;
17'ha6fd:	data_out=16'h89fe;
17'ha6fe:	data_out=16'h8a00;
17'ha6ff:	data_out=16'ha00;
17'ha700:	data_out=16'h40f;
17'ha701:	data_out=16'h4ab;
17'ha702:	data_out=16'h3b2;
17'ha703:	data_out=16'h8a00;
17'ha704:	data_out=16'h12f;
17'ha705:	data_out=16'h6a;
17'ha706:	data_out=16'h88ad;
17'ha707:	data_out=16'h8a00;
17'ha708:	data_out=16'h80bf;
17'ha709:	data_out=16'h8a00;
17'ha70a:	data_out=16'h9d2;
17'ha70b:	data_out=16'h8a00;
17'ha70c:	data_out=16'h8a00;
17'ha70d:	data_out=16'h8a00;
17'ha70e:	data_out=16'h683;
17'ha70f:	data_out=16'h8402;
17'ha710:	data_out=16'h8a00;
17'ha711:	data_out=16'h8133;
17'ha712:	data_out=16'h8a00;
17'ha713:	data_out=16'h89fc;
17'ha714:	data_out=16'h8767;
17'ha715:	data_out=16'h2c4;
17'ha716:	data_out=16'h8474;
17'ha717:	data_out=16'h8a00;
17'ha718:	data_out=16'h6c;
17'ha719:	data_out=16'h89fd;
17'ha71a:	data_out=16'h4c;
17'ha71b:	data_out=16'h8a00;
17'ha71c:	data_out=16'h9ff;
17'ha71d:	data_out=16'h84f6;
17'ha71e:	data_out=16'h891c;
17'ha71f:	data_out=16'h8704;
17'ha720:	data_out=16'h89d6;
17'ha721:	data_out=16'h648;
17'ha722:	data_out=16'h8a00;
17'ha723:	data_out=16'h550;
17'ha724:	data_out=16'h552;
17'ha725:	data_out=16'h89f7;
17'ha726:	data_out=16'h89fc;
17'ha727:	data_out=16'h89cb;
17'ha728:	data_out=16'h529;
17'ha729:	data_out=16'h86e3;
17'ha72a:	data_out=16'h89fb;
17'ha72b:	data_out=16'h89ff;
17'ha72c:	data_out=16'h8309;
17'ha72d:	data_out=16'h844b;
17'ha72e:	data_out=16'h8a00;
17'ha72f:	data_out=16'h89fd;
17'ha730:	data_out=16'h743;
17'ha731:	data_out=16'h8227;
17'ha732:	data_out=16'h77d;
17'ha733:	data_out=16'h8811;
17'ha734:	data_out=16'h92;
17'ha735:	data_out=16'h85f8;
17'ha736:	data_out=16'h89f2;
17'ha737:	data_out=16'h259;
17'ha738:	data_out=16'ha00;
17'ha739:	data_out=16'h8717;
17'ha73a:	data_out=16'h8a00;
17'ha73b:	data_out=16'h81a9;
17'ha73c:	data_out=16'h18c;
17'ha73d:	data_out=16'h82b3;
17'ha73e:	data_out=16'h515;
17'ha73f:	data_out=16'he6;
17'ha740:	data_out=16'h89d1;
17'ha741:	data_out=16'h84e5;
17'ha742:	data_out=16'h8835;
17'ha743:	data_out=16'h8a00;
17'ha744:	data_out=16'h845a;
17'ha745:	data_out=16'h202;
17'ha746:	data_out=16'h571;
17'ha747:	data_out=16'h8a00;
17'ha748:	data_out=16'h8a00;
17'ha749:	data_out=16'h89f9;
17'ha74a:	data_out=16'h8a00;
17'ha74b:	data_out=16'h8a00;
17'ha74c:	data_out=16'h89eb;
17'ha74d:	data_out=16'h8a00;
17'ha74e:	data_out=16'h89fb;
17'ha74f:	data_out=16'h8a00;
17'ha750:	data_out=16'h8890;
17'ha751:	data_out=16'h41d;
17'ha752:	data_out=16'h67e;
17'ha753:	data_out=16'h89fc;
17'ha754:	data_out=16'h8905;
17'ha755:	data_out=16'h16f;
17'ha756:	data_out=16'h370;
17'ha757:	data_out=16'h18a;
17'ha758:	data_out=16'h9fe;
17'ha759:	data_out=16'h80c6;
17'ha75a:	data_out=16'h89fd;
17'ha75b:	data_out=16'ha00;
17'ha75c:	data_out=16'h897a;
17'ha75d:	data_out=16'h8344;
17'ha75e:	data_out=16'h89ff;
17'ha75f:	data_out=16'h80b1;
17'ha760:	data_out=16'h8536;
17'ha761:	data_out=16'ha00;
17'ha762:	data_out=16'h8a00;
17'ha763:	data_out=16'h88a5;
17'ha764:	data_out=16'h893e;
17'ha765:	data_out=16'h89fc;
17'ha766:	data_out=16'h89ff;
17'ha767:	data_out=16'h8a00;
17'ha768:	data_out=16'h5f6;
17'ha769:	data_out=16'h81e6;
17'ha76a:	data_out=16'h6ae;
17'ha76b:	data_out=16'h80f5;
17'ha76c:	data_out=16'h7cf;
17'ha76d:	data_out=16'h8878;
17'ha76e:	data_out=16'h6ad;
17'ha76f:	data_out=16'h88be;
17'ha770:	data_out=16'h697;
17'ha771:	data_out=16'h8538;
17'ha772:	data_out=16'ha00;
17'ha773:	data_out=16'h37b;
17'ha774:	data_out=16'h765;
17'ha775:	data_out=16'ha00;
17'ha776:	data_out=16'h89fe;
17'ha777:	data_out=16'h8a00;
17'ha778:	data_out=16'h8a00;
17'ha779:	data_out=16'h8986;
17'ha77a:	data_out=16'h88af;
17'ha77b:	data_out=16'h4f1;
17'ha77c:	data_out=16'h17f;
17'ha77d:	data_out=16'h89fc;
17'ha77e:	data_out=16'h89ff;
17'ha77f:	data_out=16'h6b;
17'ha780:	data_out=16'h8058;
17'ha781:	data_out=16'h9c;
17'ha782:	data_out=16'h8035;
17'ha783:	data_out=16'h8110;
17'ha784:	data_out=16'h8048;
17'ha785:	data_out=16'h80ac;
17'ha786:	data_out=16'h8011;
17'ha787:	data_out=16'h821f;
17'ha788:	data_out=16'h810b;
17'ha789:	data_out=16'h82e0;
17'ha78a:	data_out=16'h77;
17'ha78b:	data_out=16'h81eb;
17'ha78c:	data_out=16'h81e4;
17'ha78d:	data_out=16'h8131;
17'ha78e:	data_out=16'h39;
17'ha78f:	data_out=16'h802e;
17'ha790:	data_out=16'h81db;
17'ha791:	data_out=16'h80a3;
17'ha792:	data_out=16'h814a;
17'ha793:	data_out=16'h812b;
17'ha794:	data_out=16'h808d;
17'ha795:	data_out=16'h8005;
17'ha796:	data_out=16'h80bd;
17'ha797:	data_out=16'h8090;
17'ha798:	data_out=16'h8093;
17'ha799:	data_out=16'h80fb;
17'ha79a:	data_out=16'h808c;
17'ha79b:	data_out=16'h8193;
17'ha79c:	data_out=16'h801c;
17'ha79d:	data_out=16'h80b5;
17'ha79e:	data_out=16'h8115;
17'ha79f:	data_out=16'h8185;
17'ha7a0:	data_out=16'h8152;
17'ha7a1:	data_out=16'h34;
17'ha7a2:	data_out=16'h81ad;
17'ha7a3:	data_out=16'hde;
17'ha7a4:	data_out=16'hd7;
17'ha7a5:	data_out=16'h811c;
17'ha7a6:	data_out=16'h81e6;
17'ha7a7:	data_out=16'h8118;
17'ha7a8:	data_out=16'h28;
17'ha7a9:	data_out=16'h80a4;
17'ha7aa:	data_out=16'h8184;
17'ha7ab:	data_out=16'h81b2;
17'ha7ac:	data_out=16'h80bb;
17'ha7ad:	data_out=16'h78;
17'ha7ae:	data_out=16'h81b0;
17'ha7af:	data_out=16'h8121;
17'ha7b0:	data_out=16'h9;
17'ha7b1:	data_out=16'h8078;
17'ha7b2:	data_out=16'he;
17'ha7b3:	data_out=16'h80e9;
17'ha7b4:	data_out=16'h8031;
17'ha7b5:	data_out=16'h817a;
17'ha7b6:	data_out=16'h808c;
17'ha7b7:	data_out=16'h8034;
17'ha7b8:	data_out=16'h2a4;
17'ha7b9:	data_out=16'h8113;
17'ha7ba:	data_out=16'h81fe;
17'ha7bb:	data_out=16'h810d;
17'ha7bc:	data_out=16'h1b;
17'ha7bd:	data_out=16'h8150;
17'ha7be:	data_out=16'h1e;
17'ha7bf:	data_out=16'h80b4;
17'ha7c0:	data_out=16'h80da;
17'ha7c1:	data_out=16'h80d4;
17'ha7c2:	data_out=16'h809b;
17'ha7c3:	data_out=16'h811f;
17'ha7c4:	data_out=16'h80db;
17'ha7c5:	data_out=16'h8069;
17'ha7c6:	data_out=16'h9a;
17'ha7c7:	data_out=16'h8198;
17'ha7c8:	data_out=16'h81ff;
17'ha7c9:	data_out=16'h810f;
17'ha7ca:	data_out=16'h81fe;
17'ha7cb:	data_out=16'h8139;
17'ha7cc:	data_out=16'h8170;
17'ha7cd:	data_out=16'h8185;
17'ha7ce:	data_out=16'h819c;
17'ha7cf:	data_out=16'h8160;
17'ha7d0:	data_out=16'h811a;
17'ha7d1:	data_out=16'hd;
17'ha7d2:	data_out=16'h104;
17'ha7d3:	data_out=16'h8169;
17'ha7d4:	data_out=16'h808b;
17'ha7d5:	data_out=16'h80a6;
17'ha7d6:	data_out=16'h805b;
17'ha7d7:	data_out=16'h8051;
17'ha7d8:	data_out=16'h8022;
17'ha7d9:	data_out=16'h8075;
17'ha7da:	data_out=16'h80af;
17'ha7db:	data_out=16'h1f3;
17'ha7dc:	data_out=16'h80c1;
17'ha7dd:	data_out=16'h8046;
17'ha7de:	data_out=16'h813d;
17'ha7df:	data_out=16'h8098;
17'ha7e0:	data_out=16'h80c1;
17'ha7e1:	data_out=16'hc;
17'ha7e2:	data_out=16'h80d6;
17'ha7e3:	data_out=16'h80dc;
17'ha7e4:	data_out=16'h8131;
17'ha7e5:	data_out=16'h8221;
17'ha7e6:	data_out=16'h81b3;
17'ha7e7:	data_out=16'h812b;
17'ha7e8:	data_out=16'h28;
17'ha7e9:	data_out=16'h808f;
17'ha7ea:	data_out=16'h46;
17'ha7eb:	data_out=16'h8119;
17'ha7ec:	data_out=16'hcb;
17'ha7ed:	data_out=16'h80e2;
17'ha7ee:	data_out=16'h4f;
17'ha7ef:	data_out=16'h80d2;
17'ha7f0:	data_out=16'h37;
17'ha7f1:	data_out=16'h8171;
17'ha7f2:	data_out=16'h4b;
17'ha7f3:	data_out=16'h8028;
17'ha7f4:	data_out=16'h6;
17'ha7f5:	data_out=16'h13d;
17'ha7f6:	data_out=16'h8202;
17'ha7f7:	data_out=16'h816a;
17'ha7f8:	data_out=16'h8108;
17'ha7f9:	data_out=16'h815f;
17'ha7fa:	data_out=16'h80b2;
17'ha7fb:	data_out=16'h17;
17'ha7fc:	data_out=16'h8017;
17'ha7fd:	data_out=16'h8091;
17'ha7fe:	data_out=16'h8272;
17'ha7ff:	data_out=16'h8157;
17'ha800:	data_out=16'h46;
17'ha801:	data_out=16'h48;
17'ha802:	data_out=16'h20;
17'ha803:	data_out=16'h34;
17'ha804:	data_out=16'h4e;
17'ha805:	data_out=16'h4b;
17'ha806:	data_out=16'h29;
17'ha807:	data_out=16'h45;
17'ha808:	data_out=16'h22;
17'ha809:	data_out=16'h1a;
17'ha80a:	data_out=16'h46;
17'ha80b:	data_out=16'h1c;
17'ha80c:	data_out=16'h5c;
17'ha80d:	data_out=16'h35;
17'ha80e:	data_out=16'h18;
17'ha80f:	data_out=16'h2d;
17'ha810:	data_out=16'h8004;
17'ha811:	data_out=16'h62;
17'ha812:	data_out=16'h34;
17'ha813:	data_out=16'h37;
17'ha814:	data_out=16'h42;
17'ha815:	data_out=16'h41;
17'ha816:	data_out=16'h41;
17'ha817:	data_out=16'h4c;
17'ha818:	data_out=16'h1a;
17'ha819:	data_out=16'h36;
17'ha81a:	data_out=16'h62;
17'ha81b:	data_out=16'h2b;
17'ha81c:	data_out=16'h50;
17'ha81d:	data_out=16'h3f;
17'ha81e:	data_out=16'h30;
17'ha81f:	data_out=16'h27;
17'ha820:	data_out=16'h4a;
17'ha821:	data_out=16'h17;
17'ha822:	data_out=16'he;
17'ha823:	data_out=16'h24;
17'ha824:	data_out=16'h22;
17'ha825:	data_out=16'h30;
17'ha826:	data_out=16'h13;
17'ha827:	data_out=16'h35;
17'ha828:	data_out=16'h11;
17'ha829:	data_out=16'h2e;
17'ha82a:	data_out=16'h37;
17'ha82b:	data_out=16'h2b;
17'ha82c:	data_out=16'h48;
17'ha82d:	data_out=16'h2c;
17'ha82e:	data_out=16'h17;
17'ha82f:	data_out=16'h3a;
17'ha830:	data_out=16'h70;
17'ha831:	data_out=16'h56;
17'ha832:	data_out=16'h6e;
17'ha833:	data_out=16'h3f;
17'ha834:	data_out=16'h42;
17'ha835:	data_out=16'h68;
17'ha836:	data_out=16'h1c;
17'ha837:	data_out=16'h2f;
17'ha838:	data_out=16'h4a;
17'ha839:	data_out=16'h2a;
17'ha83a:	data_out=16'h29;
17'ha83b:	data_out=16'h49;
17'ha83c:	data_out=16'h1d;
17'ha83d:	data_out=16'h45;
17'ha83e:	data_out=16'hc;
17'ha83f:	data_out=16'h4e;
17'ha840:	data_out=16'h5d;
17'ha841:	data_out=16'h33;
17'ha842:	data_out=16'h42;
17'ha843:	data_out=16'h1e;
17'ha844:	data_out=16'h4f;
17'ha845:	data_out=16'h2a;
17'ha846:	data_out=16'hd;
17'ha847:	data_out=16'h40;
17'ha848:	data_out=16'h16;
17'ha849:	data_out=16'h3e;
17'ha84a:	data_out=16'h56;
17'ha84b:	data_out=16'h58;
17'ha84c:	data_out=16'h47;
17'ha84d:	data_out=16'h19;
17'ha84e:	data_out=16'h45;
17'ha84f:	data_out=16'h49;
17'ha850:	data_out=16'h45;
17'ha851:	data_out=16'h32;
17'ha852:	data_out=16'h2f;
17'ha853:	data_out=16'h42;
17'ha854:	data_out=16'h54;
17'ha855:	data_out=16'h16;
17'ha856:	data_out=16'h4f;
17'ha857:	data_out=16'h11;
17'ha858:	data_out=16'h18;
17'ha859:	data_out=16'h2d;
17'ha85a:	data_out=16'h8;
17'ha85b:	data_out=16'h53;
17'ha85c:	data_out=16'h48;
17'ha85d:	data_out=16'h3f;
17'ha85e:	data_out=16'h46;
17'ha85f:	data_out=16'h2c;
17'ha860:	data_out=16'h25;
17'ha861:	data_out=16'h62;
17'ha862:	data_out=16'h21;
17'ha863:	data_out=16'h3e;
17'ha864:	data_out=16'h52;
17'ha865:	data_out=16'h46;
17'ha866:	data_out=16'h3a;
17'ha867:	data_out=16'h19;
17'ha868:	data_out=16'hb;
17'ha869:	data_out=16'h26;
17'ha86a:	data_out=16'h17;
17'ha86b:	data_out=16'h5d;
17'ha86c:	data_out=16'h3d;
17'ha86d:	data_out=16'h46;
17'ha86e:	data_out=16'ha;
17'ha86f:	data_out=16'h54;
17'ha870:	data_out=16'h12;
17'ha871:	data_out=16'h28;
17'ha872:	data_out=16'h3e;
17'ha873:	data_out=16'h5b;
17'ha874:	data_out=16'h68;
17'ha875:	data_out=16'h42;
17'ha876:	data_out=16'h2f;
17'ha877:	data_out=16'h39;
17'ha878:	data_out=16'h2d;
17'ha879:	data_out=16'h15;
17'ha87a:	data_out=16'h46;
17'ha87b:	data_out=16'he;
17'ha87c:	data_out=16'hf;
17'ha87d:	data_out=16'h39;
17'ha87e:	data_out=16'hb;
17'ha87f:	data_out=16'h44;
17'ha880:	data_out=16'h56e;
17'ha881:	data_out=16'h68f;
17'ha882:	data_out=16'h1be;
17'ha883:	data_out=16'h17f;
17'ha884:	data_out=16'h8775;
17'ha885:	data_out=16'h85c6;
17'ha886:	data_out=16'h87ff;
17'ha887:	data_out=16'h8326;
17'ha888:	data_out=16'h234;
17'ha889:	data_out=16'h8145;
17'ha88a:	data_out=16'h801d;
17'ha88b:	data_out=16'h44;
17'ha88c:	data_out=16'h84c1;
17'ha88d:	data_out=16'h215;
17'ha88e:	data_out=16'h8161;
17'ha88f:	data_out=16'h17b;
17'ha890:	data_out=16'h3e7;
17'ha891:	data_out=16'h8762;
17'ha892:	data_out=16'h601;
17'ha893:	data_out=16'h8019;
17'ha894:	data_out=16'h30c;
17'ha895:	data_out=16'h823c;
17'ha896:	data_out=16'h8222;
17'ha897:	data_out=16'h50a;
17'ha898:	data_out=16'h80b2;
17'ha899:	data_out=16'h82c3;
17'ha89a:	data_out=16'h8873;
17'ha89b:	data_out=16'h6d4;
17'ha89c:	data_out=16'h8597;
17'ha89d:	data_out=16'h472;
17'ha89e:	data_out=16'h56d;
17'ha89f:	data_out=16'h893f;
17'ha8a0:	data_out=16'h987;
17'ha8a1:	data_out=16'h8156;
17'ha8a2:	data_out=16'h648;
17'ha8a3:	data_out=16'h82ec;
17'ha8a4:	data_out=16'h82ec;
17'ha8a5:	data_out=16'h34;
17'ha8a6:	data_out=16'h834b;
17'ha8a7:	data_out=16'h559;
17'ha8a8:	data_out=16'h8161;
17'ha8a9:	data_out=16'h41d;
17'ha8aa:	data_out=16'h71a;
17'ha8ab:	data_out=16'hbc;
17'ha8ac:	data_out=16'h8231;
17'ha8ad:	data_out=16'h991;
17'ha8ae:	data_out=16'h52a;
17'ha8af:	data_out=16'ha00;
17'ha8b0:	data_out=16'h883b;
17'ha8b1:	data_out=16'h8053;
17'ha8b2:	data_out=16'h880e;
17'ha8b3:	data_out=16'h344;
17'ha8b4:	data_out=16'h8019;
17'ha8b5:	data_out=16'h8894;
17'ha8b6:	data_out=16'h6c9;
17'ha8b7:	data_out=16'h1bc;
17'ha8b8:	data_out=16'h8425;
17'ha8b9:	data_out=16'h3a1;
17'ha8ba:	data_out=16'h721;
17'ha8bb:	data_out=16'h8729;
17'ha8bc:	data_out=16'h56e;
17'ha8bd:	data_out=16'h8252;
17'ha8be:	data_out=16'h815e;
17'ha8bf:	data_out=16'h877b;
17'ha8c0:	data_out=16'h866c;
17'ha8c1:	data_out=16'h1db;
17'ha8c2:	data_out=16'h846;
17'ha8c3:	data_out=16'h8956;
17'ha8c4:	data_out=16'h8698;
17'ha8c5:	data_out=16'h82e9;
17'ha8c6:	data_out=16'h426;
17'ha8c7:	data_out=16'h138;
17'ha8c8:	data_out=16'h5d2;
17'ha8c9:	data_out=16'h80b6;
17'ha8ca:	data_out=16'h80d3;
17'ha8cb:	data_out=16'h623;
17'ha8cc:	data_out=16'h3bb;
17'ha8cd:	data_out=16'h706;
17'ha8ce:	data_out=16'h52d;
17'ha8cf:	data_out=16'h18c;
17'ha8d0:	data_out=16'h8672;
17'ha8d1:	data_out=16'h86be;
17'ha8d2:	data_out=16'h8417;
17'ha8d3:	data_out=16'ha00;
17'ha8d4:	data_out=16'ha00;
17'ha8d5:	data_out=16'h80df;
17'ha8d6:	data_out=16'h8422;
17'ha8d7:	data_out=16'h8380;
17'ha8d8:	data_out=16'h8012;
17'ha8d9:	data_out=16'h8514;
17'ha8da:	data_out=16'h708;
17'ha8db:	data_out=16'h89fe;
17'ha8dc:	data_out=16'h203;
17'ha8dd:	data_out=16'h760;
17'ha8de:	data_out=16'ha00;
17'ha8df:	data_out=16'h45d;
17'ha8e0:	data_out=16'h8240;
17'ha8e1:	data_out=16'h88f2;
17'ha8e2:	data_out=16'h162;
17'ha8e3:	data_out=16'h367;
17'ha8e4:	data_out=16'h82aa;
17'ha8e5:	data_out=16'h82ab;
17'ha8e6:	data_out=16'h8379;
17'ha8e7:	data_out=16'h2eb;
17'ha8e8:	data_out=16'h8162;
17'ha8e9:	data_out=16'h257;
17'ha8ea:	data_out=16'h8164;
17'ha8eb:	data_out=16'h87e7;
17'ha8ec:	data_out=16'ha00;
17'ha8ed:	data_out=16'h37f;
17'ha8ee:	data_out=16'h8169;
17'ha8ef:	data_out=16'h8268;
17'ha8f0:	data_out=16'h8163;
17'ha8f1:	data_out=16'h4f;
17'ha8f2:	data_out=16'h87e3;
17'ha8f3:	data_out=16'h8724;
17'ha8f4:	data_out=16'h883f;
17'ha8f5:	data_out=16'h8818;
17'ha8f6:	data_out=16'h817b;
17'ha8f7:	data_out=16'h877c;
17'ha8f8:	data_out=16'h89bf;
17'ha8f9:	data_out=16'h4d5;
17'ha8fa:	data_out=16'h36d;
17'ha8fb:	data_out=16'h815c;
17'ha8fc:	data_out=16'h97;
17'ha8fd:	data_out=16'h89b2;
17'ha8fe:	data_out=16'h83e1;
17'ha8ff:	data_out=16'h872c;
17'ha900:	data_out=16'ha00;
17'ha901:	data_out=16'ha00;
17'ha902:	data_out=16'h54b;
17'ha903:	data_out=16'h7bb;
17'ha904:	data_out=16'h89fd;
17'ha905:	data_out=16'h89fb;
17'ha906:	data_out=16'h8a00;
17'ha907:	data_out=16'h846d;
17'ha908:	data_out=16'ha00;
17'ha909:	data_out=16'h811a;
17'ha90a:	data_out=16'h2cf;
17'ha90b:	data_out=16'h23d;
17'ha90c:	data_out=16'h88a7;
17'ha90d:	data_out=16'h9cf;
17'ha90e:	data_out=16'h82cc;
17'ha90f:	data_out=16'ha00;
17'ha910:	data_out=16'h9e5;
17'ha911:	data_out=16'h89fe;
17'ha912:	data_out=16'ha00;
17'ha913:	data_out=16'h536;
17'ha914:	data_out=16'h883;
17'ha915:	data_out=16'h8301;
17'ha916:	data_out=16'h8172;
17'ha917:	data_out=16'ha00;
17'ha918:	data_out=16'h86;
17'ha919:	data_out=16'h86ab;
17'ha91a:	data_out=16'h89fc;
17'ha91b:	data_out=16'h9ff;
17'ha91c:	data_out=16'h8a00;
17'ha91d:	data_out=16'ha00;
17'ha91e:	data_out=16'ha00;
17'ha91f:	data_out=16'h8a00;
17'ha920:	data_out=16'ha00;
17'ha921:	data_out=16'h82c6;
17'ha922:	data_out=16'ha00;
17'ha923:	data_out=16'h8692;
17'ha924:	data_out=16'h8694;
17'ha925:	data_out=16'hc2;
17'ha926:	data_out=16'h8754;
17'ha927:	data_out=16'ha00;
17'ha928:	data_out=16'h82ba;
17'ha929:	data_out=16'ha00;
17'ha92a:	data_out=16'ha00;
17'ha92b:	data_out=16'h42e;
17'ha92c:	data_out=16'h83a0;
17'ha92d:	data_out=16'ha00;
17'ha92e:	data_out=16'ha00;
17'ha92f:	data_out=16'ha00;
17'ha930:	data_out=16'h89fd;
17'ha931:	data_out=16'h619;
17'ha932:	data_out=16'h89fb;
17'ha933:	data_out=16'h997;
17'ha934:	data_out=16'h538;
17'ha935:	data_out=16'h89fa;
17'ha936:	data_out=16'ha00;
17'ha937:	data_out=16'h526;
17'ha938:	data_out=16'h829e;
17'ha939:	data_out=16'ha00;
17'ha93a:	data_out=16'h9ff;
17'ha93b:	data_out=16'h89fd;
17'ha93c:	data_out=16'h9cc;
17'ha93d:	data_out=16'h802c;
17'ha93e:	data_out=16'h82ac;
17'ha93f:	data_out=16'h89fb;
17'ha940:	data_out=16'h89fa;
17'ha941:	data_out=16'h5e6;
17'ha942:	data_out=16'ha00;
17'ha943:	data_out=16'h8a00;
17'ha944:	data_out=16'h89fc;
17'ha945:	data_out=16'h84be;
17'ha946:	data_out=16'ha00;
17'ha947:	data_out=16'h536;
17'ha948:	data_out=16'ha00;
17'ha949:	data_out=16'h81f9;
17'ha94a:	data_out=16'h32c;
17'ha94b:	data_out=16'ha00;
17'ha94c:	data_out=16'ha00;
17'ha94d:	data_out=16'ha00;
17'ha94e:	data_out=16'ha00;
17'ha94f:	data_out=16'h975;
17'ha950:	data_out=16'h89fd;
17'ha951:	data_out=16'h8a00;
17'ha952:	data_out=16'h8926;
17'ha953:	data_out=16'ha00;
17'ha954:	data_out=16'ha00;
17'ha955:	data_out=16'h832c;
17'ha956:	data_out=16'h8a00;
17'ha957:	data_out=16'h8a00;
17'ha958:	data_out=16'h80ec;
17'ha959:	data_out=16'h89fa;
17'ha95a:	data_out=16'ha00;
17'ha95b:	data_out=16'h89fc;
17'ha95c:	data_out=16'h9fa;
17'ha95d:	data_out=16'ha00;
17'ha95e:	data_out=16'ha00;
17'ha95f:	data_out=16'ha00;
17'ha960:	data_out=16'h837e;
17'ha961:	data_out=16'h89fb;
17'ha962:	data_out=16'h467;
17'ha963:	data_out=16'h9f4;
17'ha964:	data_out=16'h831f;
17'ha965:	data_out=16'h81c5;
17'ha966:	data_out=16'h8a00;
17'ha967:	data_out=16'h7c3;
17'ha968:	data_out=16'h82c2;
17'ha969:	data_out=16'ha00;
17'ha96a:	data_out=16'h82ec;
17'ha96b:	data_out=16'h89f9;
17'ha96c:	data_out=16'ha00;
17'ha96d:	data_out=16'ha00;
17'ha96e:	data_out=16'h82f5;
17'ha96f:	data_out=16'h8260;
17'ha970:	data_out=16'h82cc;
17'ha971:	data_out=16'h378;
17'ha972:	data_out=16'h89f9;
17'ha973:	data_out=16'h89fa;
17'ha974:	data_out=16'h89fb;
17'ha975:	data_out=16'h8a00;
17'ha976:	data_out=16'h82b1;
17'ha977:	data_out=16'h88a2;
17'ha978:	data_out=16'h8a00;
17'ha979:	data_out=16'ha00;
17'ha97a:	data_out=16'h9d6;
17'ha97b:	data_out=16'h82af;
17'ha97c:	data_out=16'h4ad;
17'ha97d:	data_out=16'h8a00;
17'ha97e:	data_out=16'h8a00;
17'ha97f:	data_out=16'h89ff;
17'ha980:	data_out=16'ha00;
17'ha981:	data_out=16'ha00;
17'ha982:	data_out=16'h9f8;
17'ha983:	data_out=16'h234;
17'ha984:	data_out=16'h8a00;
17'ha985:	data_out=16'h8a00;
17'ha986:	data_out=16'h89ff;
17'ha987:	data_out=16'h88c8;
17'ha988:	data_out=16'ha00;
17'ha989:	data_out=16'h885b;
17'ha98a:	data_out=16'h8690;
17'ha98b:	data_out=16'h752;
17'ha98c:	data_out=16'h8963;
17'ha98d:	data_out=16'h954;
17'ha98e:	data_out=16'h856e;
17'ha98f:	data_out=16'h9fe;
17'ha990:	data_out=16'h948;
17'ha991:	data_out=16'h89f7;
17'ha992:	data_out=16'ha00;
17'ha993:	data_out=16'h2a8;
17'ha994:	data_out=16'h985;
17'ha995:	data_out=16'h8a00;
17'ha996:	data_out=16'h8a00;
17'ha997:	data_out=16'h9f5;
17'ha998:	data_out=16'h121;
17'ha999:	data_out=16'h872d;
17'ha99a:	data_out=16'h8a00;
17'ha99b:	data_out=16'h9f4;
17'ha99c:	data_out=16'h89ea;
17'ha99d:	data_out=16'ha00;
17'ha99e:	data_out=16'h9f8;
17'ha99f:	data_out=16'h8a00;
17'ha9a0:	data_out=16'ha00;
17'ha9a1:	data_out=16'h856f;
17'ha9a2:	data_out=16'h9e5;
17'ha9a3:	data_out=16'h8a00;
17'ha9a4:	data_out=16'h8a00;
17'ha9a5:	data_out=16'h85cf;
17'ha9a6:	data_out=16'h8a00;
17'ha9a7:	data_out=16'h9fb;
17'ha9a8:	data_out=16'h858a;
17'ha9a9:	data_out=16'ha00;
17'ha9aa:	data_out=16'ha00;
17'ha9ab:	data_out=16'ha00;
17'ha9ac:	data_out=16'h8a00;
17'ha9ad:	data_out=16'ha00;
17'ha9ae:	data_out=16'h9f2;
17'ha9af:	data_out=16'ha00;
17'ha9b0:	data_out=16'h89f8;
17'ha9b1:	data_out=16'h84a6;
17'ha9b2:	data_out=16'h8a00;
17'ha9b3:	data_out=16'h9fa;
17'ha9b4:	data_out=16'ha00;
17'ha9b5:	data_out=16'h8a00;
17'ha9b6:	data_out=16'ha00;
17'ha9b7:	data_out=16'h9f4;
17'ha9b8:	data_out=16'h4cc;
17'ha9b9:	data_out=16'h9fc;
17'ha9ba:	data_out=16'h977;
17'ha9bb:	data_out=16'h8a00;
17'ha9bc:	data_out=16'h9fb;
17'ha9bd:	data_out=16'h87b1;
17'ha9be:	data_out=16'h858c;
17'ha9bf:	data_out=16'h8a00;
17'ha9c0:	data_out=16'h8a00;
17'ha9c1:	data_out=16'h9cb;
17'ha9c2:	data_out=16'h9d0;
17'ha9c3:	data_out=16'h8a00;
17'ha9c4:	data_out=16'h8a00;
17'ha9c5:	data_out=16'h8a00;
17'ha9c6:	data_out=16'ha00;
17'ha9c7:	data_out=16'h80ec;
17'ha9c8:	data_out=16'ha00;
17'ha9c9:	data_out=16'h8a00;
17'ha9ca:	data_out=16'h510;
17'ha9cb:	data_out=16'h9fe;
17'ha9cc:	data_out=16'h9f8;
17'ha9cd:	data_out=16'ha00;
17'ha9ce:	data_out=16'ha00;
17'ha9cf:	data_out=16'h40e;
17'ha9d0:	data_out=16'h8a00;
17'ha9d1:	data_out=16'h89ff;
17'ha9d2:	data_out=16'h8a00;
17'ha9d3:	data_out=16'ha00;
17'ha9d4:	data_out=16'ha00;
17'ha9d5:	data_out=16'h588;
17'ha9d6:	data_out=16'h8a00;
17'ha9d7:	data_out=16'h8a00;
17'ha9d8:	data_out=16'h98b;
17'ha9d9:	data_out=16'h8a00;
17'ha9da:	data_out=16'h9fa;
17'ha9db:	data_out=16'h8a00;
17'ha9dc:	data_out=16'h9f7;
17'ha9dd:	data_out=16'ha00;
17'ha9de:	data_out=16'ha00;
17'ha9df:	data_out=16'ha00;
17'ha9e0:	data_out=16'h8a00;
17'ha9e1:	data_out=16'h8a00;
17'ha9e2:	data_out=16'h9e8;
17'ha9e3:	data_out=16'h9fe;
17'ha9e4:	data_out=16'h9b;
17'ha9e5:	data_out=16'h89fc;
17'ha9e6:	data_out=16'h8a00;
17'ha9e7:	data_out=16'ha00;
17'ha9e8:	data_out=16'h8580;
17'ha9e9:	data_out=16'ha00;
17'ha9ea:	data_out=16'h857b;
17'ha9eb:	data_out=16'h8a00;
17'ha9ec:	data_out=16'ha00;
17'ha9ed:	data_out=16'h9fe;
17'ha9ee:	data_out=16'h857b;
17'ha9ef:	data_out=16'h8a00;
17'ha9f0:	data_out=16'h8575;
17'ha9f1:	data_out=16'h7fe;
17'ha9f2:	data_out=16'h8a00;
17'ha9f3:	data_out=16'h8a00;
17'ha9f4:	data_out=16'h89f3;
17'ha9f5:	data_out=16'h8a00;
17'ha9f6:	data_out=16'h88ab;
17'ha9f7:	data_out=16'h8913;
17'ha9f8:	data_out=16'h8a00;
17'ha9f9:	data_out=16'ha00;
17'ha9fa:	data_out=16'h9fa;
17'ha9fb:	data_out=16'h858c;
17'ha9fc:	data_out=16'h7a3;
17'ha9fd:	data_out=16'h8a00;
17'ha9fe:	data_out=16'h8a00;
17'ha9ff:	data_out=16'h89ff;
17'haa00:	data_out=16'h861a;
17'haa01:	data_out=16'h8942;
17'haa02:	data_out=16'h63b;
17'haa03:	data_out=16'h821c;
17'haa04:	data_out=16'h89f8;
17'haa05:	data_out=16'h89ff;
17'haa06:	data_out=16'h89ff;
17'haa07:	data_out=16'h89f3;
17'haa08:	data_out=16'h8051;
17'haa09:	data_out=16'h89ed;
17'haa0a:	data_out=16'h8a00;
17'haa0b:	data_out=16'h3c5;
17'haa0c:	data_out=16'h89ec;
17'haa0d:	data_out=16'h832;
17'haa0e:	data_out=16'h8153;
17'haa0f:	data_out=16'h362;
17'haa10:	data_out=16'h931;
17'haa11:	data_out=16'h89f1;
17'haa12:	data_out=16'ha00;
17'haa13:	data_out=16'h83dc;
17'haa14:	data_out=16'h770;
17'haa15:	data_out=16'h8a00;
17'haa16:	data_out=16'h89ff;
17'haa17:	data_out=16'h8d9;
17'haa18:	data_out=16'h811c;
17'haa19:	data_out=16'h8428;
17'haa1a:	data_out=16'h89ff;
17'haa1b:	data_out=16'h9a8;
17'haa1c:	data_out=16'h898a;
17'haa1d:	data_out=16'h89e6;
17'haa1e:	data_out=16'h816;
17'haa1f:	data_out=16'h89ff;
17'haa20:	data_out=16'h866b;
17'haa21:	data_out=16'h80f6;
17'haa22:	data_out=16'h9f3;
17'haa23:	data_out=16'h89c1;
17'haa24:	data_out=16'h89c1;
17'haa25:	data_out=16'h89ff;
17'haa26:	data_out=16'h8a00;
17'haa27:	data_out=16'h89e7;
17'haa28:	data_out=16'h80b5;
17'haa29:	data_out=16'h9d1;
17'haa2a:	data_out=16'h783;
17'haa2b:	data_out=16'ha00;
17'haa2c:	data_out=16'h89ff;
17'haa2d:	data_out=16'ha00;
17'haa2e:	data_out=16'h886;
17'haa2f:	data_out=16'h9fb;
17'haa30:	data_out=16'h8967;
17'haa31:	data_out=16'h89fa;
17'haa32:	data_out=16'h8a00;
17'haa33:	data_out=16'h919;
17'haa34:	data_out=16'h8893;
17'haa35:	data_out=16'h89fc;
17'haa36:	data_out=16'ha00;
17'haa37:	data_out=16'h5f8;
17'haa38:	data_out=16'h39b;
17'haa39:	data_out=16'h984;
17'haa3a:	data_out=16'h8398;
17'haa3b:	data_out=16'h8a00;
17'haa3c:	data_out=16'h9e9;
17'haa3d:	data_out=16'h89f0;
17'haa3e:	data_out=16'h80b7;
17'haa3f:	data_out=16'h89ff;
17'haa40:	data_out=16'h89ff;
17'haa41:	data_out=16'h8c1;
17'haa42:	data_out=16'h8054;
17'haa43:	data_out=16'h8a00;
17'haa44:	data_out=16'h89f9;
17'haa45:	data_out=16'h8a00;
17'haa46:	data_out=16'h9ff;
17'haa47:	data_out=16'h898b;
17'haa48:	data_out=16'ha00;
17'haa49:	data_out=16'h8a00;
17'haa4a:	data_out=16'h8738;
17'haa4b:	data_out=16'h8090;
17'haa4c:	data_out=16'h88f6;
17'haa4d:	data_out=16'ha00;
17'haa4e:	data_out=16'ha00;
17'haa4f:	data_out=16'h89c5;
17'haa50:	data_out=16'h89ff;
17'haa51:	data_out=16'h88a8;
17'haa52:	data_out=16'h8938;
17'haa53:	data_out=16'ha00;
17'haa54:	data_out=16'ha00;
17'haa55:	data_out=16'h6ca;
17'haa56:	data_out=16'h8a00;
17'haa57:	data_out=16'h8a00;
17'haa58:	data_out=16'h9e9;
17'haa59:	data_out=16'h89fc;
17'haa5a:	data_out=16'h9ec;
17'haa5b:	data_out=16'h89f8;
17'haa5c:	data_out=16'h89fe;
17'haa5d:	data_out=16'h9f1;
17'haa5e:	data_out=16'h9f1;
17'haa5f:	data_out=16'ha00;
17'haa60:	data_out=16'h89f7;
17'haa61:	data_out=16'h8a00;
17'haa62:	data_out=16'h757;
17'haa63:	data_out=16'h99a;
17'haa64:	data_out=16'h846e;
17'haa65:	data_out=16'h89f7;
17'haa66:	data_out=16'h89fb;
17'haa67:	data_out=16'h4bd;
17'haa68:	data_out=16'h80d3;
17'haa69:	data_out=16'h855c;
17'haa6a:	data_out=16'h81af;
17'haa6b:	data_out=16'h89fd;
17'haa6c:	data_out=16'h9ff;
17'haa6d:	data_out=16'h992;
17'haa6e:	data_out=16'h81ad;
17'haa6f:	data_out=16'h8a00;
17'haa70:	data_out=16'h8179;
17'haa71:	data_out=16'h898f;
17'haa72:	data_out=16'h8a00;
17'haa73:	data_out=16'h8a00;
17'haa74:	data_out=16'h895c;
17'haa75:	data_out=16'h8a00;
17'haa76:	data_out=16'h89f7;
17'haa77:	data_out=16'h8946;
17'haa78:	data_out=16'h8a00;
17'haa79:	data_out=16'h96b;
17'haa7a:	data_out=16'h8cf;
17'haa7b:	data_out=16'h80b7;
17'haa7c:	data_out=16'hd9;
17'haa7d:	data_out=16'h89fe;
17'haa7e:	data_out=16'h8a00;
17'haa7f:	data_out=16'h89fb;
17'haa80:	data_out=16'h89ef;
17'haa81:	data_out=16'h8a00;
17'haa82:	data_out=16'h89a2;
17'haa83:	data_out=16'h8a00;
17'haa84:	data_out=16'h89fa;
17'haa85:	data_out=16'h8a00;
17'haa86:	data_out=16'h89ff;
17'haa87:	data_out=16'h8431;
17'haa88:	data_out=16'h143;
17'haa89:	data_out=16'h866e;
17'haa8a:	data_out=16'h89da;
17'haa8b:	data_out=16'h1ff;
17'haa8c:	data_out=16'h9f1;
17'haa8d:	data_out=16'h82c9;
17'haa8e:	data_out=16'h6d1;
17'haa8f:	data_out=16'h89fd;
17'haa90:	data_out=16'h8a00;
17'haa91:	data_out=16'h8a00;
17'haa92:	data_out=16'h2b8;
17'haa93:	data_out=16'h86b8;
17'haa94:	data_out=16'h8a00;
17'haa95:	data_out=16'h8a00;
17'haa96:	data_out=16'h8a00;
17'haa97:	data_out=16'h8a00;
17'haa98:	data_out=16'h89ff;
17'haa99:	data_out=16'ha00;
17'haa9a:	data_out=16'h89fe;
17'haa9b:	data_out=16'h89ff;
17'haa9c:	data_out=16'h8a00;
17'haa9d:	data_out=16'h89ff;
17'haa9e:	data_out=16'h8a00;
17'haa9f:	data_out=16'h8a00;
17'haaa0:	data_out=16'h8a00;
17'haaa1:	data_out=16'h73f;
17'haaa2:	data_out=16'h972;
17'haaa3:	data_out=16'ha00;
17'haaa4:	data_out=16'ha00;
17'haaa5:	data_out=16'h85b7;
17'haaa6:	data_out=16'h9f8;
17'haaa7:	data_out=16'h8a00;
17'haaa8:	data_out=16'h72e;
17'haaa9:	data_out=16'h8c4;
17'haaaa:	data_out=16'h89fe;
17'haaab:	data_out=16'ha00;
17'haaac:	data_out=16'h8a00;
17'haaad:	data_out=16'h9ff;
17'haaae:	data_out=16'h893b;
17'haaaf:	data_out=16'h8a00;
17'haab0:	data_out=16'h85d2;
17'haab1:	data_out=16'h8a00;
17'haab2:	data_out=16'h89fb;
17'haab3:	data_out=16'h8a00;
17'haab4:	data_out=16'h89e2;
17'haab5:	data_out=16'h8a00;
17'haab6:	data_out=16'h89fc;
17'haab7:	data_out=16'h87e4;
17'haab8:	data_out=16'h8a00;
17'haab9:	data_out=16'h8a00;
17'haaba:	data_out=16'h89f5;
17'haabb:	data_out=16'h89fc;
17'haabc:	data_out=16'h8099;
17'haabd:	data_out=16'h8a00;
17'haabe:	data_out=16'h72a;
17'haabf:	data_out=16'h8a00;
17'haac0:	data_out=16'h89fb;
17'haac1:	data_out=16'h89ff;
17'haac2:	data_out=16'h9fe;
17'haac3:	data_out=16'h8a00;
17'haac4:	data_out=16'h8a00;
17'haac5:	data_out=16'h8a00;
17'haac6:	data_out=16'h9f9;
17'haac7:	data_out=16'h82c6;
17'haac8:	data_out=16'h89f5;
17'haac9:	data_out=16'h89ff;
17'haaca:	data_out=16'h89d5;
17'haacb:	data_out=16'h9fe;
17'haacc:	data_out=16'ha00;
17'haacd:	data_out=16'h9e1;
17'haace:	data_out=16'h8357;
17'haacf:	data_out=16'h3de;
17'haad0:	data_out=16'h8a00;
17'haad1:	data_out=16'h164;
17'haad2:	data_out=16'ha00;
17'haad3:	data_out=16'h8a00;
17'haad4:	data_out=16'h89fd;
17'haad5:	data_out=16'h30c;
17'haad6:	data_out=16'h8a00;
17'haad7:	data_out=16'h8a00;
17'haad8:	data_out=16'h806;
17'haad9:	data_out=16'h8a00;
17'haada:	data_out=16'h89ff;
17'haadb:	data_out=16'h8a00;
17'haadc:	data_out=16'h8a00;
17'haadd:	data_out=16'h89ff;
17'haade:	data_out=16'h8a00;
17'haadf:	data_out=16'h89fc;
17'haae0:	data_out=16'h9fe;
17'haae1:	data_out=16'h8a00;
17'haae2:	data_out=16'hd;
17'haae3:	data_out=16'h8a00;
17'haae4:	data_out=16'h8924;
17'haae5:	data_out=16'h8a00;
17'haae6:	data_out=16'h89fb;
17'haae7:	data_out=16'h82cb;
17'haae8:	data_out=16'h757;
17'haae9:	data_out=16'h993;
17'haaea:	data_out=16'h66e;
17'haaeb:	data_out=16'h8a00;
17'haaec:	data_out=16'h89dc;
17'haaed:	data_out=16'h8a00;
17'haaee:	data_out=16'h673;
17'haaef:	data_out=16'h89fe;
17'haaf0:	data_out=16'h6b4;
17'haaf1:	data_out=16'h89fa;
17'haaf2:	data_out=16'h8a00;
17'haaf3:	data_out=16'h8a00;
17'haaf4:	data_out=16'h854b;
17'haaf5:	data_out=16'h8a00;
17'haaf6:	data_out=16'h8971;
17'haaf7:	data_out=16'h8864;
17'haaf8:	data_out=16'h897b;
17'haaf9:	data_out=16'h8767;
17'haafa:	data_out=16'h8a00;
17'haafb:	data_out=16'h72c;
17'haafc:	data_out=16'h89ff;
17'haafd:	data_out=16'h8a00;
17'haafe:	data_out=16'h8a00;
17'haaff:	data_out=16'h8a00;
17'hab00:	data_out=16'h89ee;
17'hab01:	data_out=16'h8a00;
17'hab02:	data_out=16'h8ef;
17'hab03:	data_out=16'h8418;
17'hab04:	data_out=16'h89f2;
17'hab05:	data_out=16'h8a00;
17'hab06:	data_out=16'h89ff;
17'hab07:	data_out=16'ha00;
17'hab08:	data_out=16'h807b;
17'hab09:	data_out=16'h9c6;
17'hab0a:	data_out=16'h89cf;
17'hab0b:	data_out=16'h198;
17'hab0c:	data_out=16'ha00;
17'hab0d:	data_out=16'h9e0;
17'hab0e:	data_out=16'h9ec;
17'hab0f:	data_out=16'h350;
17'hab10:	data_out=16'h8a00;
17'hab11:	data_out=16'h8a00;
17'hab12:	data_out=16'h8106;
17'hab13:	data_out=16'h9ea;
17'hab14:	data_out=16'h89fe;
17'hab15:	data_out=16'h8a00;
17'hab16:	data_out=16'h89f5;
17'hab17:	data_out=16'h8788;
17'hab18:	data_out=16'h8822;
17'hab19:	data_out=16'ha00;
17'hab1a:	data_out=16'h8a00;
17'hab1b:	data_out=16'h82b1;
17'hab1c:	data_out=16'h8a00;
17'hab1d:	data_out=16'h8a00;
17'hab1e:	data_out=16'h89ff;
17'hab1f:	data_out=16'h8a00;
17'hab20:	data_out=16'h8a00;
17'hab21:	data_out=16'h9f4;
17'hab22:	data_out=16'h8fc;
17'hab23:	data_out=16'ha00;
17'hab24:	data_out=16'ha00;
17'hab25:	data_out=16'h9ca;
17'hab26:	data_out=16'ha00;
17'hab27:	data_out=16'h8a00;
17'hab28:	data_out=16'h9e5;
17'hab29:	data_out=16'h9f0;
17'hab2a:	data_out=16'h825c;
17'hab2b:	data_out=16'h881a;
17'hab2c:	data_out=16'h89fc;
17'hab2d:	data_out=16'ha00;
17'hab2e:	data_out=16'h89fe;
17'hab2f:	data_out=16'h8a00;
17'hab30:	data_out=16'h802b;
17'hab31:	data_out=16'h8a00;
17'hab32:	data_out=16'h89e9;
17'hab33:	data_out=16'h8a00;
17'hab34:	data_out=16'h8a00;
17'hab35:	data_out=16'h89fe;
17'hab36:	data_out=16'h89fa;
17'hab37:	data_out=16'h8f9;
17'hab38:	data_out=16'h8a00;
17'hab39:	data_out=16'h8a00;
17'hab3a:	data_out=16'h8616;
17'hab3b:	data_out=16'h89e9;
17'hab3c:	data_out=16'h4d3;
17'hab3d:	data_out=16'h8a00;
17'hab3e:	data_out=16'h9e4;
17'hab3f:	data_out=16'h8a00;
17'hab40:	data_out=16'h89f4;
17'hab41:	data_out=16'h8697;
17'hab42:	data_out=16'ha00;
17'hab43:	data_out=16'h8a00;
17'hab44:	data_out=16'h8a00;
17'hab45:	data_out=16'h8a00;
17'hab46:	data_out=16'ha00;
17'hab47:	data_out=16'h9f2;
17'hab48:	data_out=16'h89f9;
17'hab49:	data_out=16'h9d3;
17'hab4a:	data_out=16'h89e4;
17'hab4b:	data_out=16'ha00;
17'hab4c:	data_out=16'ha00;
17'hab4d:	data_out=16'h7fb;
17'hab4e:	data_out=16'h51d;
17'hab4f:	data_out=16'ha00;
17'hab50:	data_out=16'h8a00;
17'hab51:	data_out=16'h9a2;
17'hab52:	data_out=16'ha00;
17'hab53:	data_out=16'h89ff;
17'hab54:	data_out=16'h8a00;
17'hab55:	data_out=16'h9a9;
17'hab56:	data_out=16'h924;
17'hab57:	data_out=16'h8a00;
17'hab58:	data_out=16'h9b6;
17'hab59:	data_out=16'h89ff;
17'hab5a:	data_out=16'h89ec;
17'hab5b:	data_out=16'h8a00;
17'hab5c:	data_out=16'h8a00;
17'hab5d:	data_out=16'h8a00;
17'hab5e:	data_out=16'h8a00;
17'hab5f:	data_out=16'h89ff;
17'hab60:	data_out=16'ha00;
17'hab61:	data_out=16'h8a00;
17'hab62:	data_out=16'h65c;
17'hab63:	data_out=16'h8a00;
17'hab64:	data_out=16'h89fc;
17'hab65:	data_out=16'h8a00;
17'hab66:	data_out=16'h89cd;
17'hab67:	data_out=16'h39;
17'hab68:	data_out=16'h9f4;
17'hab69:	data_out=16'h9c2;
17'hab6a:	data_out=16'h9e0;
17'hab6b:	data_out=16'h8a00;
17'hab6c:	data_out=16'h89e0;
17'hab6d:	data_out=16'h8a00;
17'hab6e:	data_out=16'h9e1;
17'hab6f:	data_out=16'h89f0;
17'hab70:	data_out=16'h9e9;
17'hab71:	data_out=16'h88c7;
17'hab72:	data_out=16'h8a00;
17'hab73:	data_out=16'h8a00;
17'hab74:	data_out=16'h11b;
17'hab75:	data_out=16'h8a00;
17'hab76:	data_out=16'h858c;
17'hab77:	data_out=16'h9e1;
17'hab78:	data_out=16'h89fe;
17'hab79:	data_out=16'h37b;
17'hab7a:	data_out=16'h89ff;
17'hab7b:	data_out=16'h9e4;
17'hab7c:	data_out=16'h8a00;
17'hab7d:	data_out=16'h8a00;
17'hab7e:	data_out=16'h89f3;
17'hab7f:	data_out=16'h8a00;
17'hab80:	data_out=16'h89f8;
17'hab81:	data_out=16'h89ff;
17'hab82:	data_out=16'h9f8;
17'hab83:	data_out=16'h899;
17'hab84:	data_out=16'h8a00;
17'hab85:	data_out=16'h8a00;
17'hab86:	data_out=16'h8a00;
17'hab87:	data_out=16'ha00;
17'hab88:	data_out=16'h4b6;
17'hab89:	data_out=16'ha00;
17'hab8a:	data_out=16'h89f6;
17'hab8b:	data_out=16'h6f8;
17'hab8c:	data_out=16'ha00;
17'hab8d:	data_out=16'ha00;
17'hab8e:	data_out=16'h9fd;
17'hab8f:	data_out=16'ha00;
17'hab90:	data_out=16'h89ff;
17'hab91:	data_out=16'h8a00;
17'hab92:	data_out=16'h8006;
17'hab93:	data_out=16'ha00;
17'hab94:	data_out=16'h89dd;
17'hab95:	data_out=16'h8a00;
17'hab96:	data_out=16'h89b3;
17'hab97:	data_out=16'h543;
17'hab98:	data_out=16'h878d;
17'hab99:	data_out=16'h5b8;
17'hab9a:	data_out=16'h8a00;
17'hab9b:	data_out=16'h887;
17'hab9c:	data_out=16'h89f5;
17'hab9d:	data_out=16'h8a00;
17'hab9e:	data_out=16'h8981;
17'hab9f:	data_out=16'h8a00;
17'haba0:	data_out=16'h8a00;
17'haba1:	data_out=16'h9fc;
17'haba2:	data_out=16'h857;
17'haba3:	data_out=16'ha00;
17'haba4:	data_out=16'ha00;
17'haba5:	data_out=16'h9de;
17'haba6:	data_out=16'ha00;
17'haba7:	data_out=16'h89ff;
17'haba8:	data_out=16'h9f8;
17'haba9:	data_out=16'h9fc;
17'habaa:	data_out=16'ha00;
17'habab:	data_out=16'h8905;
17'habac:	data_out=16'h89f9;
17'habad:	data_out=16'ha00;
17'habae:	data_out=16'h51e;
17'habaf:	data_out=16'h89f9;
17'habb0:	data_out=16'h55c;
17'habb1:	data_out=16'h8a00;
17'habb2:	data_out=16'h8a00;
17'habb3:	data_out=16'h89f6;
17'habb4:	data_out=16'h89fe;
17'habb5:	data_out=16'h89f5;
17'habb6:	data_out=16'h88e3;
17'habb7:	data_out=16'h9f9;
17'habb8:	data_out=16'h8a00;
17'habb9:	data_out=16'h89fb;
17'habba:	data_out=16'h3a8;
17'habbb:	data_out=16'h89f3;
17'habbc:	data_out=16'h9fd;
17'habbd:	data_out=16'h8a00;
17'habbe:	data_out=16'h9f8;
17'habbf:	data_out=16'h8a00;
17'habc0:	data_out=16'h8a00;
17'habc1:	data_out=16'h803a;
17'habc2:	data_out=16'ha00;
17'habc3:	data_out=16'h8a00;
17'habc4:	data_out=16'h8a00;
17'habc5:	data_out=16'h8a00;
17'habc6:	data_out=16'ha00;
17'habc7:	data_out=16'ha00;
17'habc8:	data_out=16'h89f7;
17'habc9:	data_out=16'h9ec;
17'habca:	data_out=16'h89f3;
17'habcb:	data_out=16'ha00;
17'habcc:	data_out=16'h9ff;
17'habcd:	data_out=16'h2c9;
17'habce:	data_out=16'ha00;
17'habcf:	data_out=16'ha00;
17'habd0:	data_out=16'h8a00;
17'habd1:	data_out=16'h9f5;
17'habd2:	data_out=16'ha00;
17'habd3:	data_out=16'h89fb;
17'habd4:	data_out=16'h89fe;
17'habd5:	data_out=16'ha00;
17'habd6:	data_out=16'h9ed;
17'habd7:	data_out=16'h8242;
17'habd8:	data_out=16'h9f4;
17'habd9:	data_out=16'h8a00;
17'habda:	data_out=16'h83e0;
17'habdb:	data_out=16'h8a00;
17'habdc:	data_out=16'h89fe;
17'habdd:	data_out=16'h89f9;
17'habde:	data_out=16'h89fa;
17'habdf:	data_out=16'h89fa;
17'habe0:	data_out=16'ha00;
17'habe1:	data_out=16'h8a00;
17'habe2:	data_out=16'h9f2;
17'habe3:	data_out=16'h89f9;
17'habe4:	data_out=16'h89fc;
17'habe5:	data_out=16'h8a00;
17'habe6:	data_out=16'h899e;
17'habe7:	data_out=16'h902;
17'habe8:	data_out=16'h9fc;
17'habe9:	data_out=16'h9fc;
17'habea:	data_out=16'h9fc;
17'habeb:	data_out=16'h8a00;
17'habec:	data_out=16'h89ac;
17'habed:	data_out=16'h89f9;
17'habee:	data_out=16'h9fc;
17'habef:	data_out=16'h89ff;
17'habf0:	data_out=16'h9fc;
17'habf1:	data_out=16'h4bf;
17'habf2:	data_out=16'h8a00;
17'habf3:	data_out=16'h8a00;
17'habf4:	data_out=16'h6f7;
17'habf5:	data_out=16'h8a00;
17'habf6:	data_out=16'h9e5;
17'habf7:	data_out=16'ha00;
17'habf8:	data_out=16'h8a00;
17'habf9:	data_out=16'h9e7;
17'habfa:	data_out=16'h89ec;
17'habfb:	data_out=16'h9f8;
17'habfc:	data_out=16'h8a00;
17'habfd:	data_out=16'h8a00;
17'habfe:	data_out=16'h800b;
17'habff:	data_out=16'h8a00;
17'hac00:	data_out=16'h89f2;
17'hac01:	data_out=16'h8a00;
17'hac02:	data_out=16'ha00;
17'hac03:	data_out=16'ha00;
17'hac04:	data_out=16'h8a00;
17'hac05:	data_out=16'h8a00;
17'hac06:	data_out=16'h89fe;
17'hac07:	data_out=16'ha00;
17'hac08:	data_out=16'h109;
17'hac09:	data_out=16'ha00;
17'hac0a:	data_out=16'h8957;
17'hac0b:	data_out=16'h879b;
17'hac0c:	data_out=16'ha00;
17'hac0d:	data_out=16'ha00;
17'hac0e:	data_out=16'ha00;
17'hac0f:	data_out=16'ha00;
17'hac10:	data_out=16'h89f0;
17'hac11:	data_out=16'h8a00;
17'hac12:	data_out=16'h8290;
17'hac13:	data_out=16'ha00;
17'hac14:	data_out=16'h86b2;
17'hac15:	data_out=16'h89fd;
17'hac16:	data_out=16'h88f9;
17'hac17:	data_out=16'h3d;
17'hac18:	data_out=16'he8;
17'hac19:	data_out=16'h8578;
17'hac1a:	data_out=16'h8a00;
17'hac1b:	data_out=16'ha00;
17'hac1c:	data_out=16'h89da;
17'hac1d:	data_out=16'h8a00;
17'hac1e:	data_out=16'h85c1;
17'hac1f:	data_out=16'h89fa;
17'hac20:	data_out=16'h8a00;
17'hac21:	data_out=16'ha00;
17'hac22:	data_out=16'h9d1;
17'hac23:	data_out=16'ha00;
17'hac24:	data_out=16'ha00;
17'hac25:	data_out=16'ha00;
17'hac26:	data_out=16'ha00;
17'hac27:	data_out=16'h89ff;
17'hac28:	data_out=16'ha00;
17'hac29:	data_out=16'ha00;
17'hac2a:	data_out=16'ha00;
17'hac2b:	data_out=16'h89f5;
17'hac2c:	data_out=16'h89cb;
17'hac2d:	data_out=16'ha00;
17'hac2e:	data_out=16'h3ea;
17'hac2f:	data_out=16'h89f7;
17'hac30:	data_out=16'ha00;
17'hac31:	data_out=16'h8a00;
17'hac32:	data_out=16'h89fa;
17'hac33:	data_out=16'h89eb;
17'hac34:	data_out=16'h8a00;
17'hac35:	data_out=16'h89eb;
17'hac36:	data_out=16'h8769;
17'hac37:	data_out=16'ha00;
17'hac38:	data_out=16'h8a00;
17'hac39:	data_out=16'h89f2;
17'hac3a:	data_out=16'h776;
17'hac3b:	data_out=16'h89f4;
17'hac3c:	data_out=16'h7e1;
17'hac3d:	data_out=16'h89fe;
17'hac3e:	data_out=16'ha00;
17'hac3f:	data_out=16'h8a00;
17'hac40:	data_out=16'h89f0;
17'hac41:	data_out=16'h8160;
17'hac42:	data_out=16'ha00;
17'hac43:	data_out=16'h89ff;
17'hac44:	data_out=16'h8a00;
17'hac45:	data_out=16'h89fc;
17'hac46:	data_out=16'h9f2;
17'hac47:	data_out=16'ha00;
17'hac48:	data_out=16'h89c6;
17'hac49:	data_out=16'ha00;
17'hac4a:	data_out=16'h89f9;
17'hac4b:	data_out=16'h9e6;
17'hac4c:	data_out=16'ha00;
17'hac4d:	data_out=16'h825d;
17'hac4e:	data_out=16'ha00;
17'hac4f:	data_out=16'ha00;
17'hac50:	data_out=16'h89fc;
17'hac51:	data_out=16'ha00;
17'hac52:	data_out=16'ha00;
17'hac53:	data_out=16'h89fd;
17'hac54:	data_out=16'h89fe;
17'hac55:	data_out=16'ha00;
17'hac56:	data_out=16'ha00;
17'hac57:	data_out=16'h9c9;
17'hac58:	data_out=16'h9d9;
17'hac59:	data_out=16'h89e4;
17'hac5a:	data_out=16'h84f9;
17'hac5b:	data_out=16'h8a00;
17'hac5c:	data_out=16'h8a00;
17'hac5d:	data_out=16'h89bf;
17'hac5e:	data_out=16'h89f4;
17'hac5f:	data_out=16'h89eb;
17'hac60:	data_out=16'ha00;
17'hac61:	data_out=16'h8a00;
17'hac62:	data_out=16'h9ef;
17'hac63:	data_out=16'h89ee;
17'hac64:	data_out=16'h8a00;
17'hac65:	data_out=16'h8a00;
17'hac66:	data_out=16'h825d;
17'hac67:	data_out=16'ha00;
17'hac68:	data_out=16'ha00;
17'hac69:	data_out=16'h9fb;
17'hac6a:	data_out=16'ha00;
17'hac6b:	data_out=16'h8a00;
17'hac6c:	data_out=16'h89b0;
17'hac6d:	data_out=16'h89ee;
17'hac6e:	data_out=16'ha00;
17'hac6f:	data_out=16'h89fd;
17'hac70:	data_out=16'ha00;
17'hac71:	data_out=16'h99c;
17'hac72:	data_out=16'h8a00;
17'hac73:	data_out=16'h8a00;
17'hac74:	data_out=16'ha00;
17'hac75:	data_out=16'h8a00;
17'hac76:	data_out=16'h9f3;
17'hac77:	data_out=16'ha00;
17'hac78:	data_out=16'h8a00;
17'hac79:	data_out=16'h9d5;
17'hac7a:	data_out=16'h89da;
17'hac7b:	data_out=16'ha00;
17'hac7c:	data_out=16'h89fd;
17'hac7d:	data_out=16'h8a00;
17'hac7e:	data_out=16'h809c;
17'hac7f:	data_out=16'h8a00;
17'hac80:	data_out=16'h89e4;
17'hac81:	data_out=16'h8a00;
17'hac82:	data_out=16'ha00;
17'hac83:	data_out=16'ha00;
17'hac84:	data_out=16'h89de;
17'hac85:	data_out=16'h8a00;
17'hac86:	data_out=16'h89f7;
17'hac87:	data_out=16'ha00;
17'hac88:	data_out=16'h828c;
17'hac89:	data_out=16'ha00;
17'hac8a:	data_out=16'h5c;
17'hac8b:	data_out=16'h89d2;
17'hac8c:	data_out=16'ha00;
17'hac8d:	data_out=16'ha00;
17'hac8e:	data_out=16'ha00;
17'hac8f:	data_out=16'ha00;
17'hac90:	data_out=16'h89f3;
17'hac91:	data_out=16'h8a00;
17'hac92:	data_out=16'h84a8;
17'hac93:	data_out=16'h8196;
17'hac94:	data_out=16'h85d5;
17'hac95:	data_out=16'h89e3;
17'hac96:	data_out=16'h8701;
17'hac97:	data_out=16'h8281;
17'hac98:	data_out=16'h92a;
17'hac99:	data_out=16'h89fd;
17'hac9a:	data_out=16'h8a00;
17'hac9b:	data_out=16'ha00;
17'hac9c:	data_out=16'h899a;
17'hac9d:	data_out=16'h8a00;
17'hac9e:	data_out=16'h8521;
17'hac9f:	data_out=16'h89f5;
17'haca0:	data_out=16'h8a00;
17'haca1:	data_out=16'ha00;
17'haca2:	data_out=16'h8561;
17'haca3:	data_out=16'ha00;
17'haca4:	data_out=16'ha00;
17'haca5:	data_out=16'ha00;
17'haca6:	data_out=16'ha00;
17'haca7:	data_out=16'h8a00;
17'haca8:	data_out=16'ha00;
17'haca9:	data_out=16'h9ff;
17'hacaa:	data_out=16'ha00;
17'hacab:	data_out=16'h8a00;
17'hacac:	data_out=16'h88c8;
17'hacad:	data_out=16'h89e3;
17'hacae:	data_out=16'h4e;
17'hacaf:	data_out=16'h8a00;
17'hacb0:	data_out=16'ha00;
17'hacb1:	data_out=16'h8a00;
17'hacb2:	data_out=16'h875c;
17'hacb3:	data_out=16'h89f4;
17'hacb4:	data_out=16'h8a00;
17'hacb5:	data_out=16'h8909;
17'hacb6:	data_out=16'h889a;
17'hacb7:	data_out=16'ha00;
17'hacb8:	data_out=16'h8a00;
17'hacb9:	data_out=16'h89f7;
17'hacba:	data_out=16'h541;
17'hacbb:	data_out=16'h8990;
17'hacbc:	data_out=16'hb2;
17'hacbd:	data_out=16'h89ed;
17'hacbe:	data_out=16'ha00;
17'hacbf:	data_out=16'h8a00;
17'hacc0:	data_out=16'h8999;
17'hacc1:	data_out=16'ha00;
17'hacc2:	data_out=16'ha00;
17'hacc3:	data_out=16'h89ff;
17'hacc4:	data_out=16'h8a00;
17'hacc5:	data_out=16'h89e0;
17'hacc6:	data_out=16'h9ce;
17'hacc7:	data_out=16'h9d7;
17'hacc8:	data_out=16'h89c5;
17'hacc9:	data_out=16'ha00;
17'hacca:	data_out=16'h89ff;
17'haccb:	data_out=16'ha00;
17'haccc:	data_out=16'ha00;
17'haccd:	data_out=16'h89ef;
17'hacce:	data_out=16'h9f7;
17'haccf:	data_out=16'ha00;
17'hacd0:	data_out=16'h89f6;
17'hacd1:	data_out=16'ha00;
17'hacd2:	data_out=16'ha00;
17'hacd3:	data_out=16'h89ff;
17'hacd4:	data_out=16'h8a00;
17'hacd5:	data_out=16'ha00;
17'hacd6:	data_out=16'ha00;
17'hacd7:	data_out=16'h9fc;
17'hacd8:	data_out=16'h9f4;
17'hacd9:	data_out=16'h898c;
17'hacda:	data_out=16'h8697;
17'hacdb:	data_out=16'h8a00;
17'hacdc:	data_out=16'h89fd;
17'hacdd:	data_out=16'h8973;
17'hacde:	data_out=16'h89c2;
17'hacdf:	data_out=16'h89fa;
17'hace0:	data_out=16'ha00;
17'hace1:	data_out=16'h8985;
17'hace2:	data_out=16'h39a;
17'hace3:	data_out=16'h89fa;
17'hace4:	data_out=16'h8a00;
17'hace5:	data_out=16'h8a00;
17'hace6:	data_out=16'h89e9;
17'hace7:	data_out=16'ha00;
17'hace8:	data_out=16'ha00;
17'hace9:	data_out=16'h9e8;
17'hacea:	data_out=16'ha00;
17'haceb:	data_out=16'h8a00;
17'hacec:	data_out=16'h8998;
17'haced:	data_out=16'h89f9;
17'hacee:	data_out=16'ha00;
17'hacef:	data_out=16'h89be;
17'hacf0:	data_out=16'ha00;
17'hacf1:	data_out=16'h9fe;
17'hacf2:	data_out=16'h89da;
17'hacf3:	data_out=16'h89b4;
17'hacf4:	data_out=16'ha00;
17'hacf5:	data_out=16'h89fe;
17'hacf6:	data_out=16'h9d8;
17'hacf7:	data_out=16'ha00;
17'hacf8:	data_out=16'h8a00;
17'hacf9:	data_out=16'h9f8;
17'hacfa:	data_out=16'h89db;
17'hacfb:	data_out=16'ha00;
17'hacfc:	data_out=16'h8a00;
17'hacfd:	data_out=16'h8a00;
17'hacfe:	data_out=16'h89b5;
17'hacff:	data_out=16'h8a00;
17'had00:	data_out=16'h89dd;
17'had01:	data_out=16'h89fa;
17'had02:	data_out=16'ha00;
17'had03:	data_out=16'h9ff;
17'had04:	data_out=16'h89d8;
17'had05:	data_out=16'h89d2;
17'had06:	data_out=16'h892a;
17'had07:	data_out=16'ha00;
17'had08:	data_out=16'h9ed;
17'had09:	data_out=16'ha00;
17'had0a:	data_out=16'h1c3;
17'had0b:	data_out=16'h89fd;
17'had0c:	data_out=16'ha00;
17'had0d:	data_out=16'ha00;
17'had0e:	data_out=16'ha00;
17'had0f:	data_out=16'ha00;
17'had10:	data_out=16'h8a00;
17'had11:	data_out=16'h8a00;
17'had12:	data_out=16'h9c8;
17'had13:	data_out=16'h27f;
17'had14:	data_out=16'hf8;
17'had15:	data_out=16'h8610;
17'had16:	data_out=16'h9fe;
17'had17:	data_out=16'h3a4;
17'had18:	data_out=16'h9eb;
17'had19:	data_out=16'h8a00;
17'had1a:	data_out=16'h8a00;
17'had1b:	data_out=16'ha00;
17'had1c:	data_out=16'h884f;
17'had1d:	data_out=16'h8a00;
17'had1e:	data_out=16'h7bb;
17'had1f:	data_out=16'h926;
17'had20:	data_out=16'h8a00;
17'had21:	data_out=16'ha00;
17'had22:	data_out=16'h887e;
17'had23:	data_out=16'ha00;
17'had24:	data_out=16'ha00;
17'had25:	data_out=16'ha00;
17'had26:	data_out=16'ha00;
17'had27:	data_out=16'h8a00;
17'had28:	data_out=16'ha00;
17'had29:	data_out=16'ha00;
17'had2a:	data_out=16'h9ff;
17'had2b:	data_out=16'h8a00;
17'had2c:	data_out=16'h30;
17'had2d:	data_out=16'h8a00;
17'had2e:	data_out=16'h9eb;
17'had2f:	data_out=16'h89f3;
17'had30:	data_out=16'h9ff;
17'had31:	data_out=16'h8a00;
17'had32:	data_out=16'h289;
17'had33:	data_out=16'h89f6;
17'had34:	data_out=16'h8a00;
17'had35:	data_out=16'h350;
17'had36:	data_out=16'h9fc;
17'had37:	data_out=16'ha00;
17'had38:	data_out=16'h8a00;
17'had39:	data_out=16'h89fa;
17'had3a:	data_out=16'ha00;
17'had3b:	data_out=16'h9df;
17'had3c:	data_out=16'h9c7;
17'had3d:	data_out=16'h89e6;
17'had3e:	data_out=16'ha00;
17'had3f:	data_out=16'h89d0;
17'had40:	data_out=16'h89b0;
17'had41:	data_out=16'ha00;
17'had42:	data_out=16'ha00;
17'had43:	data_out=16'h8a00;
17'had44:	data_out=16'h8a00;
17'had45:	data_out=16'h84fc;
17'had46:	data_out=16'h9bc;
17'had47:	data_out=16'h99c;
17'had48:	data_out=16'h857c;
17'had49:	data_out=16'ha00;
17'had4a:	data_out=16'h89fe;
17'had4b:	data_out=16'h31f;
17'had4c:	data_out=16'ha00;
17'had4d:	data_out=16'h8a00;
17'had4e:	data_out=16'ha00;
17'had4f:	data_out=16'ha00;
17'had50:	data_out=16'h89e4;
17'had51:	data_out=16'ha00;
17'had52:	data_out=16'ha00;
17'had53:	data_out=16'h8a00;
17'had54:	data_out=16'h8a00;
17'had55:	data_out=16'ha00;
17'had56:	data_out=16'ha00;
17'had57:	data_out=16'h9fe;
17'had58:	data_out=16'ha00;
17'had59:	data_out=16'h89b3;
17'had5a:	data_out=16'h9be;
17'had5b:	data_out=16'h8a00;
17'had5c:	data_out=16'h883b;
17'had5d:	data_out=16'h84e8;
17'had5e:	data_out=16'h878d;
17'had5f:	data_out=16'h8a00;
17'had60:	data_out=16'ha00;
17'had61:	data_out=16'h88eb;
17'had62:	data_out=16'h9ff;
17'had63:	data_out=16'h89f5;
17'had64:	data_out=16'h8a00;
17'had65:	data_out=16'h8a00;
17'had66:	data_out=16'h89fc;
17'had67:	data_out=16'h9da;
17'had68:	data_out=16'ha00;
17'had69:	data_out=16'ha00;
17'had6a:	data_out=16'ha00;
17'had6b:	data_out=16'h89ff;
17'had6c:	data_out=16'h8963;
17'had6d:	data_out=16'h89f6;
17'had6e:	data_out=16'ha00;
17'had6f:	data_out=16'h8926;
17'had70:	data_out=16'ha00;
17'had71:	data_out=16'ha00;
17'had72:	data_out=16'h89d2;
17'had73:	data_out=16'h89cc;
17'had74:	data_out=16'h9ff;
17'had75:	data_out=16'h9cf;
17'had76:	data_out=16'h886;
17'had77:	data_out=16'ha00;
17'had78:	data_out=16'h8a00;
17'had79:	data_out=16'ha00;
17'had7a:	data_out=16'h8619;
17'had7b:	data_out=16'ha00;
17'had7c:	data_out=16'h24d;
17'had7d:	data_out=16'h89fc;
17'had7e:	data_out=16'h89d9;
17'had7f:	data_out=16'h8a00;
17'had80:	data_out=16'h89e8;
17'had81:	data_out=16'h89f4;
17'had82:	data_out=16'ha00;
17'had83:	data_out=16'h8583;
17'had84:	data_out=16'h89e3;
17'had85:	data_out=16'h8999;
17'had86:	data_out=16'h887a;
17'had87:	data_out=16'ha00;
17'had88:	data_out=16'h9f3;
17'had89:	data_out=16'ha00;
17'had8a:	data_out=16'h8366;
17'had8b:	data_out=16'h8a00;
17'had8c:	data_out=16'ha00;
17'had8d:	data_out=16'ha00;
17'had8e:	data_out=16'ha00;
17'had8f:	data_out=16'ha00;
17'had90:	data_out=16'h8a00;
17'had91:	data_out=16'h8a00;
17'had92:	data_out=16'h9f0;
17'had93:	data_out=16'h330;
17'had94:	data_out=16'h89a1;
17'had95:	data_out=16'h8432;
17'had96:	data_out=16'h9fc;
17'had97:	data_out=16'h888d;
17'had98:	data_out=16'ha00;
17'had99:	data_out=16'h8a00;
17'had9a:	data_out=16'h8a00;
17'had9b:	data_out=16'ha00;
17'had9c:	data_out=16'h89b2;
17'had9d:	data_out=16'h8a00;
17'had9e:	data_out=16'h8397;
17'had9f:	data_out=16'h8f4;
17'hada0:	data_out=16'h8a00;
17'hada1:	data_out=16'ha00;
17'hada2:	data_out=16'h89f2;
17'hada3:	data_out=16'ha00;
17'hada4:	data_out=16'ha00;
17'hada5:	data_out=16'ha00;
17'hada6:	data_out=16'ha00;
17'hada7:	data_out=16'h8a00;
17'hada8:	data_out=16'ha00;
17'hada9:	data_out=16'h329;
17'hadaa:	data_out=16'h9ff;
17'hadab:	data_out=16'h8a00;
17'hadac:	data_out=16'h270;
17'hadad:	data_out=16'h8a00;
17'hadae:	data_out=16'h9e7;
17'hadaf:	data_out=16'h89fd;
17'hadb0:	data_out=16'h9fc;
17'hadb1:	data_out=16'h8a00;
17'hadb2:	data_out=16'h86c6;
17'hadb3:	data_out=16'h8a00;
17'hadb4:	data_out=16'h89ef;
17'hadb5:	data_out=16'h15b;
17'hadb6:	data_out=16'h9fb;
17'hadb7:	data_out=16'ha00;
17'hadb8:	data_out=16'h8a00;
17'hadb9:	data_out=16'h8a00;
17'hadba:	data_out=16'h207;
17'hadbb:	data_out=16'h9fc;
17'hadbc:	data_out=16'h88e2;
17'hadbd:	data_out=16'h8a00;
17'hadbe:	data_out=16'ha00;
17'hadbf:	data_out=16'h8972;
17'hadc0:	data_out=16'h89d0;
17'hadc1:	data_out=16'ha00;
17'hadc2:	data_out=16'ha00;
17'hadc3:	data_out=16'h8a00;
17'hadc4:	data_out=16'h8a00;
17'hadc5:	data_out=16'h8364;
17'hadc6:	data_out=16'h89e8;
17'hadc7:	data_out=16'h96f;
17'hadc8:	data_out=16'h8392;
17'hadc9:	data_out=16'ha00;
17'hadca:	data_out=16'h220;
17'hadcb:	data_out=16'h886b;
17'hadcc:	data_out=16'ha00;
17'hadcd:	data_out=16'h8a00;
17'hadce:	data_out=16'ha00;
17'hadcf:	data_out=16'ha00;
17'hadd0:	data_out=16'h8a00;
17'hadd1:	data_out=16'ha00;
17'hadd2:	data_out=16'ha00;
17'hadd3:	data_out=16'h8a00;
17'hadd4:	data_out=16'h8a00;
17'hadd5:	data_out=16'ha00;
17'hadd6:	data_out=16'ha00;
17'hadd7:	data_out=16'h9ff;
17'hadd8:	data_out=16'ha00;
17'hadd9:	data_out=16'h89db;
17'hadda:	data_out=16'h9b4;
17'haddb:	data_out=16'h8a00;
17'haddc:	data_out=16'hfd;
17'haddd:	data_out=16'h80e6;
17'hadde:	data_out=16'h8562;
17'haddf:	data_out=16'h8a00;
17'hade0:	data_out=16'ha00;
17'hade1:	data_out=16'h89d5;
17'hade2:	data_out=16'h8853;
17'hade3:	data_out=16'h8a00;
17'hade4:	data_out=16'h8a00;
17'hade5:	data_out=16'h8a00;
17'hade6:	data_out=16'h8a00;
17'hade7:	data_out=16'h8a00;
17'hade8:	data_out=16'ha00;
17'hade9:	data_out=16'ha00;
17'hadea:	data_out=16'ha00;
17'hadeb:	data_out=16'h89ff;
17'hadec:	data_out=16'h83;
17'haded:	data_out=16'h8a00;
17'hadee:	data_out=16'ha00;
17'hadef:	data_out=16'h87a1;
17'hadf0:	data_out=16'ha00;
17'hadf1:	data_out=16'ha00;
17'hadf2:	data_out=16'h89de;
17'hadf3:	data_out=16'h89ee;
17'hadf4:	data_out=16'h9fe;
17'hadf5:	data_out=16'ha00;
17'hadf6:	data_out=16'h8a00;
17'hadf7:	data_out=16'ha00;
17'hadf8:	data_out=16'h8a00;
17'hadf9:	data_out=16'ha00;
17'hadfa:	data_out=16'h89fb;
17'hadfb:	data_out=16'ha00;
17'hadfc:	data_out=16'h9e8;
17'hadfd:	data_out=16'h89fc;
17'hadfe:	data_out=16'h89fd;
17'hadff:	data_out=16'h8a00;
17'hae00:	data_out=16'h8a00;
17'hae01:	data_out=16'h8a00;
17'hae02:	data_out=16'ha00;
17'hae03:	data_out=16'h89ad;
17'hae04:	data_out=16'h89de;
17'hae05:	data_out=16'h9df;
17'hae06:	data_out=16'h8959;
17'hae07:	data_out=16'ha00;
17'hae08:	data_out=16'h97e;
17'hae09:	data_out=16'h89cd;
17'hae0a:	data_out=16'h80d9;
17'hae0b:	data_out=16'h8a00;
17'hae0c:	data_out=16'h9f0;
17'hae0d:	data_out=16'ha00;
17'hae0e:	data_out=16'ha00;
17'hae0f:	data_out=16'ha00;
17'hae10:	data_out=16'h8a00;
17'hae11:	data_out=16'h8a00;
17'hae12:	data_out=16'h89f9;
17'hae13:	data_out=16'h841e;
17'hae14:	data_out=16'h8a00;
17'hae15:	data_out=16'h89d6;
17'hae16:	data_out=16'h8543;
17'hae17:	data_out=16'h89fe;
17'hae18:	data_out=16'h9e5;
17'hae19:	data_out=16'h8a00;
17'hae1a:	data_out=16'h89fc;
17'hae1b:	data_out=16'h2dd;
17'hae1c:	data_out=16'h89af;
17'hae1d:	data_out=16'h8a00;
17'hae1e:	data_out=16'h89fd;
17'hae1f:	data_out=16'h89fe;
17'hae20:	data_out=16'h8a00;
17'hae21:	data_out=16'ha00;
17'hae22:	data_out=16'h89fd;
17'hae23:	data_out=16'ha00;
17'hae24:	data_out=16'ha00;
17'hae25:	data_out=16'h85a6;
17'hae26:	data_out=16'ha00;
17'hae27:	data_out=16'h8a00;
17'hae28:	data_out=16'ha00;
17'hae29:	data_out=16'h89e2;
17'hae2a:	data_out=16'h1d7;
17'hae2b:	data_out=16'h8a00;
17'hae2c:	data_out=16'h8961;
17'hae2d:	data_out=16'h8a00;
17'hae2e:	data_out=16'h89f0;
17'hae2f:	data_out=16'h8a00;
17'hae30:	data_out=16'h9fd;
17'hae31:	data_out=16'h83cb;
17'hae32:	data_out=16'h984;
17'hae33:	data_out=16'h8a00;
17'hae34:	data_out=16'h89fe;
17'hae35:	data_out=16'h89f9;
17'hae36:	data_out=16'h8849;
17'hae37:	data_out=16'ha00;
17'hae38:	data_out=16'h89eb;
17'hae39:	data_out=16'h8a00;
17'hae3a:	data_out=16'h8a00;
17'hae3b:	data_out=16'ha00;
17'hae3c:	data_out=16'h89b4;
17'hae3d:	data_out=16'h8a00;
17'hae3e:	data_out=16'ha00;
17'hae3f:	data_out=16'h9e7;
17'hae40:	data_out=16'h89e4;
17'hae41:	data_out=16'ha00;
17'hae42:	data_out=16'h865a;
17'hae43:	data_out=16'h8a00;
17'hae44:	data_out=16'h8a00;
17'hae45:	data_out=16'h89d3;
17'hae46:	data_out=16'h89ac;
17'hae47:	data_out=16'h8a00;
17'hae48:	data_out=16'h89ee;
17'hae49:	data_out=16'h894e;
17'hae4a:	data_out=16'h82c4;
17'hae4b:	data_out=16'h89e3;
17'hae4c:	data_out=16'ha00;
17'hae4d:	data_out=16'h8a00;
17'hae4e:	data_out=16'h81c8;
17'hae4f:	data_out=16'h89a3;
17'hae50:	data_out=16'h8a00;
17'hae51:	data_out=16'ha00;
17'hae52:	data_out=16'ha00;
17'hae53:	data_out=16'h8a00;
17'hae54:	data_out=16'h8a00;
17'hae55:	data_out=16'ha00;
17'hae56:	data_out=16'ha00;
17'hae57:	data_out=16'h8924;
17'hae58:	data_out=16'ha00;
17'hae59:	data_out=16'h8a00;
17'hae5a:	data_out=16'h9ca;
17'hae5b:	data_out=16'h8a00;
17'hae5c:	data_out=16'h9ff;
17'hae5d:	data_out=16'h8859;
17'hae5e:	data_out=16'h8806;
17'hae5f:	data_out=16'h8a00;
17'hae60:	data_out=16'h9e4;
17'hae61:	data_out=16'h85c2;
17'hae62:	data_out=16'h89f1;
17'hae63:	data_out=16'h8a00;
17'hae64:	data_out=16'h8a00;
17'hae65:	data_out=16'h8a00;
17'hae66:	data_out=16'h8a00;
17'hae67:	data_out=16'h8a00;
17'hae68:	data_out=16'ha00;
17'hae69:	data_out=16'h9a7;
17'hae6a:	data_out=16'ha00;
17'hae6b:	data_out=16'h8a00;
17'hae6c:	data_out=16'h12a;
17'hae6d:	data_out=16'h8a00;
17'hae6e:	data_out=16'ha00;
17'hae6f:	data_out=16'h81b7;
17'hae70:	data_out=16'ha00;
17'hae71:	data_out=16'h9f1;
17'hae72:	data_out=16'h89c8;
17'hae73:	data_out=16'h89d8;
17'hae74:	data_out=16'ha00;
17'hae75:	data_out=16'ha00;
17'hae76:	data_out=16'h8a00;
17'hae77:	data_out=16'h89cb;
17'hae78:	data_out=16'h8a00;
17'hae79:	data_out=16'ha00;
17'hae7a:	data_out=16'h8a00;
17'hae7b:	data_out=16'ha00;
17'hae7c:	data_out=16'h72;
17'hae7d:	data_out=16'h8a00;
17'hae7e:	data_out=16'h89fc;
17'hae7f:	data_out=16'h8a00;
17'hae80:	data_out=16'h89e8;
17'hae81:	data_out=16'h813f;
17'hae82:	data_out=16'h9be;
17'hae83:	data_out=16'h89d1;
17'hae84:	data_out=16'h89f5;
17'hae85:	data_out=16'ha00;
17'hae86:	data_out=16'h89e7;
17'hae87:	data_out=16'h975;
17'hae88:	data_out=16'h89b2;
17'hae89:	data_out=16'h8a00;
17'hae8a:	data_out=16'h3d0;
17'hae8b:	data_out=16'h8a00;
17'hae8c:	data_out=16'h158;
17'hae8d:	data_out=16'h9ff;
17'hae8e:	data_out=16'ha00;
17'hae8f:	data_out=16'h89fb;
17'hae90:	data_out=16'h8a00;
17'hae91:	data_out=16'h8a00;
17'hae92:	data_out=16'h8a00;
17'hae93:	data_out=16'h8581;
17'hae94:	data_out=16'h8a00;
17'hae95:	data_out=16'h89e7;
17'hae96:	data_out=16'h8114;
17'hae97:	data_out=16'h89c9;
17'hae98:	data_out=16'h8a00;
17'hae99:	data_out=16'h8a00;
17'hae9a:	data_out=16'h9f3;
17'hae9b:	data_out=16'h8446;
17'hae9c:	data_out=16'h93e;
17'hae9d:	data_out=16'h8a00;
17'hae9e:	data_out=16'h8a00;
17'hae9f:	data_out=16'h8a00;
17'haea0:	data_out=16'h8a00;
17'haea1:	data_out=16'ha00;
17'haea2:	data_out=16'h8a00;
17'haea3:	data_out=16'h993;
17'haea4:	data_out=16'h995;
17'haea5:	data_out=16'h8a00;
17'haea6:	data_out=16'h89d0;
17'haea7:	data_out=16'h8a00;
17'haea8:	data_out=16'ha00;
17'haea9:	data_out=16'h8a00;
17'haeaa:	data_out=16'h89fc;
17'haeab:	data_out=16'h8a00;
17'haeac:	data_out=16'h84af;
17'haead:	data_out=16'h8a00;
17'haeae:	data_out=16'h89ff;
17'haeaf:	data_out=16'h89f7;
17'haeb0:	data_out=16'ha00;
17'haeb1:	data_out=16'h9dc;
17'haeb2:	data_out=16'h968;
17'haeb3:	data_out=16'h8a00;
17'haeb4:	data_out=16'h89be;
17'haeb5:	data_out=16'h8a00;
17'haeb6:	data_out=16'h89fb;
17'haeb7:	data_out=16'h396;
17'haeb8:	data_out=16'ha00;
17'haeb9:	data_out=16'h8a00;
17'haeba:	data_out=16'h8a00;
17'haebb:	data_out=16'h98c;
17'haebc:	data_out=16'h949;
17'haebd:	data_out=16'h8a00;
17'haebe:	data_out=16'ha00;
17'haebf:	data_out=16'ha00;
17'haec0:	data_out=16'h89a1;
17'haec1:	data_out=16'ha00;
17'haec2:	data_out=16'h89c3;
17'haec3:	data_out=16'h8a00;
17'haec4:	data_out=16'h89fa;
17'haec5:	data_out=16'h89e3;
17'haec6:	data_out=16'h33b;
17'haec7:	data_out=16'h8a00;
17'haec8:	data_out=16'h89f7;
17'haec9:	data_out=16'h8a00;
17'haeca:	data_out=16'h89ff;
17'haecb:	data_out=16'h8a00;
17'haecc:	data_out=16'h89b8;
17'haecd:	data_out=16'h8a00;
17'haece:	data_out=16'h89f1;
17'haecf:	data_out=16'h8a00;
17'haed0:	data_out=16'h8a00;
17'haed1:	data_out=16'h9fd;
17'haed2:	data_out=16'h170;
17'haed3:	data_out=16'h89f9;
17'haed4:	data_out=16'h8a00;
17'haed5:	data_out=16'h89b8;
17'haed6:	data_out=16'h87a9;
17'haed7:	data_out=16'h8a00;
17'haed8:	data_out=16'ha00;
17'haed9:	data_out=16'h8a00;
17'haeda:	data_out=16'h9ff;
17'haedb:	data_out=16'h8a00;
17'haedc:	data_out=16'ha00;
17'haedd:	data_out=16'h89e9;
17'haede:	data_out=16'h891d;
17'haedf:	data_out=16'h8a00;
17'haee0:	data_out=16'h8a00;
17'haee1:	data_out=16'h9d7;
17'haee2:	data_out=16'h89e6;
17'haee3:	data_out=16'h8a00;
17'haee4:	data_out=16'h8a00;
17'haee5:	data_out=16'h8a00;
17'haee6:	data_out=16'h8a00;
17'haee7:	data_out=16'h8a00;
17'haee8:	data_out=16'ha00;
17'haee9:	data_out=16'h89f7;
17'haeea:	data_out=16'ha00;
17'haeeb:	data_out=16'h89f6;
17'haeec:	data_out=16'h85d9;
17'haeed:	data_out=16'h8a00;
17'haeee:	data_out=16'ha00;
17'haeef:	data_out=16'ha00;
17'haef0:	data_out=16'ha00;
17'haef1:	data_out=16'h89f8;
17'haef2:	data_out=16'h899b;
17'haef3:	data_out=16'h9de;
17'haef4:	data_out=16'ha00;
17'haef5:	data_out=16'ha00;
17'haef6:	data_out=16'h8a00;
17'haef7:	data_out=16'h89ff;
17'haef8:	data_out=16'h8a00;
17'haef9:	data_out=16'h8255;
17'haefa:	data_out=16'h89fd;
17'haefb:	data_out=16'ha00;
17'haefc:	data_out=16'h89ff;
17'haefd:	data_out=16'h8a00;
17'haefe:	data_out=16'h8a00;
17'haeff:	data_out=16'h860c;
17'haf00:	data_out=16'h89ed;
17'haf01:	data_out=16'h8525;
17'haf02:	data_out=16'h89f9;
17'haf03:	data_out=16'h843a;
17'haf04:	data_out=16'h8a00;
17'haf05:	data_out=16'ha00;
17'haf06:	data_out=16'h8906;
17'haf07:	data_out=16'h8a00;
17'haf08:	data_out=16'h89e6;
17'haf09:	data_out=16'h8a00;
17'haf0a:	data_out=16'h8a00;
17'haf0b:	data_out=16'h8a00;
17'haf0c:	data_out=16'h8a00;
17'haf0d:	data_out=16'h9ff;
17'haf0e:	data_out=16'h9ff;
17'haf0f:	data_out=16'h8a00;
17'haf10:	data_out=16'h8a00;
17'haf11:	data_out=16'h8a00;
17'haf12:	data_out=16'h89f8;
17'haf13:	data_out=16'h1c8;
17'haf14:	data_out=16'h765;
17'haf15:	data_out=16'h89fb;
17'haf16:	data_out=16'h82f;
17'haf17:	data_out=16'h9f5;
17'haf18:	data_out=16'h8a00;
17'haf19:	data_out=16'h8a00;
17'haf1a:	data_out=16'ha00;
17'haf1b:	data_out=16'h65d;
17'haf1c:	data_out=16'ha00;
17'haf1d:	data_out=16'h8a00;
17'haf1e:	data_out=16'h89fb;
17'haf1f:	data_out=16'h89f4;
17'haf20:	data_out=16'h89ef;
17'haf21:	data_out=16'ha00;
17'haf22:	data_out=16'h8a00;
17'haf23:	data_out=16'h8a00;
17'haf24:	data_out=16'h8a00;
17'haf25:	data_out=16'h8a00;
17'haf26:	data_out=16'h8a00;
17'haf27:	data_out=16'h8a00;
17'haf28:	data_out=16'ha00;
17'haf29:	data_out=16'h8a00;
17'haf2a:	data_out=16'h8a00;
17'haf2b:	data_out=16'h89ff;
17'haf2c:	data_out=16'h7a0;
17'haf2d:	data_out=16'h8a00;
17'haf2e:	data_out=16'h89f9;
17'haf2f:	data_out=16'h8901;
17'haf30:	data_out=16'h86b;
17'haf31:	data_out=16'h31b;
17'haf32:	data_out=16'h8a00;
17'haf33:	data_out=16'h8997;
17'haf34:	data_out=16'h8953;
17'haf35:	data_out=16'h8a00;
17'haf36:	data_out=16'h89fd;
17'haf37:	data_out=16'h8a00;
17'haf38:	data_out=16'ha00;
17'haf39:	data_out=16'h89ca;
17'haf3a:	data_out=16'h8a00;
17'haf3b:	data_out=16'h8a00;
17'haf3c:	data_out=16'h9e2;
17'haf3d:	data_out=16'h8a00;
17'haf3e:	data_out=16'ha00;
17'haf3f:	data_out=16'ha00;
17'haf40:	data_out=16'h8a00;
17'haf41:	data_out=16'h9fe;
17'haf42:	data_out=16'h8a00;
17'haf43:	data_out=16'h8a00;
17'haf44:	data_out=16'h89f4;
17'haf45:	data_out=16'h89fa;
17'haf46:	data_out=16'h859e;
17'haf47:	data_out=16'h8a00;
17'haf48:	data_out=16'h89f1;
17'haf49:	data_out=16'h8a00;
17'haf4a:	data_out=16'h8a00;
17'haf4b:	data_out=16'h8a00;
17'haf4c:	data_out=16'h8a00;
17'haf4d:	data_out=16'h8a00;
17'haf4e:	data_out=16'h8a00;
17'haf4f:	data_out=16'h8a00;
17'haf50:	data_out=16'h8442;
17'haf51:	data_out=16'ha00;
17'haf52:	data_out=16'h8a00;
17'haf53:	data_out=16'h89b3;
17'haf54:	data_out=16'h89f7;
17'haf55:	data_out=16'h85bf;
17'haf56:	data_out=16'h8a00;
17'haf57:	data_out=16'h8a00;
17'haf58:	data_out=16'ha00;
17'haf59:	data_out=16'h8a00;
17'haf5a:	data_out=16'ha00;
17'haf5b:	data_out=16'h8a00;
17'haf5c:	data_out=16'ha00;
17'haf5d:	data_out=16'h89f9;
17'haf5e:	data_out=16'h8872;
17'haf5f:	data_out=16'h8a00;
17'haf60:	data_out=16'h8a00;
17'haf61:	data_out=16'h91c;
17'haf62:	data_out=16'h8992;
17'haf63:	data_out=16'h84b7;
17'haf64:	data_out=16'h8a00;
17'haf65:	data_out=16'h8a00;
17'haf66:	data_out=16'h89f3;
17'haf67:	data_out=16'h8a00;
17'haf68:	data_out=16'ha00;
17'haf69:	data_out=16'h8a00;
17'haf6a:	data_out=16'h9ff;
17'haf6b:	data_out=16'h89b2;
17'haf6c:	data_out=16'h893d;
17'haf6d:	data_out=16'h879f;
17'haf6e:	data_out=16'h9ff;
17'haf6f:	data_out=16'ha00;
17'haf70:	data_out=16'h9ff;
17'haf71:	data_out=16'h89fd;
17'haf72:	data_out=16'h89fd;
17'haf73:	data_out=16'h9d2;
17'haf74:	data_out=16'h9f4;
17'haf75:	data_out=16'ha00;
17'haf76:	data_out=16'h8a00;
17'haf77:	data_out=16'h8a00;
17'haf78:	data_out=16'h80e;
17'haf79:	data_out=16'h8939;
17'haf7a:	data_out=16'h210;
17'haf7b:	data_out=16'ha00;
17'haf7c:	data_out=16'h89ff;
17'haf7d:	data_out=16'h89ef;
17'haf7e:	data_out=16'h89e6;
17'haf7f:	data_out=16'ha00;
17'haf80:	data_out=16'h89fd;
17'haf81:	data_out=16'h8a00;
17'haf82:	data_out=16'h8a00;
17'haf83:	data_out=16'h41b;
17'haf84:	data_out=16'h8a00;
17'haf85:	data_out=16'h9c2;
17'haf86:	data_out=16'hd0;
17'haf87:	data_out=16'h8a00;
17'haf88:	data_out=16'h8a00;
17'haf89:	data_out=16'h8a00;
17'haf8a:	data_out=16'h8a00;
17'haf8b:	data_out=16'h8a00;
17'haf8c:	data_out=16'h8a00;
17'haf8d:	data_out=16'h9f2;
17'haf8e:	data_out=16'h9f9;
17'haf8f:	data_out=16'h8a00;
17'haf90:	data_out=16'h8a00;
17'haf91:	data_out=16'h8a00;
17'haf92:	data_out=16'h9f5;
17'haf93:	data_out=16'h9fa;
17'haf94:	data_out=16'h9f3;
17'haf95:	data_out=16'h8a00;
17'haf96:	data_out=16'h89ff;
17'haf97:	data_out=16'ha00;
17'haf98:	data_out=16'h89fb;
17'haf99:	data_out=16'h8a00;
17'haf9a:	data_out=16'h89f8;
17'haf9b:	data_out=16'h79f;
17'haf9c:	data_out=16'h9d6;
17'haf9d:	data_out=16'h8a00;
17'haf9e:	data_out=16'h87e6;
17'haf9f:	data_out=16'had;
17'hafa0:	data_out=16'h89f0;
17'hafa1:	data_out=16'h9fe;
17'hafa2:	data_out=16'h89ec;
17'hafa3:	data_out=16'h8a00;
17'hafa4:	data_out=16'h8a00;
17'hafa5:	data_out=16'h8a00;
17'hafa6:	data_out=16'h8a00;
17'hafa7:	data_out=16'h8a00;
17'hafa8:	data_out=16'h9ff;
17'hafa9:	data_out=16'h8a00;
17'hafaa:	data_out=16'h8a00;
17'hafab:	data_out=16'h89d1;
17'hafac:	data_out=16'h89ff;
17'hafad:	data_out=16'h8a00;
17'hafae:	data_out=16'h8978;
17'hafaf:	data_out=16'h884b;
17'hafb0:	data_out=16'h8a00;
17'hafb1:	data_out=16'h8a00;
17'hafb2:	data_out=16'h8a00;
17'hafb3:	data_out=16'ha00;
17'hafb4:	data_out=16'h89ff;
17'hafb5:	data_out=16'h8a00;
17'hafb6:	data_out=16'h8a00;
17'hafb7:	data_out=16'h8a00;
17'hafb8:	data_out=16'ha00;
17'hafb9:	data_out=16'ha00;
17'hafba:	data_out=16'h8a00;
17'hafbb:	data_out=16'h8a00;
17'hafbc:	data_out=16'h949;
17'hafbd:	data_out=16'h8a00;
17'hafbe:	data_out=16'h9ff;
17'hafbf:	data_out=16'h9bf;
17'hafc0:	data_out=16'h8a00;
17'hafc1:	data_out=16'h94b;
17'hafc2:	data_out=16'h8a00;
17'hafc3:	data_out=16'h385;
17'hafc4:	data_out=16'h8a00;
17'hafc5:	data_out=16'h8a00;
17'hafc6:	data_out=16'h8a00;
17'hafc7:	data_out=16'h8a00;
17'hafc8:	data_out=16'h8944;
17'hafc9:	data_out=16'h8a00;
17'hafca:	data_out=16'h8a00;
17'hafcb:	data_out=16'h8a00;
17'hafcc:	data_out=16'h8a00;
17'hafcd:	data_out=16'h8a00;
17'hafce:	data_out=16'h279;
17'hafcf:	data_out=16'h8a00;
17'hafd0:	data_out=16'ha;
17'hafd1:	data_out=16'ha00;
17'hafd2:	data_out=16'h8a00;
17'hafd3:	data_out=16'h87b3;
17'hafd4:	data_out=16'h89f1;
17'hafd5:	data_out=16'h85e4;
17'hafd6:	data_out=16'h8a00;
17'hafd7:	data_out=16'h8a00;
17'hafd8:	data_out=16'ha00;
17'hafd9:	data_out=16'h8a00;
17'hafda:	data_out=16'ha00;
17'hafdb:	data_out=16'h8a00;
17'hafdc:	data_out=16'ha00;
17'hafdd:	data_out=16'h89f8;
17'hafde:	data_out=16'h8806;
17'hafdf:	data_out=16'h89ff;
17'hafe0:	data_out=16'h8a00;
17'hafe1:	data_out=16'h8a00;
17'hafe2:	data_out=16'h64b;
17'hafe3:	data_out=16'ha00;
17'hafe4:	data_out=16'h8a00;
17'hafe5:	data_out=16'h8a00;
17'hafe6:	data_out=16'h89fa;
17'hafe7:	data_out=16'h8a00;
17'hafe8:	data_out=16'h9ff;
17'hafe9:	data_out=16'h8a00;
17'hafea:	data_out=16'h9d1;
17'hafeb:	data_out=16'h8a00;
17'hafec:	data_out=16'h89f1;
17'hafed:	data_out=16'ha00;
17'hafee:	data_out=16'h9d4;
17'hafef:	data_out=16'h38c;
17'haff0:	data_out=16'h9f7;
17'haff1:	data_out=16'h89f5;
17'haff2:	data_out=16'h8a00;
17'haff3:	data_out=16'h8a00;
17'haff4:	data_out=16'h8a00;
17'haff5:	data_out=16'ha00;
17'haff6:	data_out=16'h8a00;
17'haff7:	data_out=16'h8a00;
17'haff8:	data_out=16'ha00;
17'haff9:	data_out=16'h89a3;
17'haffa:	data_out=16'h9ff;
17'haffb:	data_out=16'h9ff;
17'haffc:	data_out=16'h89f6;
17'haffd:	data_out=16'h8946;
17'haffe:	data_out=16'h89b1;
17'hafff:	data_out=16'ha00;
17'hb000:	data_out=16'h8a00;
17'hb001:	data_out=16'h8a00;
17'hb002:	data_out=16'h8a00;
17'hb003:	data_out=16'h6b6;
17'hb004:	data_out=16'h8a00;
17'hb005:	data_out=16'h8a00;
17'hb006:	data_out=16'h9f7;
17'hb007:	data_out=16'h8a00;
17'hb008:	data_out=16'h8a00;
17'hb009:	data_out=16'h8a00;
17'hb00a:	data_out=16'h8a00;
17'hb00b:	data_out=16'h323;
17'hb00c:	data_out=16'h8a00;
17'hb00d:	data_out=16'h965;
17'hb00e:	data_out=16'h9a1;
17'hb00f:	data_out=16'h89fe;
17'hb010:	data_out=16'h89fb;
17'hb011:	data_out=16'h8a00;
17'hb012:	data_out=16'h9f6;
17'hb013:	data_out=16'h845a;
17'hb014:	data_out=16'h9e6;
17'hb015:	data_out=16'h8a00;
17'hb016:	data_out=16'h8a00;
17'hb017:	data_out=16'h9fc;
17'hb018:	data_out=16'h89fa;
17'hb019:	data_out=16'h89ec;
17'hb01a:	data_out=16'h8a00;
17'hb01b:	data_out=16'h94f;
17'hb01c:	data_out=16'h996;
17'hb01d:	data_out=16'h8a00;
17'hb01e:	data_out=16'h22b;
17'hb01f:	data_out=16'h956;
17'hb020:	data_out=16'h89ff;
17'hb021:	data_out=16'h9fe;
17'hb022:	data_out=16'h8977;
17'hb023:	data_out=16'h8a00;
17'hb024:	data_out=16'h8a00;
17'hb025:	data_out=16'h8a00;
17'hb026:	data_out=16'h8a00;
17'hb027:	data_out=16'h8a00;
17'hb028:	data_out=16'h9ff;
17'hb029:	data_out=16'h9a6;
17'hb02a:	data_out=16'h8a00;
17'hb02b:	data_out=16'h9d2;
17'hb02c:	data_out=16'h8a00;
17'hb02d:	data_out=16'h89fd;
17'hb02e:	data_out=16'h9dc;
17'hb02f:	data_out=16'h8457;
17'hb030:	data_out=16'h8a00;
17'hb031:	data_out=16'h8a00;
17'hb032:	data_out=16'h8a00;
17'hb033:	data_out=16'ha00;
17'hb034:	data_out=16'h8a00;
17'hb035:	data_out=16'h8a00;
17'hb036:	data_out=16'h8a00;
17'hb037:	data_out=16'h83c0;
17'hb038:	data_out=16'h53e;
17'hb039:	data_out=16'ha00;
17'hb03a:	data_out=16'h8a00;
17'hb03b:	data_out=16'h8a00;
17'hb03c:	data_out=16'h771;
17'hb03d:	data_out=16'h8a00;
17'hb03e:	data_out=16'h9ff;
17'hb03f:	data_out=16'h8a00;
17'hb040:	data_out=16'h8a00;
17'hb041:	data_out=16'h8a00;
17'hb042:	data_out=16'h8a00;
17'hb043:	data_out=16'h9ea;
17'hb044:	data_out=16'h8a00;
17'hb045:	data_out=16'h8a00;
17'hb046:	data_out=16'h8a00;
17'hb047:	data_out=16'h8a00;
17'hb048:	data_out=16'h9f9;
17'hb049:	data_out=16'h8a00;
17'hb04a:	data_out=16'h89f7;
17'hb04b:	data_out=16'h8a00;
17'hb04c:	data_out=16'h8a00;
17'hb04d:	data_out=16'h8981;
17'hb04e:	data_out=16'h99e;
17'hb04f:	data_out=16'h8a00;
17'hb050:	data_out=16'h229;
17'hb051:	data_out=16'h974;
17'hb052:	data_out=16'h8a00;
17'hb053:	data_out=16'h2b6;
17'hb054:	data_out=16'h89f3;
17'hb055:	data_out=16'h854e;
17'hb056:	data_out=16'h8a00;
17'hb057:	data_out=16'h8a00;
17'hb058:	data_out=16'h9fb;
17'hb059:	data_out=16'h8a00;
17'hb05a:	data_out=16'ha00;
17'hb05b:	data_out=16'h8a00;
17'hb05c:	data_out=16'ha00;
17'hb05d:	data_out=16'h89fb;
17'hb05e:	data_out=16'h8673;
17'hb05f:	data_out=16'h89fb;
17'hb060:	data_out=16'h8a00;
17'hb061:	data_out=16'h8a00;
17'hb062:	data_out=16'h9d0;
17'hb063:	data_out=16'ha00;
17'hb064:	data_out=16'h8a00;
17'hb065:	data_out=16'h8a00;
17'hb066:	data_out=16'h89c6;
17'hb067:	data_out=16'h89c2;
17'hb068:	data_out=16'h9ff;
17'hb069:	data_out=16'h8a00;
17'hb06a:	data_out=16'h8cf;
17'hb06b:	data_out=16'h8a00;
17'hb06c:	data_out=16'h8a00;
17'hb06d:	data_out=16'ha00;
17'hb06e:	data_out=16'h8d2;
17'hb06f:	data_out=16'h89f1;
17'hb070:	data_out=16'h94a;
17'hb071:	data_out=16'h85a4;
17'hb072:	data_out=16'h8a00;
17'hb073:	data_out=16'h8a00;
17'hb074:	data_out=16'h8a00;
17'hb075:	data_out=16'h9bd;
17'hb076:	data_out=16'h85d7;
17'hb077:	data_out=16'h8a00;
17'hb078:	data_out=16'ha00;
17'hb079:	data_out=16'h89c6;
17'hb07a:	data_out=16'h9fe;
17'hb07b:	data_out=16'h9ff;
17'hb07c:	data_out=16'h89f7;
17'hb07d:	data_out=16'h1f1;
17'hb07e:	data_out=16'h1f3;
17'hb07f:	data_out=16'h875e;
17'hb080:	data_out=16'h8a00;
17'hb081:	data_out=16'h8a00;
17'hb082:	data_out=16'h989;
17'hb083:	data_out=16'h86f8;
17'hb084:	data_out=16'h8a00;
17'hb085:	data_out=16'h8a00;
17'hb086:	data_out=16'h9ed;
17'hb087:	data_out=16'h8a00;
17'hb088:	data_out=16'h86e0;
17'hb089:	data_out=16'h89f0;
17'hb08a:	data_out=16'h8a00;
17'hb08b:	data_out=16'ha00;
17'hb08c:	data_out=16'h89de;
17'hb08d:	data_out=16'h8a00;
17'hb08e:	data_out=16'h9fb;
17'hb08f:	data_out=16'h86e5;
17'hb090:	data_out=16'h8540;
17'hb091:	data_out=16'h8a00;
17'hb092:	data_out=16'h989;
17'hb093:	data_out=16'h8758;
17'hb094:	data_out=16'h9ec;
17'hb095:	data_out=16'h8a00;
17'hb096:	data_out=16'h8a00;
17'hb097:	data_out=16'h9f3;
17'hb098:	data_out=16'h8a00;
17'hb099:	data_out=16'h9f8;
17'hb09a:	data_out=16'h8a00;
17'hb09b:	data_out=16'h9e8;
17'hb09c:	data_out=16'h84c3;
17'hb09d:	data_out=16'h8a00;
17'hb09e:	data_out=16'h86d8;
17'hb09f:	data_out=16'h7b2;
17'hb0a0:	data_out=16'h8a00;
17'hb0a1:	data_out=16'h9fe;
17'hb0a2:	data_out=16'h9f1;
17'hb0a3:	data_out=16'h8a00;
17'hb0a4:	data_out=16'h8a00;
17'hb0a5:	data_out=16'h8a00;
17'hb0a6:	data_out=16'h89fd;
17'hb0a7:	data_out=16'h8a00;
17'hb0a8:	data_out=16'ha00;
17'hb0a9:	data_out=16'h9ee;
17'hb0aa:	data_out=16'h8a00;
17'hb0ab:	data_out=16'ha00;
17'hb0ac:	data_out=16'h8a00;
17'hb0ad:	data_out=16'h9f7;
17'hb0ae:	data_out=16'h9ce;
17'hb0af:	data_out=16'h8678;
17'hb0b0:	data_out=16'h8a00;
17'hb0b1:	data_out=16'h8a00;
17'hb0b2:	data_out=16'h8a00;
17'hb0b3:	data_out=16'h9fa;
17'hb0b4:	data_out=16'h8a00;
17'hb0b5:	data_out=16'h8a00;
17'hb0b6:	data_out=16'h89ad;
17'hb0b7:	data_out=16'h9a2;
17'hb0b8:	data_out=16'h88bb;
17'hb0b9:	data_out=16'h9f9;
17'hb0ba:	data_out=16'h8a00;
17'hb0bb:	data_out=16'h8a00;
17'hb0bc:	data_out=16'h9d8;
17'hb0bd:	data_out=16'h8a00;
17'hb0be:	data_out=16'ha00;
17'hb0bf:	data_out=16'h8a00;
17'hb0c0:	data_out=16'h8a00;
17'hb0c1:	data_out=16'h8a00;
17'hb0c2:	data_out=16'h89ff;
17'hb0c3:	data_out=16'h9f4;
17'hb0c4:	data_out=16'h8a00;
17'hb0c5:	data_out=16'h8a00;
17'hb0c6:	data_out=16'h9f9;
17'hb0c7:	data_out=16'h8a00;
17'hb0c8:	data_out=16'h9ea;
17'hb0c9:	data_out=16'h8a00;
17'hb0ca:	data_out=16'h8742;
17'hb0cb:	data_out=16'h89fa;
17'hb0cc:	data_out=16'h89fe;
17'hb0cd:	data_out=16'h9f1;
17'hb0ce:	data_out=16'h9d7;
17'hb0cf:	data_out=16'h8a00;
17'hb0d0:	data_out=16'h899f;
17'hb0d1:	data_out=16'h8876;
17'hb0d2:	data_out=16'h8a00;
17'hb0d3:	data_out=16'h8c6;
17'hb0d4:	data_out=16'h89a1;
17'hb0d5:	data_out=16'h7bf;
17'hb0d6:	data_out=16'h8a00;
17'hb0d7:	data_out=16'h8a00;
17'hb0d8:	data_out=16'h465;
17'hb0d9:	data_out=16'h8a00;
17'hb0da:	data_out=16'h9ff;
17'hb0db:	data_out=16'h8a00;
17'hb0dc:	data_out=16'h9fb;
17'hb0dd:	data_out=16'h89a3;
17'hb0de:	data_out=16'h84bf;
17'hb0df:	data_out=16'h89e9;
17'hb0e0:	data_out=16'h89fe;
17'hb0e1:	data_out=16'h8a00;
17'hb0e2:	data_out=16'h9e9;
17'hb0e3:	data_out=16'h9f9;
17'hb0e4:	data_out=16'h8a00;
17'hb0e5:	data_out=16'h8873;
17'hb0e6:	data_out=16'h9d6;
17'hb0e7:	data_out=16'h898b;
17'hb0e8:	data_out=16'ha00;
17'hb0e9:	data_out=16'h884e;
17'hb0ea:	data_out=16'h9d1;
17'hb0eb:	data_out=16'h8a00;
17'hb0ec:	data_out=16'h8a00;
17'hb0ed:	data_out=16'h9f9;
17'hb0ee:	data_out=16'h9d2;
17'hb0ef:	data_out=16'h89b5;
17'hb0f0:	data_out=16'h9f9;
17'hb0f1:	data_out=16'h89ef;
17'hb0f2:	data_out=16'h8a00;
17'hb0f3:	data_out=16'h8a00;
17'hb0f4:	data_out=16'h8a00;
17'hb0f5:	data_out=16'h9c4;
17'hb0f6:	data_out=16'ha00;
17'hb0f7:	data_out=16'h89b2;
17'hb0f8:	data_out=16'ha00;
17'hb0f9:	data_out=16'h88fa;
17'hb0fa:	data_out=16'h9f6;
17'hb0fb:	data_out=16'ha00;
17'hb0fc:	data_out=16'h8a00;
17'hb0fd:	data_out=16'h8455;
17'hb0fe:	data_out=16'h9ff;
17'hb0ff:	data_out=16'h8a00;
17'hb100:	data_out=16'h8a00;
17'hb101:	data_out=16'h89c8;
17'hb102:	data_out=16'h28d;
17'hb103:	data_out=16'h85ba;
17'hb104:	data_out=16'h8a00;
17'hb105:	data_out=16'h89de;
17'hb106:	data_out=16'h9eb;
17'hb107:	data_out=16'h8a00;
17'hb108:	data_out=16'h892d;
17'hb109:	data_out=16'h601;
17'hb10a:	data_out=16'h89ba;
17'hb10b:	data_out=16'ha00;
17'hb10c:	data_out=16'h882d;
17'hb10d:	data_out=16'h8a00;
17'hb10e:	data_out=16'h9ed;
17'hb10f:	data_out=16'h89f8;
17'hb110:	data_out=16'h229;
17'hb111:	data_out=16'h1c0;
17'hb112:	data_out=16'h8a4;
17'hb113:	data_out=16'h8501;
17'hb114:	data_out=16'ha00;
17'hb115:	data_out=16'h8a00;
17'hb116:	data_out=16'h8a00;
17'hb117:	data_out=16'ha00;
17'hb118:	data_out=16'h8a00;
17'hb119:	data_out=16'ha00;
17'hb11a:	data_out=16'h89c2;
17'hb11b:	data_out=16'h9fb;
17'hb11c:	data_out=16'h88b4;
17'hb11d:	data_out=16'h8964;
17'hb11e:	data_out=16'h8557;
17'hb11f:	data_out=16'h97c;
17'hb120:	data_out=16'h899c;
17'hb121:	data_out=16'h9f2;
17'hb122:	data_out=16'h9f0;
17'hb123:	data_out=16'h89ff;
17'hb124:	data_out=16'h89ff;
17'hb125:	data_out=16'h89c0;
17'hb126:	data_out=16'h53;
17'hb127:	data_out=16'h8927;
17'hb128:	data_out=16'h9fb;
17'hb129:	data_out=16'h9f2;
17'hb12a:	data_out=16'h89ff;
17'hb12b:	data_out=16'ha00;
17'hb12c:	data_out=16'h8a00;
17'hb12d:	data_out=16'ha00;
17'hb12e:	data_out=16'h9e5;
17'hb12f:	data_out=16'h87ac;
17'hb130:	data_out=16'h8428;
17'hb131:	data_out=16'h89d4;
17'hb132:	data_out=16'h8997;
17'hb133:	data_out=16'h9ff;
17'hb134:	data_out=16'h89db;
17'hb135:	data_out=16'h89a1;
17'hb136:	data_out=16'h88f4;
17'hb137:	data_out=16'h9af;
17'hb138:	data_out=16'h8996;
17'hb139:	data_out=16'h6fe;
17'hb13a:	data_out=16'h88c9;
17'hb13b:	data_out=16'h89b3;
17'hb13c:	data_out=16'ha00;
17'hb13d:	data_out=16'h8a00;
17'hb13e:	data_out=16'h9fc;
17'hb13f:	data_out=16'h89e4;
17'hb140:	data_out=16'h8990;
17'hb141:	data_out=16'h89d7;
17'hb142:	data_out=16'h89e1;
17'hb143:	data_out=16'h9ec;
17'hb144:	data_out=16'h89d9;
17'hb145:	data_out=16'h8a00;
17'hb146:	data_out=16'ha00;
17'hb147:	data_out=16'h87f6;
17'hb148:	data_out=16'h9f8;
17'hb149:	data_out=16'h8985;
17'hb14a:	data_out=16'h877c;
17'hb14b:	data_out=16'h89df;
17'hb14c:	data_out=16'h89fd;
17'hb14d:	data_out=16'h9f6;
17'hb14e:	data_out=16'h9f5;
17'hb14f:	data_out=16'h89f7;
17'hb150:	data_out=16'h890b;
17'hb151:	data_out=16'h89f5;
17'hb152:	data_out=16'h89ff;
17'hb153:	data_out=16'h346;
17'hb154:	data_out=16'h896a;
17'hb155:	data_out=16'h996;
17'hb156:	data_out=16'h89ea;
17'hb157:	data_out=16'h89f3;
17'hb158:	data_out=16'h8477;
17'hb159:	data_out=16'h89b8;
17'hb15a:	data_out=16'h9f9;
17'hb15b:	data_out=16'h899e;
17'hb15c:	data_out=16'h860f;
17'hb15d:	data_out=16'h89a6;
17'hb15e:	data_out=16'h8652;
17'hb15f:	data_out=16'h89f5;
17'hb160:	data_out=16'h8001;
17'hb161:	data_out=16'h89f4;
17'hb162:	data_out=16'h9ff;
17'hb163:	data_out=16'ha00;
17'hb164:	data_out=16'h89e4;
17'hb165:	data_out=16'h9ff;
17'hb166:	data_out=16'h9fb;
17'hb167:	data_out=16'h9e5;
17'hb168:	data_out=16'h9f7;
17'hb169:	data_out=16'h8724;
17'hb16a:	data_out=16'h952;
17'hb16b:	data_out=16'h8955;
17'hb16c:	data_out=16'h8a00;
17'hb16d:	data_out=16'ha00;
17'hb16e:	data_out=16'h953;
17'hb16f:	data_out=16'h8974;
17'hb170:	data_out=16'h9b3;
17'hb171:	data_out=16'h89ff;
17'hb172:	data_out=16'h89ed;
17'hb173:	data_out=16'h89f8;
17'hb174:	data_out=16'h850f;
17'hb175:	data_out=16'h8936;
17'hb176:	data_out=16'ha00;
17'hb177:	data_out=16'h88a8;
17'hb178:	data_out=16'h9fb;
17'hb179:	data_out=16'h89d9;
17'hb17a:	data_out=16'ha00;
17'hb17b:	data_out=16'h9fc;
17'hb17c:	data_out=16'h8a00;
17'hb17d:	data_out=16'h52;
17'hb17e:	data_out=16'h958;
17'hb17f:	data_out=16'h8a00;
17'hb180:	data_out=16'h89fb;
17'hb181:	data_out=16'h89a6;
17'hb182:	data_out=16'h89f7;
17'hb183:	data_out=16'h867b;
17'hb184:	data_out=16'h8a00;
17'hb185:	data_out=16'h8a00;
17'hb186:	data_out=16'h555;
17'hb187:	data_out=16'h130;
17'hb188:	data_out=16'h89c1;
17'hb189:	data_out=16'h9ff;
17'hb18a:	data_out=16'h8968;
17'hb18b:	data_out=16'ha00;
17'hb18c:	data_out=16'h895a;
17'hb18d:	data_out=16'h8a00;
17'hb18e:	data_out=16'h89f1;
17'hb18f:	data_out=16'h89f9;
17'hb190:	data_out=16'ha00;
17'hb191:	data_out=16'ha00;
17'hb192:	data_out=16'h8a00;
17'hb193:	data_out=16'h86ce;
17'hb194:	data_out=16'h8111;
17'hb195:	data_out=16'h8a00;
17'hb196:	data_out=16'h8a00;
17'hb197:	data_out=16'h81fe;
17'hb198:	data_out=16'h8a00;
17'hb199:	data_out=16'ha00;
17'hb19a:	data_out=16'h8a00;
17'hb19b:	data_out=16'h8532;
17'hb19c:	data_out=16'h897c;
17'hb19d:	data_out=16'h9fe;
17'hb19e:	data_out=16'h8866;
17'hb19f:	data_out=16'h8838;
17'hb1a0:	data_out=16'h89cc;
17'hb1a1:	data_out=16'h89f0;
17'hb1a2:	data_out=16'ha00;
17'hb1a3:	data_out=16'h9fd;
17'hb1a4:	data_out=16'h9fd;
17'hb1a5:	data_out=16'h9de;
17'hb1a6:	data_out=16'h9ee;
17'hb1a7:	data_out=16'h88f4;
17'hb1a8:	data_out=16'h89d0;
17'hb1a9:	data_out=16'h9fa;
17'hb1aa:	data_out=16'h89e8;
17'hb1ab:	data_out=16'ha00;
17'hb1ac:	data_out=16'h8a00;
17'hb1ad:	data_out=16'ha00;
17'hb1ae:	data_out=16'h95;
17'hb1af:	data_out=16'h897a;
17'hb1b0:	data_out=16'h8483;
17'hb1b1:	data_out=16'h89dd;
17'hb1b2:	data_out=16'h89bb;
17'hb1b3:	data_out=16'h82ec;
17'hb1b4:	data_out=16'h8929;
17'hb1b5:	data_out=16'h89bb;
17'hb1b6:	data_out=16'h89ae;
17'hb1b7:	data_out=16'h8915;
17'hb1b8:	data_out=16'h89c2;
17'hb1b9:	data_out=16'h860a;
17'hb1ba:	data_out=16'h9fc;
17'hb1bb:	data_out=16'h89e8;
17'hb1bc:	data_out=16'ha00;
17'hb1bd:	data_out=16'h89eb;
17'hb1be:	data_out=16'h89cf;
17'hb1bf:	data_out=16'h8a00;
17'hb1c0:	data_out=16'h89d8;
17'hb1c1:	data_out=16'h89ec;
17'hb1c2:	data_out=16'h897f;
17'hb1c3:	data_out=16'h79f;
17'hb1c4:	data_out=16'h89e9;
17'hb1c5:	data_out=16'h8a00;
17'hb1c6:	data_out=16'ha00;
17'hb1c7:	data_out=16'h822c;
17'hb1c8:	data_out=16'h9ee;
17'hb1c9:	data_out=16'h9ed;
17'hb1ca:	data_out=16'h89b1;
17'hb1cb:	data_out=16'h89b0;
17'hb1cc:	data_out=16'h89fd;
17'hb1cd:	data_out=16'ha00;
17'hb1ce:	data_out=16'h870;
17'hb1cf:	data_out=16'h8441;
17'hb1d0:	data_out=16'h8988;
17'hb1d1:	data_out=16'h8a00;
17'hb1d2:	data_out=16'h357;
17'hb1d3:	data_out=16'h878c;
17'hb1d4:	data_out=16'h8992;
17'hb1d5:	data_out=16'h8290;
17'hb1d6:	data_out=16'h8912;
17'hb1d7:	data_out=16'h8996;
17'hb1d8:	data_out=16'h89e2;
17'hb1d9:	data_out=16'h89b4;
17'hb1da:	data_out=16'h661;
17'hb1db:	data_out=16'h89d8;
17'hb1dc:	data_out=16'h89bd;
17'hb1dd:	data_out=16'h89c1;
17'hb1de:	data_out=16'h88fb;
17'hb1df:	data_out=16'h89f3;
17'hb1e0:	data_out=16'h9db;
17'hb1e1:	data_out=16'h89fc;
17'hb1e2:	data_out=16'h253;
17'hb1e3:	data_out=16'h835f;
17'hb1e4:	data_out=16'h9f9;
17'hb1e5:	data_out=16'ha00;
17'hb1e6:	data_out=16'ha00;
17'hb1e7:	data_out=16'ha00;
17'hb1e8:	data_out=16'h89e7;
17'hb1e9:	data_out=16'h89e2;
17'hb1ea:	data_out=16'h89ef;
17'hb1eb:	data_out=16'h89cb;
17'hb1ec:	data_out=16'h8a00;
17'hb1ed:	data_out=16'h8353;
17'hb1ee:	data_out=16'h89ef;
17'hb1ef:	data_out=16'h89e8;
17'hb1f0:	data_out=16'h89f1;
17'hb1f1:	data_out=16'h8a00;
17'hb1f2:	data_out=16'h89e6;
17'hb1f3:	data_out=16'h89f2;
17'hb1f4:	data_out=16'h8553;
17'hb1f5:	data_out=16'h89fb;
17'hb1f6:	data_out=16'ha00;
17'hb1f7:	data_out=16'h899b;
17'hb1f8:	data_out=16'h8569;
17'hb1f9:	data_out=16'h89fb;
17'hb1fa:	data_out=16'h83d6;
17'hb1fb:	data_out=16'h89cf;
17'hb1fc:	data_out=16'h8a00;
17'hb1fd:	data_out=16'h89fd;
17'hb1fe:	data_out=16'h95d;
17'hb1ff:	data_out=16'h8a00;
17'hb200:	data_out=16'h8a00;
17'hb201:	data_out=16'h89eb;
17'hb202:	data_out=16'h8a00;
17'hb203:	data_out=16'h867b;
17'hb204:	data_out=16'h8a00;
17'hb205:	data_out=16'h8a00;
17'hb206:	data_out=16'h8f8;
17'hb207:	data_out=16'h228;
17'hb208:	data_out=16'h89e8;
17'hb209:	data_out=16'ha00;
17'hb20a:	data_out=16'h89b5;
17'hb20b:	data_out=16'ha00;
17'hb20c:	data_out=16'h9f6;
17'hb20d:	data_out=16'h8a00;
17'hb20e:	data_out=16'h89ff;
17'hb20f:	data_out=16'h89f9;
17'hb210:	data_out=16'h9f4;
17'hb211:	data_out=16'h89dd;
17'hb212:	data_out=16'h8a00;
17'hb213:	data_out=16'h9bd;
17'hb214:	data_out=16'h86a9;
17'hb215:	data_out=16'h8a00;
17'hb216:	data_out=16'h8a00;
17'hb217:	data_out=16'h8416;
17'hb218:	data_out=16'h8a00;
17'hb219:	data_out=16'ha00;
17'hb21a:	data_out=16'h8a00;
17'hb21b:	data_out=16'h87fa;
17'hb21c:	data_out=16'h89fc;
17'hb21d:	data_out=16'h8302;
17'hb21e:	data_out=16'h89ed;
17'hb21f:	data_out=16'h89f5;
17'hb220:	data_out=16'h8a00;
17'hb221:	data_out=16'h89ff;
17'hb222:	data_out=16'ha00;
17'hb223:	data_out=16'ha00;
17'hb224:	data_out=16'ha00;
17'hb225:	data_out=16'h9ab;
17'hb226:	data_out=16'h9ff;
17'hb227:	data_out=16'h89f5;
17'hb228:	data_out=16'h89ff;
17'hb229:	data_out=16'ha00;
17'hb22a:	data_out=16'h8983;
17'hb22b:	data_out=16'ha00;
17'hb22c:	data_out=16'h8a00;
17'hb22d:	data_out=16'ha00;
17'hb22e:	data_out=16'h32e;
17'hb22f:	data_out=16'h89e2;
17'hb230:	data_out=16'h893b;
17'hb231:	data_out=16'h8a00;
17'hb232:	data_out=16'h89c3;
17'hb233:	data_out=16'h89ba;
17'hb234:	data_out=16'h88c6;
17'hb235:	data_out=16'h8a00;
17'hb236:	data_out=16'h89ea;
17'hb237:	data_out=16'h89d9;
17'hb238:	data_out=16'h89f8;
17'hb239:	data_out=16'h89f5;
17'hb23a:	data_out=16'ha00;
17'hb23b:	data_out=16'h8a00;
17'hb23c:	data_out=16'ha00;
17'hb23d:	data_out=16'h8a00;
17'hb23e:	data_out=16'h89ff;
17'hb23f:	data_out=16'h8a00;
17'hb240:	data_out=16'h8a00;
17'hb241:	data_out=16'h8a00;
17'hb242:	data_out=16'h9fc;
17'hb243:	data_out=16'h8570;
17'hb244:	data_out=16'h8a00;
17'hb245:	data_out=16'h8a00;
17'hb246:	data_out=16'ha00;
17'hb247:	data_out=16'h682;
17'hb248:	data_out=16'h9dd;
17'hb249:	data_out=16'h9bf;
17'hb24a:	data_out=16'h89d0;
17'hb24b:	data_out=16'h9f6;
17'hb24c:	data_out=16'h9cb;
17'hb24d:	data_out=16'ha00;
17'hb24e:	data_out=16'h80d0;
17'hb24f:	data_out=16'ha00;
17'hb250:	data_out=16'h89f0;
17'hb251:	data_out=16'h8a00;
17'hb252:	data_out=16'h609;
17'hb253:	data_out=16'h89bc;
17'hb254:	data_out=16'h89fc;
17'hb255:	data_out=16'h88cf;
17'hb256:	data_out=16'h89fd;
17'hb257:	data_out=16'h89fa;
17'hb258:	data_out=16'h8a00;
17'hb259:	data_out=16'h89fa;
17'hb25a:	data_out=16'h8944;
17'hb25b:	data_out=16'h8a00;
17'hb25c:	data_out=16'h8a00;
17'hb25d:	data_out=16'h89eb;
17'hb25e:	data_out=16'h89b7;
17'hb25f:	data_out=16'h89fc;
17'hb260:	data_out=16'h9ff;
17'hb261:	data_out=16'h8a00;
17'hb262:	data_out=16'ha00;
17'hb263:	data_out=16'h8986;
17'hb264:	data_out=16'h9fe;
17'hb265:	data_out=16'h832;
17'hb266:	data_out=16'ha00;
17'hb267:	data_out=16'ha00;
17'hb268:	data_out=16'h89ff;
17'hb269:	data_out=16'h89eb;
17'hb26a:	data_out=16'h89ff;
17'hb26b:	data_out=16'h8a00;
17'hb26c:	data_out=16'h8a00;
17'hb26d:	data_out=16'h898a;
17'hb26e:	data_out=16'h89ff;
17'hb26f:	data_out=16'h8a00;
17'hb270:	data_out=16'h89ff;
17'hb271:	data_out=16'h8a00;
17'hb272:	data_out=16'h89fe;
17'hb273:	data_out=16'h89fe;
17'hb274:	data_out=16'h8953;
17'hb275:	data_out=16'h8a00;
17'hb276:	data_out=16'ha00;
17'hb277:	data_out=16'h8980;
17'hb278:	data_out=16'h851b;
17'hb279:	data_out=16'h8a00;
17'hb27a:	data_out=16'h88af;
17'hb27b:	data_out=16'h89ff;
17'hb27c:	data_out=16'h8a00;
17'hb27d:	data_out=16'h8a00;
17'hb27e:	data_out=16'h9fd;
17'hb27f:	data_out=16'h8a00;
17'hb280:	data_out=16'h8a00;
17'hb281:	data_out=16'h89fa;
17'hb282:	data_out=16'h8a00;
17'hb283:	data_out=16'h87d5;
17'hb284:	data_out=16'h8a00;
17'hb285:	data_out=16'h8a00;
17'hb286:	data_out=16'h9e9;
17'hb287:	data_out=16'h9f8;
17'hb288:	data_out=16'h8a00;
17'hb289:	data_out=16'ha00;
17'hb28a:	data_out=16'h89b6;
17'hb28b:	data_out=16'ha00;
17'hb28c:	data_out=16'ha00;
17'hb28d:	data_out=16'h8a00;
17'hb28e:	data_out=16'h8a00;
17'hb28f:	data_out=16'h8a00;
17'hb290:	data_out=16'hf5;
17'hb291:	data_out=16'h89ff;
17'hb292:	data_out=16'h8a00;
17'hb293:	data_out=16'h9df;
17'hb294:	data_out=16'h89dc;
17'hb295:	data_out=16'h8a00;
17'hb296:	data_out=16'h8a00;
17'hb297:	data_out=16'h8709;
17'hb298:	data_out=16'h8a00;
17'hb299:	data_out=16'ha00;
17'hb29a:	data_out=16'h8a00;
17'hb29b:	data_out=16'h89ff;
17'hb29c:	data_out=16'h8a00;
17'hb29d:	data_out=16'h8995;
17'hb29e:	data_out=16'h8a00;
17'hb29f:	data_out=16'h8a00;
17'hb2a0:	data_out=16'h8a00;
17'hb2a1:	data_out=16'h8a00;
17'hb2a2:	data_out=16'ha00;
17'hb2a3:	data_out=16'ha00;
17'hb2a4:	data_out=16'ha00;
17'hb2a5:	data_out=16'h9c7;
17'hb2a6:	data_out=16'ha00;
17'hb2a7:	data_out=16'h8a00;
17'hb2a8:	data_out=16'h8a00;
17'hb2a9:	data_out=16'ha00;
17'hb2aa:	data_out=16'h8997;
17'hb2ab:	data_out=16'ha00;
17'hb2ac:	data_out=16'h8a00;
17'hb2ad:	data_out=16'ha00;
17'hb2ae:	data_out=16'h31;
17'hb2af:	data_out=16'h8a00;
17'hb2b0:	data_out=16'h89a6;
17'hb2b1:	data_out=16'h8a00;
17'hb2b2:	data_out=16'h89c1;
17'hb2b3:	data_out=16'h8a00;
17'hb2b4:	data_out=16'h81ab;
17'hb2b5:	data_out=16'h8a00;
17'hb2b6:	data_out=16'h8a00;
17'hb2b7:	data_out=16'h8a00;
17'hb2b8:	data_out=16'h89ff;
17'hb2b9:	data_out=16'h8a00;
17'hb2ba:	data_out=16'ha00;
17'hb2bb:	data_out=16'h8a00;
17'hb2bc:	data_out=16'ha00;
17'hb2bd:	data_out=16'h8a00;
17'hb2be:	data_out=16'h8a00;
17'hb2bf:	data_out=16'h8a00;
17'hb2c0:	data_out=16'h8a00;
17'hb2c1:	data_out=16'h8a00;
17'hb2c2:	data_out=16'ha00;
17'hb2c3:	data_out=16'h86d4;
17'hb2c4:	data_out=16'h8a00;
17'hb2c5:	data_out=16'h8a00;
17'hb2c6:	data_out=16'ha00;
17'hb2c7:	data_out=16'h655;
17'hb2c8:	data_out=16'h78f;
17'hb2c9:	data_out=16'h9d9;
17'hb2ca:	data_out=16'h89f9;
17'hb2cb:	data_out=16'ha00;
17'hb2cc:	data_out=16'h9ff;
17'hb2cd:	data_out=16'ha00;
17'hb2ce:	data_out=16'h8958;
17'hb2cf:	data_out=16'ha00;
17'hb2d0:	data_out=16'h89fe;
17'hb2d1:	data_out=16'h8a00;
17'hb2d2:	data_out=16'h9ff;
17'hb2d3:	data_out=16'h8a00;
17'hb2d4:	data_out=16'h8a00;
17'hb2d5:	data_out=16'h89fd;
17'hb2d6:	data_out=16'h8a00;
17'hb2d7:	data_out=16'h8a00;
17'hb2d8:	data_out=16'h8a00;
17'hb2d9:	data_out=16'h8a00;
17'hb2da:	data_out=16'h8a00;
17'hb2db:	data_out=16'h8a00;
17'hb2dc:	data_out=16'h8a00;
17'hb2dd:	data_out=16'h8a00;
17'hb2de:	data_out=16'h89f1;
17'hb2df:	data_out=16'h8a00;
17'hb2e0:	data_out=16'ha00;
17'hb2e1:	data_out=16'h8a00;
17'hb2e2:	data_out=16'ha00;
17'hb2e3:	data_out=16'h8a00;
17'hb2e4:	data_out=16'ha00;
17'hb2e5:	data_out=16'h8171;
17'hb2e6:	data_out=16'ha00;
17'hb2e7:	data_out=16'ha00;
17'hb2e8:	data_out=16'h8a00;
17'hb2e9:	data_out=16'h8a00;
17'hb2ea:	data_out=16'h8a00;
17'hb2eb:	data_out=16'h8a00;
17'hb2ec:	data_out=16'h8a00;
17'hb2ed:	data_out=16'h8a00;
17'hb2ee:	data_out=16'h8a00;
17'hb2ef:	data_out=16'h8a00;
17'hb2f0:	data_out=16'h8a00;
17'hb2f1:	data_out=16'h8a00;
17'hb2f2:	data_out=16'h8a00;
17'hb2f3:	data_out=16'h8a00;
17'hb2f4:	data_out=16'h89b4;
17'hb2f5:	data_out=16'h8a00;
17'hb2f6:	data_out=16'ha00;
17'hb2f7:	data_out=16'h8925;
17'hb2f8:	data_out=16'h9f6;
17'hb2f9:	data_out=16'h8a00;
17'hb2fa:	data_out=16'h89fd;
17'hb2fb:	data_out=16'h8a00;
17'hb2fc:	data_out=16'h8a00;
17'hb2fd:	data_out=16'h8a00;
17'hb2fe:	data_out=16'ha00;
17'hb2ff:	data_out=16'h8a00;
17'hb300:	data_out=16'h8a00;
17'hb301:	data_out=16'h8a00;
17'hb302:	data_out=16'h8a00;
17'hb303:	data_out=16'h8876;
17'hb304:	data_out=16'h8a00;
17'hb305:	data_out=16'h8a00;
17'hb306:	data_out=16'ha00;
17'hb307:	data_out=16'ha00;
17'hb308:	data_out=16'h8a00;
17'hb309:	data_out=16'ha00;
17'hb30a:	data_out=16'h83f7;
17'hb30b:	data_out=16'ha00;
17'hb30c:	data_out=16'ha00;
17'hb30d:	data_out=16'h8a00;
17'hb30e:	data_out=16'h8a00;
17'hb30f:	data_out=16'h8a00;
17'hb310:	data_out=16'h89d7;
17'hb311:	data_out=16'h8a00;
17'hb312:	data_out=16'h8a00;
17'hb313:	data_out=16'h9f7;
17'hb314:	data_out=16'h89fd;
17'hb315:	data_out=16'h8a00;
17'hb316:	data_out=16'h8a00;
17'hb317:	data_out=16'h849e;
17'hb318:	data_out=16'h8a00;
17'hb319:	data_out=16'ha00;
17'hb31a:	data_out=16'h8a00;
17'hb31b:	data_out=16'h8a00;
17'hb31c:	data_out=16'h8a00;
17'hb31d:	data_out=16'h85f6;
17'hb31e:	data_out=16'h8a00;
17'hb31f:	data_out=16'h8a00;
17'hb320:	data_out=16'h8a00;
17'hb321:	data_out=16'h8a00;
17'hb322:	data_out=16'ha00;
17'hb323:	data_out=16'ha00;
17'hb324:	data_out=16'ha00;
17'hb325:	data_out=16'h848;
17'hb326:	data_out=16'ha00;
17'hb327:	data_out=16'h8a00;
17'hb328:	data_out=16'h8a00;
17'hb329:	data_out=16'ha00;
17'hb32a:	data_out=16'h8927;
17'hb32b:	data_out=16'h9ed;
17'hb32c:	data_out=16'h8a00;
17'hb32d:	data_out=16'ha00;
17'hb32e:	data_out=16'h443;
17'hb32f:	data_out=16'h8a00;
17'hb330:	data_out=16'h92f;
17'hb331:	data_out=16'h8a00;
17'hb332:	data_out=16'h794;
17'hb333:	data_out=16'h8a00;
17'hb334:	data_out=16'h9fe;
17'hb335:	data_out=16'h8a00;
17'hb336:	data_out=16'h8a00;
17'hb337:	data_out=16'h8a00;
17'hb338:	data_out=16'h8a00;
17'hb339:	data_out=16'h8a00;
17'hb33a:	data_out=16'ha00;
17'hb33b:	data_out=16'h8a00;
17'hb33c:	data_out=16'h9ff;
17'hb33d:	data_out=16'h8a00;
17'hb33e:	data_out=16'h8a00;
17'hb33f:	data_out=16'h8a00;
17'hb340:	data_out=16'h8a00;
17'hb341:	data_out=16'h8a00;
17'hb342:	data_out=16'ha00;
17'hb343:	data_out=16'h88d7;
17'hb344:	data_out=16'h8a00;
17'hb345:	data_out=16'h8a00;
17'hb346:	data_out=16'ha00;
17'hb347:	data_out=16'ha00;
17'hb348:	data_out=16'h613;
17'hb349:	data_out=16'h76c;
17'hb34a:	data_out=16'h8a00;
17'hb34b:	data_out=16'ha00;
17'hb34c:	data_out=16'ha00;
17'hb34d:	data_out=16'h9f8;
17'hb34e:	data_out=16'h89fa;
17'hb34f:	data_out=16'ha00;
17'hb350:	data_out=16'h8a00;
17'hb351:	data_out=16'h8a00;
17'hb352:	data_out=16'ha00;
17'hb353:	data_out=16'h8a00;
17'hb354:	data_out=16'h8a00;
17'hb355:	data_out=16'h89f1;
17'hb356:	data_out=16'h8a00;
17'hb357:	data_out=16'h8a00;
17'hb358:	data_out=16'h8a00;
17'hb359:	data_out=16'h8a00;
17'hb35a:	data_out=16'h8a00;
17'hb35b:	data_out=16'h8a00;
17'hb35c:	data_out=16'h8a00;
17'hb35d:	data_out=16'h8a00;
17'hb35e:	data_out=16'h89fe;
17'hb35f:	data_out=16'h8a00;
17'hb360:	data_out=16'ha00;
17'hb361:	data_out=16'h8a00;
17'hb362:	data_out=16'ha00;
17'hb363:	data_out=16'h8a00;
17'hb364:	data_out=16'ha00;
17'hb365:	data_out=16'h9f1;
17'hb366:	data_out=16'h9f0;
17'hb367:	data_out=16'ha00;
17'hb368:	data_out=16'h8a00;
17'hb369:	data_out=16'h8a00;
17'hb36a:	data_out=16'h8a00;
17'hb36b:	data_out=16'h8a00;
17'hb36c:	data_out=16'h8a00;
17'hb36d:	data_out=16'h8a00;
17'hb36e:	data_out=16'h8a00;
17'hb36f:	data_out=16'h89fe;
17'hb370:	data_out=16'h8a00;
17'hb371:	data_out=16'h8a00;
17'hb372:	data_out=16'h8a00;
17'hb373:	data_out=16'h8a00;
17'hb374:	data_out=16'h94b;
17'hb375:	data_out=16'h8a00;
17'hb376:	data_out=16'ha00;
17'hb377:	data_out=16'h8933;
17'hb378:	data_out=16'ha00;
17'hb379:	data_out=16'h8a00;
17'hb37a:	data_out=16'h8a00;
17'hb37b:	data_out=16'h8a00;
17'hb37c:	data_out=16'h8a00;
17'hb37d:	data_out=16'h8a00;
17'hb37e:	data_out=16'ha00;
17'hb37f:	data_out=16'h8a00;
17'hb380:	data_out=16'h8a00;
17'hb381:	data_out=16'h89ff;
17'hb382:	data_out=16'h8a00;
17'hb383:	data_out=16'h8965;
17'hb384:	data_out=16'h8a00;
17'hb385:	data_out=16'h8a00;
17'hb386:	data_out=16'ha00;
17'hb387:	data_out=16'ha00;
17'hb388:	data_out=16'h8a00;
17'hb389:	data_out=16'ha00;
17'hb38a:	data_out=16'h9f0;
17'hb38b:	data_out=16'ha00;
17'hb38c:	data_out=16'ha00;
17'hb38d:	data_out=16'h8a00;
17'hb38e:	data_out=16'h8a00;
17'hb38f:	data_out=16'h89f4;
17'hb390:	data_out=16'h89ef;
17'hb391:	data_out=16'h8a00;
17'hb392:	data_out=16'h8a00;
17'hb393:	data_out=16'h9a2;
17'hb394:	data_out=16'h89f1;
17'hb395:	data_out=16'h8a00;
17'hb396:	data_out=16'h8a00;
17'hb397:	data_out=16'h85bb;
17'hb398:	data_out=16'h8a00;
17'hb399:	data_out=16'ha00;
17'hb39a:	data_out=16'h8a00;
17'hb39b:	data_out=16'h8a00;
17'hb39c:	data_out=16'h8a00;
17'hb39d:	data_out=16'h86bd;
17'hb39e:	data_out=16'h8a00;
17'hb39f:	data_out=16'h89f7;
17'hb3a0:	data_out=16'h8a00;
17'hb3a1:	data_out=16'h8a00;
17'hb3a2:	data_out=16'ha00;
17'hb3a3:	data_out=16'ha00;
17'hb3a4:	data_out=16'ha00;
17'hb3a5:	data_out=16'h9af;
17'hb3a6:	data_out=16'ha00;
17'hb3a7:	data_out=16'h8a00;
17'hb3a8:	data_out=16'h8a00;
17'hb3a9:	data_out=16'ha00;
17'hb3aa:	data_out=16'h89ba;
17'hb3ab:	data_out=16'h89de;
17'hb3ac:	data_out=16'h8a00;
17'hb3ad:	data_out=16'ha00;
17'hb3ae:	data_out=16'h5f;
17'hb3af:	data_out=16'h8a00;
17'hb3b0:	data_out=16'ha00;
17'hb3b1:	data_out=16'h8a00;
17'hb3b2:	data_out=16'ha00;
17'hb3b3:	data_out=16'h8a00;
17'hb3b4:	data_out=16'h506;
17'hb3b5:	data_out=16'h8a00;
17'hb3b6:	data_out=16'h8a00;
17'hb3b7:	data_out=16'h8a00;
17'hb3b8:	data_out=16'h8a00;
17'hb3b9:	data_out=16'h8a00;
17'hb3ba:	data_out=16'h622;
17'hb3bb:	data_out=16'h230;
17'hb3bc:	data_out=16'h9ff;
17'hb3bd:	data_out=16'h8a00;
17'hb3be:	data_out=16'h8a00;
17'hb3bf:	data_out=16'h8a00;
17'hb3c0:	data_out=16'h8964;
17'hb3c1:	data_out=16'h8a00;
17'hb3c2:	data_out=16'ha00;
17'hb3c3:	data_out=16'h5f6;
17'hb3c4:	data_out=16'h8a00;
17'hb3c5:	data_out=16'h8a00;
17'hb3c6:	data_out=16'h9e4;
17'hb3c7:	data_out=16'hc2;
17'hb3c8:	data_out=16'h333;
17'hb3c9:	data_out=16'h92e;
17'hb3ca:	data_out=16'h8a00;
17'hb3cb:	data_out=16'ha00;
17'hb3cc:	data_out=16'ha00;
17'hb3cd:	data_out=16'h936;
17'hb3ce:	data_out=16'h8a00;
17'hb3cf:	data_out=16'ha00;
17'hb3d0:	data_out=16'h89e4;
17'hb3d1:	data_out=16'h8a00;
17'hb3d2:	data_out=16'ha00;
17'hb3d3:	data_out=16'h8a00;
17'hb3d4:	data_out=16'h8a00;
17'hb3d5:	data_out=16'h89e5;
17'hb3d6:	data_out=16'h8a00;
17'hb3d7:	data_out=16'h8a00;
17'hb3d8:	data_out=16'h8a00;
17'hb3d9:	data_out=16'h89ec;
17'hb3da:	data_out=16'h8a00;
17'hb3db:	data_out=16'h8a00;
17'hb3dc:	data_out=16'h8a00;
17'hb3dd:	data_out=16'h8a00;
17'hb3de:	data_out=16'h89f4;
17'hb3df:	data_out=16'h8a00;
17'hb3e0:	data_out=16'ha00;
17'hb3e1:	data_out=16'h89f1;
17'hb3e2:	data_out=16'ha00;
17'hb3e3:	data_out=16'h8a00;
17'hb3e4:	data_out=16'h9c3;
17'hb3e5:	data_out=16'ha00;
17'hb3e6:	data_out=16'h9dd;
17'hb3e7:	data_out=16'ha00;
17'hb3e8:	data_out=16'h8a00;
17'hb3e9:	data_out=16'h8a00;
17'hb3ea:	data_out=16'h8a00;
17'hb3eb:	data_out=16'h8a00;
17'hb3ec:	data_out=16'h8a00;
17'hb3ed:	data_out=16'h8a00;
17'hb3ee:	data_out=16'h8a00;
17'hb3ef:	data_out=16'ha00;
17'hb3f0:	data_out=16'h8a00;
17'hb3f1:	data_out=16'h89f5;
17'hb3f2:	data_out=16'h89fc;
17'hb3f3:	data_out=16'h8331;
17'hb3f4:	data_out=16'ha00;
17'hb3f5:	data_out=16'h8a00;
17'hb3f6:	data_out=16'ha00;
17'hb3f7:	data_out=16'h8920;
17'hb3f8:	data_out=16'ha00;
17'hb3f9:	data_out=16'h8a00;
17'hb3fa:	data_out=16'h8a00;
17'hb3fb:	data_out=16'h8a00;
17'hb3fc:	data_out=16'h8a00;
17'hb3fd:	data_out=16'h8a00;
17'hb3fe:	data_out=16'ha00;
17'hb3ff:	data_out=16'h8a00;
17'hb400:	data_out=16'h8a00;
17'hb401:	data_out=16'h89ff;
17'hb402:	data_out=16'h8a00;
17'hb403:	data_out=16'h89fc;
17'hb404:	data_out=16'h80b3;
17'hb405:	data_out=16'h8a00;
17'hb406:	data_out=16'ha00;
17'hb407:	data_out=16'ha00;
17'hb408:	data_out=16'h8a00;
17'hb409:	data_out=16'h82ab;
17'hb40a:	data_out=16'h9fc;
17'hb40b:	data_out=16'h83b;
17'hb40c:	data_out=16'h790;
17'hb40d:	data_out=16'h8a00;
17'hb40e:	data_out=16'h8a00;
17'hb40f:	data_out=16'h8a00;
17'hb410:	data_out=16'h89f9;
17'hb411:	data_out=16'h80b8;
17'hb412:	data_out=16'h8a00;
17'hb413:	data_out=16'h89f0;
17'hb414:	data_out=16'h8a00;
17'hb415:	data_out=16'h8a00;
17'hb416:	data_out=16'h8a00;
17'hb417:	data_out=16'h89f5;
17'hb418:	data_out=16'h8a00;
17'hb419:	data_out=16'ha00;
17'hb41a:	data_out=16'h729;
17'hb41b:	data_out=16'h8a00;
17'hb41c:	data_out=16'h8a00;
17'hb41d:	data_out=16'h87f6;
17'hb41e:	data_out=16'h8a00;
17'hb41f:	data_out=16'h89f2;
17'hb420:	data_out=16'h8a00;
17'hb421:	data_out=16'h89c1;
17'hb422:	data_out=16'ha00;
17'hb423:	data_out=16'h9fb;
17'hb424:	data_out=16'h9fb;
17'hb425:	data_out=16'h9ef;
17'hb426:	data_out=16'h837c;
17'hb427:	data_out=16'h8a00;
17'hb428:	data_out=16'h8a00;
17'hb429:	data_out=16'h8785;
17'hb42a:	data_out=16'h89fd;
17'hb42b:	data_out=16'h89fe;
17'hb42c:	data_out=16'h8a00;
17'hb42d:	data_out=16'ha00;
17'hb42e:	data_out=16'h898b;
17'hb42f:	data_out=16'h8a00;
17'hb430:	data_out=16'ha00;
17'hb431:	data_out=16'h8742;
17'hb432:	data_out=16'ha00;
17'hb433:	data_out=16'h8a00;
17'hb434:	data_out=16'h44f;
17'hb435:	data_out=16'h8a00;
17'hb436:	data_out=16'h8a00;
17'hb437:	data_out=16'h8a00;
17'hb438:	data_out=16'h364;
17'hb439:	data_out=16'h8a00;
17'hb43a:	data_out=16'h8998;
17'hb43b:	data_out=16'h83eb;
17'hb43c:	data_out=16'h89ee;
17'hb43d:	data_out=16'h8a00;
17'hb43e:	data_out=16'h8a00;
17'hb43f:	data_out=16'h8a00;
17'hb440:	data_out=16'h9fe;
17'hb441:	data_out=16'h8a00;
17'hb442:	data_out=16'ha00;
17'hb443:	data_out=16'h858e;
17'hb444:	data_out=16'h8a00;
17'hb445:	data_out=16'h8a00;
17'hb446:	data_out=16'h355;
17'hb447:	data_out=16'h8417;
17'hb448:	data_out=16'h89ea;
17'hb449:	data_out=16'h96a;
17'hb44a:	data_out=16'h89fa;
17'hb44b:	data_out=16'ha00;
17'hb44c:	data_out=16'ha00;
17'hb44d:	data_out=16'h912;
17'hb44e:	data_out=16'h8a00;
17'hb44f:	data_out=16'ha00;
17'hb450:	data_out=16'h89ee;
17'hb451:	data_out=16'h8a00;
17'hb452:	data_out=16'ha00;
17'hb453:	data_out=16'h8a00;
17'hb454:	data_out=16'h8a00;
17'hb455:	data_out=16'h89fb;
17'hb456:	data_out=16'h8a00;
17'hb457:	data_out=16'h8a00;
17'hb458:	data_out=16'h8a00;
17'hb459:	data_out=16'h41c;
17'hb45a:	data_out=16'h8a00;
17'hb45b:	data_out=16'h8a00;
17'hb45c:	data_out=16'h8a00;
17'hb45d:	data_out=16'h8a00;
17'hb45e:	data_out=16'h89fd;
17'hb45f:	data_out=16'h8a00;
17'hb460:	data_out=16'ha00;
17'hb461:	data_out=16'h89ea;
17'hb462:	data_out=16'h89db;
17'hb463:	data_out=16'h8a00;
17'hb464:	data_out=16'h2e6;
17'hb465:	data_out=16'ha00;
17'hb466:	data_out=16'h728;
17'hb467:	data_out=16'h8128;
17'hb468:	data_out=16'h89d5;
17'hb469:	data_out=16'h8a00;
17'hb46a:	data_out=16'h8a00;
17'hb46b:	data_out=16'h8a00;
17'hb46c:	data_out=16'h8a00;
17'hb46d:	data_out=16'h8a00;
17'hb46e:	data_out=16'h8a00;
17'hb46f:	data_out=16'ha00;
17'hb470:	data_out=16'h8a00;
17'hb471:	data_out=16'h89ff;
17'hb472:	data_out=16'h8228;
17'hb473:	data_out=16'h66f;
17'hb474:	data_out=16'ha00;
17'hb475:	data_out=16'h8a00;
17'hb476:	data_out=16'h5f8;
17'hb477:	data_out=16'h89e7;
17'hb478:	data_out=16'ha00;
17'hb479:	data_out=16'h8a00;
17'hb47a:	data_out=16'h8a00;
17'hb47b:	data_out=16'h8a00;
17'hb47c:	data_out=16'h8a00;
17'hb47d:	data_out=16'h8a00;
17'hb47e:	data_out=16'h376;
17'hb47f:	data_out=16'h8a00;
17'hb480:	data_out=16'h3e7;
17'hb481:	data_out=16'h82fe;
17'hb482:	data_out=16'h8a00;
17'hb483:	data_out=16'h8a00;
17'hb484:	data_out=16'ha00;
17'hb485:	data_out=16'h8997;
17'hb486:	data_out=16'h89fc;
17'hb487:	data_out=16'h8a00;
17'hb488:	data_out=16'h8a00;
17'hb489:	data_out=16'h89fd;
17'hb48a:	data_out=16'h3f2;
17'hb48b:	data_out=16'h89ff;
17'hb48c:	data_out=16'h8a00;
17'hb48d:	data_out=16'h8a00;
17'hb48e:	data_out=16'h218;
17'hb48f:	data_out=16'h8a00;
17'hb490:	data_out=16'h8a00;
17'hb491:	data_out=16'h9e8;
17'hb492:	data_out=16'h8a00;
17'hb493:	data_out=16'h8a00;
17'hb494:	data_out=16'h8a00;
17'hb495:	data_out=16'h877b;
17'hb496:	data_out=16'h8a00;
17'hb497:	data_out=16'h8a00;
17'hb498:	data_out=16'h8a00;
17'hb499:	data_out=16'ha00;
17'hb49a:	data_out=16'h9ff;
17'hb49b:	data_out=16'h8a00;
17'hb49c:	data_out=16'h59;
17'hb49d:	data_out=16'h86cf;
17'hb49e:	data_out=16'h8a00;
17'hb49f:	data_out=16'h89ff;
17'hb4a0:	data_out=16'h89c1;
17'hb4a1:	data_out=16'h189;
17'hb4a2:	data_out=16'h857f;
17'hb4a3:	data_out=16'h81c4;
17'hb4a4:	data_out=16'h81c4;
17'hb4a5:	data_out=16'h89fb;
17'hb4a6:	data_out=16'h8a00;
17'hb4a7:	data_out=16'h89e3;
17'hb4a8:	data_out=16'h93;
17'hb4a9:	data_out=16'h8a00;
17'hb4aa:	data_out=16'h8a00;
17'hb4ab:	data_out=16'h2e;
17'hb4ac:	data_out=16'h8a00;
17'hb4ad:	data_out=16'h42a;
17'hb4ae:	data_out=16'h89ff;
17'hb4af:	data_out=16'h8a00;
17'hb4b0:	data_out=16'h7b5;
17'hb4b1:	data_out=16'h4e3;
17'hb4b2:	data_out=16'h98b;
17'hb4b3:	data_out=16'h8a00;
17'hb4b4:	data_out=16'h9b3;
17'hb4b5:	data_out=16'h89fe;
17'hb4b6:	data_out=16'h8a00;
17'hb4b7:	data_out=16'h8a00;
17'hb4b8:	data_out=16'ha00;
17'hb4b9:	data_out=16'h8a00;
17'hb4ba:	data_out=16'h89fe;
17'hb4bb:	data_out=16'h8a00;
17'hb4bc:	data_out=16'h8a00;
17'hb4bd:	data_out=16'h83b1;
17'hb4be:	data_out=16'h8c;
17'hb4bf:	data_out=16'h8989;
17'hb4c0:	data_out=16'h8494;
17'hb4c1:	data_out=16'h8a00;
17'hb4c2:	data_out=16'h814b;
17'hb4c3:	data_out=16'h8a00;
17'hb4c4:	data_out=16'h89ee;
17'hb4c5:	data_out=16'h8981;
17'hb4c6:	data_out=16'h80e7;
17'hb4c7:	data_out=16'h89fe;
17'hb4c8:	data_out=16'h8a00;
17'hb4c9:	data_out=16'h89fe;
17'hb4ca:	data_out=16'h89ff;
17'hb4cb:	data_out=16'h8976;
17'hb4cc:	data_out=16'h8772;
17'hb4cd:	data_out=16'h8509;
17'hb4ce:	data_out=16'h8a00;
17'hb4cf:	data_out=16'h8949;
17'hb4d0:	data_out=16'h89fe;
17'hb4d1:	data_out=16'h8a00;
17'hb4d2:	data_out=16'h8a;
17'hb4d3:	data_out=16'h8a00;
17'hb4d4:	data_out=16'h89ef;
17'hb4d5:	data_out=16'h8a00;
17'hb4d6:	data_out=16'h85b7;
17'hb4d7:	data_out=16'h8412;
17'hb4d8:	data_out=16'h8a00;
17'hb4d9:	data_out=16'h50c;
17'hb4da:	data_out=16'h8a00;
17'hb4db:	data_out=16'ha00;
17'hb4dc:	data_out=16'h8a00;
17'hb4dd:	data_out=16'h89fc;
17'hb4de:	data_out=16'h89ff;
17'hb4df:	data_out=16'h858b;
17'hb4e0:	data_out=16'h8a00;
17'hb4e1:	data_out=16'h8098;
17'hb4e2:	data_out=16'h8a00;
17'hb4e3:	data_out=16'h8a00;
17'hb4e4:	data_out=16'hff;
17'hb4e5:	data_out=16'h8852;
17'hb4e6:	data_out=16'h8101;
17'hb4e7:	data_out=16'h88dd;
17'hb4e8:	data_out=16'hdd;
17'hb4e9:	data_out=16'h8a00;
17'hb4ea:	data_out=16'h31b;
17'hb4eb:	data_out=16'h6bb;
17'hb4ec:	data_out=16'h813a;
17'hb4ed:	data_out=16'h8a00;
17'hb4ee:	data_out=16'h31b;
17'hb4ef:	data_out=16'h88fc;
17'hb4f0:	data_out=16'h25e;
17'hb4f1:	data_out=16'h8a00;
17'hb4f2:	data_out=16'ha00;
17'hb4f3:	data_out=16'h9f5;
17'hb4f4:	data_out=16'h785;
17'hb4f5:	data_out=16'h8803;
17'hb4f6:	data_out=16'h8421;
17'hb4f7:	data_out=16'h8a00;
17'hb4f8:	data_out=16'h86a9;
17'hb4f9:	data_out=16'h8a00;
17'hb4fa:	data_out=16'h8a00;
17'hb4fb:	data_out=16'h8a;
17'hb4fc:	data_out=16'h86eb;
17'hb4fd:	data_out=16'h89f3;
17'hb4fe:	data_out=16'h89fd;
17'hb4ff:	data_out=16'h851b;
17'hb500:	data_out=16'ha00;
17'hb501:	data_out=16'h6af;
17'hb502:	data_out=16'h8708;
17'hb503:	data_out=16'h8878;
17'hb504:	data_out=16'h23d;
17'hb505:	data_out=16'h818a;
17'hb506:	data_out=16'h86f5;
17'hb507:	data_out=16'h8a00;
17'hb508:	data_out=16'h89d5;
17'hb509:	data_out=16'h8a00;
17'hb50a:	data_out=16'h72d;
17'hb50b:	data_out=16'h89ff;
17'hb50c:	data_out=16'h8a00;
17'hb50d:	data_out=16'h8a00;
17'hb50e:	data_out=16'h179;
17'hb50f:	data_out=16'h8a00;
17'hb510:	data_out=16'h8a00;
17'hb511:	data_out=16'h2a4;
17'hb512:	data_out=16'h89ff;
17'hb513:	data_out=16'h89ff;
17'hb514:	data_out=16'h8590;
17'hb515:	data_out=16'h15b;
17'hb516:	data_out=16'h867c;
17'hb517:	data_out=16'h89b2;
17'hb518:	data_out=16'h8213;
17'hb519:	data_out=16'h1cc;
17'hb51a:	data_out=16'h8040;
17'hb51b:	data_out=16'h8a00;
17'hb51c:	data_out=16'h814;
17'hb51d:	data_out=16'h24c;
17'hb51e:	data_out=16'h8729;
17'hb51f:	data_out=16'h8683;
17'hb520:	data_out=16'h893;
17'hb521:	data_out=16'h137;
17'hb522:	data_out=16'h82c2;
17'hb523:	data_out=16'h801b;
17'hb524:	data_out=16'h8018;
17'hb525:	data_out=16'h88cb;
17'hb526:	data_out=16'h8a00;
17'hb527:	data_out=16'hf3;
17'hb528:	data_out=16'h75;
17'hb529:	data_out=16'h8562;
17'hb52a:	data_out=16'h89ff;
17'hb52b:	data_out=16'h732;
17'hb52c:	data_out=16'h8573;
17'hb52d:	data_out=16'h8063;
17'hb52e:	data_out=16'h89ff;
17'hb52f:	data_out=16'h84c4;
17'hb530:	data_out=16'h8412;
17'hb531:	data_out=16'h7cb;
17'hb532:	data_out=16'h831f;
17'hb533:	data_out=16'h8424;
17'hb534:	data_out=16'h9e0;
17'hb535:	data_out=16'h8948;
17'hb536:	data_out=16'h89f8;
17'hb537:	data_out=16'h8790;
17'hb538:	data_out=16'ha00;
17'hb539:	data_out=16'h8352;
17'hb53a:	data_out=16'h8a00;
17'hb53b:	data_out=16'h84a2;
17'hb53c:	data_out=16'h874d;
17'hb53d:	data_out=16'h8b7;
17'hb53e:	data_out=16'h5b;
17'hb53f:	data_out=16'h817e;
17'hb540:	data_out=16'h874a;
17'hb541:	data_out=16'h89ff;
17'hb542:	data_out=16'h8889;
17'hb543:	data_out=16'h8a00;
17'hb544:	data_out=16'h8144;
17'hb545:	data_out=16'h113;
17'hb546:	data_out=16'h370;
17'hb547:	data_out=16'h89f4;
17'hb548:	data_out=16'h8a00;
17'hb549:	data_out=16'h8988;
17'hb54a:	data_out=16'h89fc;
17'hb54b:	data_out=16'h8a00;
17'hb54c:	data_out=16'h8867;
17'hb54d:	data_out=16'h8273;
17'hb54e:	data_out=16'h8a00;
17'hb54f:	data_out=16'h87a7;
17'hb550:	data_out=16'h880a;
17'hb551:	data_out=16'h893c;
17'hb552:	data_out=16'h47;
17'hb553:	data_out=16'h850b;
17'hb554:	data_out=16'h365;
17'hb555:	data_out=16'h8a00;
17'hb556:	data_out=16'h812c;
17'hb557:	data_out=16'h8093;
17'hb558:	data_out=16'h87bf;
17'hb559:	data_out=16'h820c;
17'hb55a:	data_out=16'h87c6;
17'hb55b:	data_out=16'ha00;
17'hb55c:	data_out=16'h82ec;
17'hb55d:	data_out=16'h8398;
17'hb55e:	data_out=16'h85ee;
17'hb55f:	data_out=16'h8052;
17'hb560:	data_out=16'h8961;
17'hb561:	data_out=16'h6b0;
17'hb562:	data_out=16'h89ff;
17'hb563:	data_out=16'h84c1;
17'hb564:	data_out=16'h766;
17'hb565:	data_out=16'h89e1;
17'hb566:	data_out=16'h84b7;
17'hb567:	data_out=16'h8701;
17'hb568:	data_out=16'he9;
17'hb569:	data_out=16'h8a00;
17'hb56a:	data_out=16'h1f4;
17'hb56b:	data_out=16'h226;
17'hb56c:	data_out=16'h5ff;
17'hb56d:	data_out=16'h847b;
17'hb56e:	data_out=16'h1e8;
17'hb56f:	data_out=16'h88f5;
17'hb570:	data_out=16'h19f;
17'hb571:	data_out=16'h89ff;
17'hb572:	data_out=16'h87c;
17'hb573:	data_out=16'h5fc;
17'hb574:	data_out=16'h8460;
17'hb575:	data_out=16'h828c;
17'hb576:	data_out=16'h80ce;
17'hb577:	data_out=16'h8a00;
17'hb578:	data_out=16'h86b6;
17'hb579:	data_out=16'h89ff;
17'hb57a:	data_out=16'h85f7;
17'hb57b:	data_out=16'h43;
17'hb57c:	data_out=16'h80c5;
17'hb57d:	data_out=16'h8962;
17'hb57e:	data_out=16'h8a00;
17'hb57f:	data_out=16'h81b4;
17'hb580:	data_out=16'h23c;
17'hb581:	data_out=16'h1a8;
17'hb582:	data_out=16'h8063;
17'hb583:	data_out=16'h7a;
17'hb584:	data_out=16'h806f;
17'hb585:	data_out=16'h802b;
17'hb586:	data_out=16'h8068;
17'hb587:	data_out=16'h80b1;
17'hb588:	data_out=16'h46;
17'hb589:	data_out=16'hf;
17'hb58a:	data_out=16'h7b;
17'hb58b:	data_out=16'h8039;
17'hb58c:	data_out=16'h8206;
17'hb58d:	data_out=16'h63;
17'hb58e:	data_out=16'h8026;
17'hb58f:	data_out=16'h2b;
17'hb590:	data_out=16'h7c;
17'hb591:	data_out=16'h8019;
17'hb592:	data_out=16'h1d;
17'hb593:	data_out=16'h6c;
17'hb594:	data_out=16'h117;
17'hb595:	data_out=16'hc8;
17'hb596:	data_out=16'h6c;
17'hb597:	data_out=16'h103;
17'hb598:	data_out=16'h8076;
17'hb599:	data_out=16'h806f;
17'hb59a:	data_out=16'h80d0;
17'hb59b:	data_out=16'h17b;
17'hb59c:	data_out=16'h126;
17'hb59d:	data_out=16'h19d;
17'hb59e:	data_out=16'h138;
17'hb59f:	data_out=16'h80ed;
17'hb5a0:	data_out=16'h2ea;
17'hb5a1:	data_out=16'h8026;
17'hb5a2:	data_out=16'hc8;
17'hb5a3:	data_out=16'h810d;
17'hb5a4:	data_out=16'h8114;
17'hb5a5:	data_out=16'h8013;
17'hb5a6:	data_out=16'h8095;
17'hb5a7:	data_out=16'h1bc;
17'hb5a8:	data_out=16'h802c;
17'hb5a9:	data_out=16'h55;
17'hb5aa:	data_out=16'h8041;
17'hb5ab:	data_out=16'h274;
17'hb5ac:	data_out=16'h8009;
17'hb5ad:	data_out=16'h6e;
17'hb5ae:	data_out=16'h801d;
17'hb5af:	data_out=16'h225;
17'hb5b0:	data_out=16'h80e9;
17'hb5b1:	data_out=16'h135;
17'hb5b2:	data_out=16'h80d4;
17'hb5b3:	data_out=16'h147;
17'hb5b4:	data_out=16'h124;
17'hb5b5:	data_out=16'h8151;
17'hb5b6:	data_out=16'hb3;
17'hb5b7:	data_out=16'h802b;
17'hb5b8:	data_out=16'h1a9;
17'hb5b9:	data_out=16'h103;
17'hb5ba:	data_out=16'h58;
17'hb5bb:	data_out=16'h8069;
17'hb5bc:	data_out=16'h78;
17'hb5bd:	data_out=16'h1b3;
17'hb5be:	data_out=16'h803b;
17'hb5bf:	data_out=16'h806c;
17'hb5c0:	data_out=16'h8051;
17'hb5c1:	data_out=16'h7e;
17'hb5c2:	data_out=16'h8063;
17'hb5c3:	data_out=16'h80ea;
17'hb5c4:	data_out=16'h28;
17'hb5c5:	data_out=16'h7b;
17'hb5c6:	data_out=16'hef;
17'hb5c7:	data_out=16'h803e;
17'hb5c8:	data_out=16'h8006;
17'hb5c9:	data_out=16'h5;
17'hb5ca:	data_out=16'h80d2;
17'hb5cb:	data_out=16'h80b2;
17'hb5cc:	data_out=16'h8041;
17'hb5cd:	data_out=16'h12d;
17'hb5ce:	data_out=16'h3b;
17'hb5cf:	data_out=16'h805b;
17'hb5d0:	data_out=16'h8053;
17'hb5d1:	data_out=16'h804d;
17'hb5d2:	data_out=16'h80d4;
17'hb5d3:	data_out=16'h279;
17'hb5d4:	data_out=16'h258;
17'hb5d5:	data_out=16'h8130;
17'hb5d6:	data_out=16'h2d;
17'hb5d7:	data_out=16'h8007;
17'hb5d8:	data_out=16'h80dd;
17'hb5d9:	data_out=16'h8012;
17'hb5da:	data_out=16'h97;
17'hb5db:	data_out=16'h802c;
17'hb5dc:	data_out=16'he2;
17'hb5dd:	data_out=16'hf1;
17'hb5de:	data_out=16'h1cb;
17'hb5df:	data_out=16'h5a;
17'hb5e0:	data_out=16'h80c0;
17'hb5e1:	data_out=16'h60;
17'hb5e2:	data_out=16'h18;
17'hb5e3:	data_out=16'h13d;
17'hb5e4:	data_out=16'h125;
17'hb5e5:	data_out=16'h800f;
17'hb5e6:	data_out=16'h80cb;
17'hb5e7:	data_out=16'h8026;
17'hb5e8:	data_out=16'h8034;
17'hb5e9:	data_out=16'h8023;
17'hb5ea:	data_out=16'h8021;
17'hb5eb:	data_out=16'h4d;
17'hb5ec:	data_out=16'h229;
17'hb5ed:	data_out=16'h149;
17'hb5ee:	data_out=16'h8028;
17'hb5ef:	data_out=16'h1;
17'hb5f0:	data_out=16'h8030;
17'hb5f1:	data_out=16'h812b;
17'hb5f2:	data_out=16'h801c;
17'hb5f3:	data_out=16'h8b;
17'hb5f4:	data_out=16'h80f0;
17'hb5f5:	data_out=16'h80fd;
17'hb5f6:	data_out=16'h9b;
17'hb5f7:	data_out=16'h80b7;
17'hb5f8:	data_out=16'h8052;
17'hb5f9:	data_out=16'h8072;
17'hb5fa:	data_out=16'h130;
17'hb5fb:	data_out=16'h803f;
17'hb5fc:	data_out=16'h8038;
17'hb5fd:	data_out=16'h80d5;
17'hb5fe:	data_out=16'h38;
17'hb5ff:	data_out=16'h80a1;
17'hb600:	data_out=16'h1;
17'hb601:	data_out=16'h9;
17'hb602:	data_out=16'h8000;
17'hb603:	data_out=16'h7;
17'hb604:	data_out=16'h8001;
17'hb605:	data_out=16'hb;
17'hb606:	data_out=16'h9;
17'hb607:	data_out=16'h4;
17'hb608:	data_out=16'h7;
17'hb609:	data_out=16'h7;
17'hb60a:	data_out=16'h4;
17'hb60b:	data_out=16'h8;
17'hb60c:	data_out=16'hc;
17'hb60d:	data_out=16'hc;
17'hb60e:	data_out=16'h7;
17'hb60f:	data_out=16'h8005;
17'hb610:	data_out=16'h8;
17'hb611:	data_out=16'h0;
17'hb612:	data_out=16'hb;
17'hb613:	data_out=16'h5;
17'hb614:	data_out=16'h6;
17'hb615:	data_out=16'h8004;
17'hb616:	data_out=16'h5;
17'hb617:	data_out=16'h1;
17'hb618:	data_out=16'h2;
17'hb619:	data_out=16'h1;
17'hb61a:	data_out=16'h6;
17'hb61b:	data_out=16'hc;
17'hb61c:	data_out=16'h6;
17'hb61d:	data_out=16'hc;
17'hb61e:	data_out=16'h2;
17'hb61f:	data_out=16'hd;
17'hb620:	data_out=16'h6;
17'hb621:	data_out=16'h4;
17'hb622:	data_out=16'h7;
17'hb623:	data_out=16'h7;
17'hb624:	data_out=16'h3;
17'hb625:	data_out=16'h5;
17'hb626:	data_out=16'h8002;
17'hb627:	data_out=16'h8000;
17'hb628:	data_out=16'h8004;
17'hb629:	data_out=16'h5;
17'hb62a:	data_out=16'hf;
17'hb62b:	data_out=16'h8006;
17'hb62c:	data_out=16'h5;
17'hb62d:	data_out=16'ha;
17'hb62e:	data_out=16'h8002;
17'hb62f:	data_out=16'h8002;
17'hb630:	data_out=16'h8003;
17'hb631:	data_out=16'hc;
17'hb632:	data_out=16'hb;
17'hb633:	data_out=16'h6;
17'hb634:	data_out=16'hd;
17'hb635:	data_out=16'h4;
17'hb636:	data_out=16'h8004;
17'hb637:	data_out=16'h3;
17'hb638:	data_out=16'h6;
17'hb639:	data_out=16'h4;
17'hb63a:	data_out=16'h2;
17'hb63b:	data_out=16'h2;
17'hb63c:	data_out=16'h2;
17'hb63d:	data_out=16'hb;
17'hb63e:	data_out=16'h8002;
17'hb63f:	data_out=16'h8005;
17'hb640:	data_out=16'h5;
17'hb641:	data_out=16'hb;
17'hb642:	data_out=16'ha;
17'hb643:	data_out=16'hb;
17'hb644:	data_out=16'h5;
17'hb645:	data_out=16'ha;
17'hb646:	data_out=16'h8004;
17'hb647:	data_out=16'h7;
17'hb648:	data_out=16'h3;
17'hb649:	data_out=16'h8001;
17'hb64a:	data_out=16'ha;
17'hb64b:	data_out=16'hd;
17'hb64c:	data_out=16'hf;
17'hb64d:	data_out=16'h7;
17'hb64e:	data_out=16'h8001;
17'hb64f:	data_out=16'hf;
17'hb650:	data_out=16'h6;
17'hb651:	data_out=16'hb;
17'hb652:	data_out=16'h5;
17'hb653:	data_out=16'h4;
17'hb654:	data_out=16'h8002;
17'hb655:	data_out=16'h8;
17'hb656:	data_out=16'hd;
17'hb657:	data_out=16'hc;
17'hb658:	data_out=16'h1;
17'hb659:	data_out=16'h2;
17'hb65a:	data_out=16'h8002;
17'hb65b:	data_out=16'h7;
17'hb65c:	data_out=16'h8004;
17'hb65d:	data_out=16'h4;
17'hb65e:	data_out=16'h7;
17'hb65f:	data_out=16'h3;
17'hb660:	data_out=16'h5;
17'hb661:	data_out=16'h4;
17'hb662:	data_out=16'h1;
17'hb663:	data_out=16'h9;
17'hb664:	data_out=16'h2;
17'hb665:	data_out=16'h7;
17'hb666:	data_out=16'h3;
17'hb667:	data_out=16'h9;
17'hb668:	data_out=16'h6;
17'hb669:	data_out=16'h8003;
17'hb66a:	data_out=16'h3;
17'hb66b:	data_out=16'h8;
17'hb66c:	data_out=16'hc;
17'hb66d:	data_out=16'h5;
17'hb66e:	data_out=16'h4;
17'hb66f:	data_out=16'h1;
17'hb670:	data_out=16'h2;
17'hb671:	data_out=16'h1;
17'hb672:	data_out=16'hc;
17'hb673:	data_out=16'h8;
17'hb674:	data_out=16'h8004;
17'hb675:	data_out=16'h9;
17'hb676:	data_out=16'h6;
17'hb677:	data_out=16'h3;
17'hb678:	data_out=16'h8004;
17'hb679:	data_out=16'hd;
17'hb67a:	data_out=16'hc;
17'hb67b:	data_out=16'h8004;
17'hb67c:	data_out=16'h8001;
17'hb67d:	data_out=16'h7;
17'hb67e:	data_out=16'h7;
17'hb67f:	data_out=16'hc;
17'hb680:	data_out=16'h282;
17'hb681:	data_out=16'h274;
17'hb682:	data_out=16'h124;
17'hb683:	data_out=16'h2d;
17'hb684:	data_out=16'h84ae;
17'hb685:	data_out=16'h8426;
17'hb686:	data_out=16'h84eb;
17'hb687:	data_out=16'h8246;
17'hb688:	data_out=16'hdf;
17'hb689:	data_out=16'h80da;
17'hb68a:	data_out=16'h804e;
17'hb68b:	data_out=16'h8097;
17'hb68c:	data_out=16'h82b2;
17'hb68d:	data_out=16'h6b;
17'hb68e:	data_out=16'h80ea;
17'hb68f:	data_out=16'h12;
17'hb690:	data_out=16'h174;
17'hb691:	data_out=16'h84d9;
17'hb692:	data_out=16'h345;
17'hb693:	data_out=16'h80cf;
17'hb694:	data_out=16'h1f9;
17'hb695:	data_out=16'h81fd;
17'hb696:	data_out=16'h820d;
17'hb697:	data_out=16'h30f;
17'hb698:	data_out=16'h80c7;
17'hb699:	data_out=16'h81e7;
17'hb69a:	data_out=16'h8539;
17'hb69b:	data_out=16'h341;
17'hb69c:	data_out=16'h830c;
17'hb69d:	data_out=16'h25a;
17'hb69e:	data_out=16'h30f;
17'hb69f:	data_out=16'h858f;
17'hb6a0:	data_out=16'h47d;
17'hb6a1:	data_out=16'h80e2;
17'hb6a2:	data_out=16'h39f;
17'hb6a3:	data_out=16'h81bb;
17'hb6a4:	data_out=16'h81b8;
17'hb6a5:	data_out=16'h80ce;
17'hb6a6:	data_out=16'h8154;
17'hb6a7:	data_out=16'h2c6;
17'hb6a8:	data_out=16'h80f0;
17'hb6a9:	data_out=16'h1a4;
17'hb6aa:	data_out=16'h381;
17'hb6ab:	data_out=16'h21;
17'hb6ac:	data_out=16'h81e3;
17'hb6ad:	data_out=16'h4f3;
17'hb6ae:	data_out=16'h26d;
17'hb6af:	data_out=16'h526;
17'hb6b0:	data_out=16'h859f;
17'hb6b1:	data_out=16'h80df;
17'hb6b2:	data_out=16'h8587;
17'hb6b3:	data_out=16'h20b;
17'hb6b4:	data_out=16'h804f;
17'hb6b5:	data_out=16'h8549;
17'hb6b6:	data_out=16'h356;
17'hb6b7:	data_out=16'h122;
17'hb6b8:	data_out=16'h8323;
17'hb6b9:	data_out=16'h12f;
17'hb6ba:	data_out=16'h37d;
17'hb6bb:	data_out=16'h8460;
17'hb6bc:	data_out=16'h34e;
17'hb6bd:	data_out=16'h818e;
17'hb6be:	data_out=16'h80e2;
17'hb6bf:	data_out=16'h84fa;
17'hb6c0:	data_out=16'h8356;
17'hb6c1:	data_out=16'h14f;
17'hb6c2:	data_out=16'h3fb;
17'hb6c3:	data_out=16'h859c;
17'hb6c4:	data_out=16'h8436;
17'hb6c5:	data_out=16'h822c;
17'hb6c6:	data_out=16'h267;
17'hb6c7:	data_out=16'hba;
17'hb6c8:	data_out=16'h259;
17'hb6c9:	data_out=16'h8142;
17'hb6ca:	data_out=16'h8109;
17'hb6cb:	data_out=16'h2b3;
17'hb6cc:	data_out=16'h175;
17'hb6cd:	data_out=16'h407;
17'hb6ce:	data_out=16'h256;
17'hb6cf:	data_out=16'h30;
17'hb6d0:	data_out=16'h835c;
17'hb6d1:	data_out=16'h8426;
17'hb6d2:	data_out=16'h8247;
17'hb6d3:	data_out=16'h617;
17'hb6d4:	data_out=16'h471;
17'hb6d5:	data_out=16'h804c;
17'hb6d6:	data_out=16'h81fd;
17'hb6d7:	data_out=16'h8207;
17'hb6d8:	data_out=16'h77;
17'hb6d9:	data_out=16'h8307;
17'hb6da:	data_out=16'h393;
17'hb6db:	data_out=16'h866c;
17'hb6dc:	data_out=16'h59;
17'hb6dd:	data_out=16'h339;
17'hb6de:	data_out=16'h488;
17'hb6df:	data_out=16'h1e0;
17'hb6e0:	data_out=16'h8163;
17'hb6e1:	data_out=16'h85e4;
17'hb6e2:	data_out=16'h5c;
17'hb6e3:	data_out=16'h21e;
17'hb6e4:	data_out=16'h81e2;
17'hb6e5:	data_out=16'h8228;
17'hb6e6:	data_out=16'h825e;
17'hb6e7:	data_out=16'h170;
17'hb6e8:	data_out=16'h80e4;
17'hb6e9:	data_out=16'hfa;
17'hb6ea:	data_out=16'h80f1;
17'hb6eb:	data_out=16'h84f6;
17'hb6ec:	data_out=16'h83a;
17'hb6ed:	data_out=16'h229;
17'hb6ee:	data_out=16'h80ed;
17'hb6ef:	data_out=16'h822f;
17'hb6f0:	data_out=16'h80e3;
17'hb6f1:	data_out=16'h38;
17'hb6f2:	data_out=16'h84e0;
17'hb6f3:	data_out=16'h84af;
17'hb6f4:	data_out=16'h85a0;
17'hb6f5:	data_out=16'h8504;
17'hb6f6:	data_out=16'h80d3;
17'hb6f7:	data_out=16'h845f;
17'hb6f8:	data_out=16'h85bc;
17'hb6f9:	data_out=16'h24a;
17'hb6fa:	data_out=16'h227;
17'hb6fb:	data_out=16'h80ec;
17'hb6fc:	data_out=16'h802c;
17'hb6fd:	data_out=16'h85e2;
17'hb6fe:	data_out=16'h8203;
17'hb6ff:	data_out=16'h8465;
17'hb700:	data_out=16'ha00;
17'hb701:	data_out=16'ha00;
17'hb702:	data_out=16'h3a4;
17'hb703:	data_out=16'h588;
17'hb704:	data_out=16'h8828;
17'hb705:	data_out=16'h8572;
17'hb706:	data_out=16'h8a00;
17'hb707:	data_out=16'h817d;
17'hb708:	data_out=16'h6f8;
17'hb709:	data_out=16'h822e;
17'hb70a:	data_out=16'h480;
17'hb70b:	data_out=16'h6d;
17'hb70c:	data_out=16'h8477;
17'hb70d:	data_out=16'h5d6;
17'hb70e:	data_out=16'h81e8;
17'hb70f:	data_out=16'h5da;
17'hb710:	data_out=16'h7ac;
17'hb711:	data_out=16'h87bf;
17'hb712:	data_out=16'h8f1;
17'hb713:	data_out=16'h291;
17'hb714:	data_out=16'h4de;
17'hb715:	data_out=16'h8123;
17'hb716:	data_out=16'h1f;
17'hb717:	data_out=16'h844;
17'hb718:	data_out=16'h8045;
17'hb719:	data_out=16'h8354;
17'hb71a:	data_out=16'h8916;
17'hb71b:	data_out=16'ha00;
17'hb71c:	data_out=16'h84de;
17'hb71d:	data_out=16'ha00;
17'hb71e:	data_out=16'ha00;
17'hb71f:	data_out=16'h89fd;
17'hb720:	data_out=16'ha00;
17'hb721:	data_out=16'h81e1;
17'hb722:	data_out=16'ha00;
17'hb723:	data_out=16'h8455;
17'hb724:	data_out=16'h8455;
17'hb725:	data_out=16'h31;
17'hb726:	data_out=16'h84a8;
17'hb727:	data_out=16'ha00;
17'hb728:	data_out=16'h81e1;
17'hb729:	data_out=16'h949;
17'hb72a:	data_out=16'ha00;
17'hb72b:	data_out=16'h360;
17'hb72c:	data_out=16'h8128;
17'hb72d:	data_out=16'ha00;
17'hb72e:	data_out=16'ha00;
17'hb72f:	data_out=16'ha00;
17'hb730:	data_out=16'h87a5;
17'hb731:	data_out=16'h5e8;
17'hb732:	data_out=16'h8742;
17'hb733:	data_out=16'h5ad;
17'hb734:	data_out=16'h365;
17'hb735:	data_out=16'h8812;
17'hb736:	data_out=16'ha00;
17'hb737:	data_out=16'h38d;
17'hb738:	data_out=16'h8157;
17'hb739:	data_out=16'h756;
17'hb73a:	data_out=16'h9fe;
17'hb73b:	data_out=16'h8740;
17'hb73c:	data_out=16'h9ec;
17'hb73d:	data_out=16'hd7;
17'hb73e:	data_out=16'h81db;
17'hb73f:	data_out=16'h8700;
17'hb740:	data_out=16'h88d9;
17'hb741:	data_out=16'h3c7;
17'hb742:	data_out=16'ha00;
17'hb743:	data_out=16'h8a00;
17'hb744:	data_out=16'h8673;
17'hb745:	data_out=16'h82ea;
17'hb746:	data_out=16'h80a;
17'hb747:	data_out=16'h2a2;
17'hb748:	data_out=16'ha00;
17'hb749:	data_out=16'h8146;
17'hb74a:	data_out=16'h2ed;
17'hb74b:	data_out=16'ha00;
17'hb74c:	data_out=16'h836;
17'hb74d:	data_out=16'ha00;
17'hb74e:	data_out=16'ha00;
17'hb74f:	data_out=16'h4a6;
17'hb750:	data_out=16'h89fc;
17'hb751:	data_out=16'h8974;
17'hb752:	data_out=16'h85f9;
17'hb753:	data_out=16'ha00;
17'hb754:	data_out=16'ha00;
17'hb755:	data_out=16'h8234;
17'hb756:	data_out=16'h8726;
17'hb757:	data_out=16'h86d7;
17'hb758:	data_out=16'h8061;
17'hb759:	data_out=16'h864f;
17'hb75a:	data_out=16'h9ff;
17'hb75b:	data_out=16'h89f8;
17'hb75c:	data_out=16'h89d;
17'hb75d:	data_out=16'ha00;
17'hb75e:	data_out=16'ha00;
17'hb75f:	data_out=16'h935;
17'hb760:	data_out=16'h82b2;
17'hb761:	data_out=16'h88e1;
17'hb762:	data_out=16'h260;
17'hb763:	data_out=16'h5e2;
17'hb764:	data_out=16'h818a;
17'hb765:	data_out=16'h3b;
17'hb766:	data_out=16'h852f;
17'hb767:	data_out=16'h471;
17'hb768:	data_out=16'h81e1;
17'hb769:	data_out=16'h69e;
17'hb76a:	data_out=16'h8209;
17'hb76b:	data_out=16'h87ac;
17'hb76c:	data_out=16'ha00;
17'hb76d:	data_out=16'h61f;
17'hb76e:	data_out=16'h8202;
17'hb76f:	data_out=16'h1d;
17'hb770:	data_out=16'h81ef;
17'hb771:	data_out=16'h1db;
17'hb772:	data_out=16'h8758;
17'hb773:	data_out=16'h8611;
17'hb774:	data_out=16'h87bb;
17'hb775:	data_out=16'h898e;
17'hb776:	data_out=16'h814c;
17'hb777:	data_out=16'h8957;
17'hb778:	data_out=16'h8a00;
17'hb779:	data_out=16'ha00;
17'hb77a:	data_out=16'h5ad;
17'hb77b:	data_out=16'h81d4;
17'hb77c:	data_out=16'h25c;
17'hb77d:	data_out=16'h89fe;
17'hb77e:	data_out=16'h8767;
17'hb77f:	data_out=16'h88a2;
17'hb780:	data_out=16'ha00;
17'hb781:	data_out=16'ha00;
17'hb782:	data_out=16'h604;
17'hb783:	data_out=16'hb0;
17'hb784:	data_out=16'h8a00;
17'hb785:	data_out=16'h8a00;
17'hb786:	data_out=16'h89fd;
17'hb787:	data_out=16'h89f9;
17'hb788:	data_out=16'ha00;
17'hb789:	data_out=16'h84c0;
17'hb78a:	data_out=16'h8744;
17'hb78b:	data_out=16'h3ef;
17'hb78c:	data_out=16'h89fe;
17'hb78d:	data_out=16'h739;
17'hb78e:	data_out=16'h84ab;
17'hb78f:	data_out=16'h7ee;
17'hb790:	data_out=16'h98e;
17'hb791:	data_out=16'h89f1;
17'hb792:	data_out=16'h9ff;
17'hb793:	data_out=16'h8074;
17'hb794:	data_out=16'h9b6;
17'hb795:	data_out=16'h8a00;
17'hb796:	data_out=16'h8a00;
17'hb797:	data_out=16'h9f4;
17'hb798:	data_out=16'h15c;
17'hb799:	data_out=16'h88ec;
17'hb79a:	data_out=16'h8a00;
17'hb79b:	data_out=16'h9f6;
17'hb79c:	data_out=16'h89d5;
17'hb79d:	data_out=16'h9ff;
17'hb79e:	data_out=16'h9f6;
17'hb79f:	data_out=16'h8a00;
17'hb7a0:	data_out=16'h9ff;
17'hb7a1:	data_out=16'h84b4;
17'hb7a2:	data_out=16'h9e0;
17'hb7a3:	data_out=16'h89f0;
17'hb7a4:	data_out=16'h89f2;
17'hb7a5:	data_out=16'h8532;
17'hb7a6:	data_out=16'h8a00;
17'hb7a7:	data_out=16'h9f5;
17'hb7a8:	data_out=16'h84de;
17'hb7a9:	data_out=16'h9fc;
17'hb7aa:	data_out=16'h9fb;
17'hb7ab:	data_out=16'h823;
17'hb7ac:	data_out=16'h8a00;
17'hb7ad:	data_out=16'ha00;
17'hb7ae:	data_out=16'h9d9;
17'hb7af:	data_out=16'ha00;
17'hb7b0:	data_out=16'h89f8;
17'hb7b1:	data_out=16'h8887;
17'hb7b2:	data_out=16'h8a00;
17'hb7b3:	data_out=16'h9fc;
17'hb7b4:	data_out=16'h4da;
17'hb7b5:	data_out=16'h8a00;
17'hb7b6:	data_out=16'ha00;
17'hb7b7:	data_out=16'h603;
17'hb7b8:	data_out=16'h80fa;
17'hb7b9:	data_out=16'h9fd;
17'hb7ba:	data_out=16'h972;
17'hb7bb:	data_out=16'h8a00;
17'hb7bc:	data_out=16'h9f7;
17'hb7bd:	data_out=16'h892d;
17'hb7be:	data_out=16'h84e0;
17'hb7bf:	data_out=16'h8a00;
17'hb7c0:	data_out=16'h8a00;
17'hb7c1:	data_out=16'h900;
17'hb7c2:	data_out=16'h94e;
17'hb7c3:	data_out=16'h8a00;
17'hb7c4:	data_out=16'h89ff;
17'hb7c5:	data_out=16'h8a00;
17'hb7c6:	data_out=16'ha00;
17'hb7c7:	data_out=16'h849d;
17'hb7c8:	data_out=16'ha00;
17'hb7c9:	data_out=16'h88ed;
17'hb7ca:	data_out=16'h82bf;
17'hb7cb:	data_out=16'h244;
17'hb7cc:	data_out=16'h558;
17'hb7cd:	data_out=16'ha00;
17'hb7ce:	data_out=16'ha00;
17'hb7cf:	data_out=16'h8104;
17'hb7d0:	data_out=16'h8a00;
17'hb7d1:	data_out=16'h89fb;
17'hb7d2:	data_out=16'h8a00;
17'hb7d3:	data_out=16'ha00;
17'hb7d4:	data_out=16'ha00;
17'hb7d5:	data_out=16'h595;
17'hb7d6:	data_out=16'h8a00;
17'hb7d7:	data_out=16'h8a00;
17'hb7d8:	data_out=16'h85e;
17'hb7d9:	data_out=16'h8a00;
17'hb7da:	data_out=16'h9fa;
17'hb7db:	data_out=16'h89fe;
17'hb7dc:	data_out=16'h871;
17'hb7dd:	data_out=16'ha00;
17'hb7de:	data_out=16'ha00;
17'hb7df:	data_out=16'ha00;
17'hb7e0:	data_out=16'h8a00;
17'hb7e1:	data_out=16'h8a00;
17'hb7e2:	data_out=16'h863;
17'hb7e3:	data_out=16'h9fe;
17'hb7e4:	data_out=16'h814e;
17'hb7e5:	data_out=16'h89f6;
17'hb7e6:	data_out=16'h89fe;
17'hb7e7:	data_out=16'h477;
17'hb7e8:	data_out=16'h84c5;
17'hb7e9:	data_out=16'h9fe;
17'hb7ea:	data_out=16'h84af;
17'hb7eb:	data_out=16'h8a00;
17'hb7ec:	data_out=16'ha00;
17'hb7ed:	data_out=16'h9fe;
17'hb7ee:	data_out=16'h84af;
17'hb7ef:	data_out=16'h8a00;
17'hb7f0:	data_out=16'h84ae;
17'hb7f1:	data_out=16'h80b3;
17'hb7f2:	data_out=16'h8a00;
17'hb7f3:	data_out=16'h8a00;
17'hb7f4:	data_out=16'h89f6;
17'hb7f5:	data_out=16'h8a00;
17'hb7f6:	data_out=16'h88f7;
17'hb7f7:	data_out=16'h89bf;
17'hb7f8:	data_out=16'h8a00;
17'hb7f9:	data_out=16'h9fb;
17'hb7fa:	data_out=16'h9fb;
17'hb7fb:	data_out=16'h84e1;
17'hb7fc:	data_out=16'h657;
17'hb7fd:	data_out=16'h89ff;
17'hb7fe:	data_out=16'h8a00;
17'hb7ff:	data_out=16'h89fe;
17'hb800:	data_out=16'h8916;
17'hb801:	data_out=16'h89f7;
17'hb802:	data_out=16'h966;
17'hb803:	data_out=16'h394;
17'hb804:	data_out=16'h8a00;
17'hb805:	data_out=16'h8a00;
17'hb806:	data_out=16'h89ff;
17'hb807:	data_out=16'h8833;
17'hb808:	data_out=16'ha00;
17'hb809:	data_out=16'h7bd;
17'hb80a:	data_out=16'h8a00;
17'hb80b:	data_out=16'h9f7;
17'hb80c:	data_out=16'h119;
17'hb80d:	data_out=16'h9fc;
17'hb80e:	data_out=16'h8042;
17'hb80f:	data_out=16'h974;
17'hb810:	data_out=16'h86b;
17'hb811:	data_out=16'h89fd;
17'hb812:	data_out=16'ha00;
17'hb813:	data_out=16'h48e;
17'hb814:	data_out=16'h9a8;
17'hb815:	data_out=16'h8a00;
17'hb816:	data_out=16'h89ff;
17'hb817:	data_out=16'h9ef;
17'hb818:	data_out=16'h483;
17'hb819:	data_out=16'h898d;
17'hb81a:	data_out=16'h8a00;
17'hb81b:	data_out=16'h9fe;
17'hb81c:	data_out=16'h88f7;
17'hb81d:	data_out=16'h89f1;
17'hb81e:	data_out=16'h8d8;
17'hb81f:	data_out=16'h89ff;
17'hb820:	data_out=16'h89f0;
17'hb821:	data_out=16'h21;
17'hb822:	data_out=16'h8a0;
17'hb823:	data_out=16'h81f3;
17'hb824:	data_out=16'h81ef;
17'hb825:	data_out=16'h84f9;
17'hb826:	data_out=16'h9f8;
17'hb827:	data_out=16'h89f0;
17'hb828:	data_out=16'h6e;
17'hb829:	data_out=16'h9fa;
17'hb82a:	data_out=16'h905;
17'hb82b:	data_out=16'ha00;
17'hb82c:	data_out=16'h8a00;
17'hb82d:	data_out=16'ha00;
17'hb82e:	data_out=16'h7e7;
17'hb82f:	data_out=16'h89ee;
17'hb830:	data_out=16'h89c9;
17'hb831:	data_out=16'h89ff;
17'hb832:	data_out=16'h8a00;
17'hb833:	data_out=16'h9b8;
17'hb834:	data_out=16'h89e7;
17'hb835:	data_out=16'h8a00;
17'hb836:	data_out=16'h9f4;
17'hb837:	data_out=16'h8e4;
17'hb838:	data_out=16'h89f0;
17'hb839:	data_out=16'h9d0;
17'hb83a:	data_out=16'h2ce;
17'hb83b:	data_out=16'h89fc;
17'hb83c:	data_out=16'h9e8;
17'hb83d:	data_out=16'h89ff;
17'hb83e:	data_out=16'h6d;
17'hb83f:	data_out=16'h8a00;
17'hb840:	data_out=16'h8a00;
17'hb841:	data_out=16'h9f7;
17'hb842:	data_out=16'h9f3;
17'hb843:	data_out=16'h8a00;
17'hb844:	data_out=16'h89fe;
17'hb845:	data_out=16'h8a00;
17'hb846:	data_out=16'ha00;
17'hb847:	data_out=16'h85ae;
17'hb848:	data_out=16'h93e;
17'hb849:	data_out=16'h8a00;
17'hb84a:	data_out=16'h894d;
17'hb84b:	data_out=16'h41b;
17'hb84c:	data_out=16'h866a;
17'hb84d:	data_out=16'h9f3;
17'hb84e:	data_out=16'ha00;
17'hb84f:	data_out=16'h89f6;
17'hb850:	data_out=16'h8a00;
17'hb851:	data_out=16'h9e7;
17'hb852:	data_out=16'h846f;
17'hb853:	data_out=16'h875e;
17'hb854:	data_out=16'h89df;
17'hb855:	data_out=16'h9e8;
17'hb856:	data_out=16'h89ff;
17'hb857:	data_out=16'h8a00;
17'hb858:	data_out=16'h9fa;
17'hb859:	data_out=16'h8a00;
17'hb85a:	data_out=16'h9fe;
17'hb85b:	data_out=16'h8a00;
17'hb85c:	data_out=16'h89fd;
17'hb85d:	data_out=16'h89f5;
17'hb85e:	data_out=16'h89f2;
17'hb85f:	data_out=16'h32a;
17'hb860:	data_out=16'h9fb;
17'hb861:	data_out=16'h8a00;
17'hb862:	data_out=16'h95f;
17'hb863:	data_out=16'h9cc;
17'hb864:	data_out=16'h87bd;
17'hb865:	data_out=16'h8a00;
17'hb866:	data_out=16'h89f5;
17'hb867:	data_out=16'h271;
17'hb868:	data_out=16'h4e;
17'hb869:	data_out=16'ha00;
17'hb86a:	data_out=16'h80a0;
17'hb86b:	data_out=16'h8a00;
17'hb86c:	data_out=16'h89d2;
17'hb86d:	data_out=16'h9c4;
17'hb86e:	data_out=16'h809e;
17'hb86f:	data_out=16'h8a00;
17'hb870:	data_out=16'h8069;
17'hb871:	data_out=16'h86ba;
17'hb872:	data_out=16'h8a00;
17'hb873:	data_out=16'h8a00;
17'hb874:	data_out=16'h89af;
17'hb875:	data_out=16'h8a00;
17'hb876:	data_out=16'h89fc;
17'hb877:	data_out=16'h8451;
17'hb878:	data_out=16'h8a00;
17'hb879:	data_out=16'ha00;
17'hb87a:	data_out=16'h9bd;
17'hb87b:	data_out=16'h6e;
17'hb87c:	data_out=16'h810d;
17'hb87d:	data_out=16'h8a00;
17'hb87e:	data_out=16'h2c7;
17'hb87f:	data_out=16'h8a00;
17'hb880:	data_out=16'h89fd;
17'hb881:	data_out=16'h8a00;
17'hb882:	data_out=16'h41e;
17'hb883:	data_out=16'h856b;
17'hb884:	data_out=16'h8a00;
17'hb885:	data_out=16'h8a00;
17'hb886:	data_out=16'h89fe;
17'hb887:	data_out=16'ha00;
17'hb888:	data_out=16'h926;
17'hb889:	data_out=16'h9e2;
17'hb88a:	data_out=16'h8a00;
17'hb88b:	data_out=16'h9ea;
17'hb88c:	data_out=16'ha00;
17'hb88d:	data_out=16'h9e9;
17'hb88e:	data_out=16'h22f;
17'hb88f:	data_out=16'h605;
17'hb890:	data_out=16'h851f;
17'hb891:	data_out=16'h8a00;
17'hb892:	data_out=16'h9aa;
17'hb893:	data_out=16'h9e7;
17'hb894:	data_out=16'h8a00;
17'hb895:	data_out=16'h8a00;
17'hb896:	data_out=16'h8a00;
17'hb897:	data_out=16'h2ff;
17'hb898:	data_out=16'h82cf;
17'hb899:	data_out=16'h8337;
17'hb89a:	data_out=16'h8a00;
17'hb89b:	data_out=16'h800d;
17'hb89c:	data_out=16'h8a00;
17'hb89d:	data_out=16'h8a00;
17'hb89e:	data_out=16'h8a00;
17'hb89f:	data_out=16'h8a00;
17'hb8a0:	data_out=16'h8a00;
17'hb8a1:	data_out=16'h2ed;
17'hb8a2:	data_out=16'h5b4;
17'hb8a3:	data_out=16'ha00;
17'hb8a4:	data_out=16'ha00;
17'hb8a5:	data_out=16'h8f1;
17'hb8a6:	data_out=16'h9fe;
17'hb8a7:	data_out=16'h8a00;
17'hb8a8:	data_out=16'h33b;
17'hb8a9:	data_out=16'h92a;
17'hb8aa:	data_out=16'h25c;
17'hb8ab:	data_out=16'h6a0;
17'hb8ac:	data_out=16'h8a00;
17'hb8ad:	data_out=16'ha00;
17'hb8ae:	data_out=16'h171;
17'hb8af:	data_out=16'h8a00;
17'hb8b0:	data_out=16'h866f;
17'hb8b1:	data_out=16'h8a00;
17'hb8b2:	data_out=16'h89f8;
17'hb8b3:	data_out=16'h8a00;
17'hb8b4:	data_out=16'h8a00;
17'hb8b5:	data_out=16'h8a00;
17'hb8b6:	data_out=16'h89fd;
17'hb8b7:	data_out=16'h759;
17'hb8b8:	data_out=16'h8a00;
17'hb8b9:	data_out=16'h8a00;
17'hb8ba:	data_out=16'h7bf;
17'hb8bb:	data_out=16'h89b0;
17'hb8bc:	data_out=16'h82b8;
17'hb8bd:	data_out=16'h8a00;
17'hb8be:	data_out=16'h33a;
17'hb8bf:	data_out=16'h8a00;
17'hb8c0:	data_out=16'h8a00;
17'hb8c1:	data_out=16'h7ce;
17'hb8c2:	data_out=16'ha00;
17'hb8c3:	data_out=16'h8a00;
17'hb8c4:	data_out=16'h8a00;
17'hb8c5:	data_out=16'h8a00;
17'hb8c6:	data_out=16'h9f9;
17'hb8c7:	data_out=16'h9ea;
17'hb8c8:	data_out=16'h89f6;
17'hb8c9:	data_out=16'h952;
17'hb8ca:	data_out=16'h82f4;
17'hb8cb:	data_out=16'ha00;
17'hb8cc:	data_out=16'h9fd;
17'hb8cd:	data_out=16'h6b0;
17'hb8ce:	data_out=16'h814a;
17'hb8cf:	data_out=16'ha00;
17'hb8d0:	data_out=16'h8a00;
17'hb8d1:	data_out=16'h9ab;
17'hb8d2:	data_out=16'ha00;
17'hb8d3:	data_out=16'h8a00;
17'hb8d4:	data_out=16'h8a00;
17'hb8d5:	data_out=16'h9ae;
17'hb8d6:	data_out=16'h89fe;
17'hb8d7:	data_out=16'h8a00;
17'hb8d8:	data_out=16'h9c0;
17'hb8d9:	data_out=16'h8a00;
17'hb8da:	data_out=16'h811b;
17'hb8db:	data_out=16'h8a00;
17'hb8dc:	data_out=16'h8a00;
17'hb8dd:	data_out=16'h8a00;
17'hb8de:	data_out=16'h8a00;
17'hb8df:	data_out=16'h8a00;
17'hb8e0:	data_out=16'ha00;
17'hb8e1:	data_out=16'h8a00;
17'hb8e2:	data_out=16'h83e;
17'hb8e3:	data_out=16'h8a00;
17'hb8e4:	data_out=16'h89f0;
17'hb8e5:	data_out=16'h8a00;
17'hb8e6:	data_out=16'h8848;
17'hb8e7:	data_out=16'h8425;
17'hb8e8:	data_out=16'h334;
17'hb8e9:	data_out=16'h9d9;
17'hb8ea:	data_out=16'h180;
17'hb8eb:	data_out=16'h8a00;
17'hb8ec:	data_out=16'h8a00;
17'hb8ed:	data_out=16'h8a00;
17'hb8ee:	data_out=16'h186;
17'hb8ef:	data_out=16'h89ff;
17'hb8f0:	data_out=16'h1f2;
17'hb8f1:	data_out=16'h89f7;
17'hb8f2:	data_out=16'h8a00;
17'hb8f3:	data_out=16'h8a00;
17'hb8f4:	data_out=16'h8580;
17'hb8f5:	data_out=16'h8a00;
17'hb8f6:	data_out=16'h847b;
17'hb8f7:	data_out=16'h9e2;
17'hb8f8:	data_out=16'h89fd;
17'hb8f9:	data_out=16'h83c8;
17'hb8fa:	data_out=16'h8a00;
17'hb8fb:	data_out=16'h33e;
17'hb8fc:	data_out=16'h8a00;
17'hb8fd:	data_out=16'h8a00;
17'hb8fe:	data_out=16'h298;
17'hb8ff:	data_out=16'h8a00;
17'hb900:	data_out=16'h8a00;
17'hb901:	data_out=16'h8a00;
17'hb902:	data_out=16'h856;
17'hb903:	data_out=16'h5da;
17'hb904:	data_out=16'h8a00;
17'hb905:	data_out=16'h8a00;
17'hb906:	data_out=16'h8107;
17'hb907:	data_out=16'ha00;
17'hb908:	data_out=16'h26c;
17'hb909:	data_out=16'h9fd;
17'hb90a:	data_out=16'h8a00;
17'hb90b:	data_out=16'h9ff;
17'hb90c:	data_out=16'ha00;
17'hb90d:	data_out=16'ha00;
17'hb90e:	data_out=16'h2d2;
17'hb90f:	data_out=16'h9c0;
17'hb910:	data_out=16'h8a00;
17'hb911:	data_out=16'h8a00;
17'hb912:	data_out=16'h82e;
17'hb913:	data_out=16'h9f4;
17'hb914:	data_out=16'h84cf;
17'hb915:	data_out=16'h8a00;
17'hb916:	data_out=16'h89fd;
17'hb917:	data_out=16'h9c7;
17'hb918:	data_out=16'h86da;
17'hb919:	data_out=16'hb7;
17'hb91a:	data_out=16'h8a00;
17'hb91b:	data_out=16'h9e7;
17'hb91c:	data_out=16'h8a00;
17'hb91d:	data_out=16'h8a00;
17'hb91e:	data_out=16'h89ff;
17'hb91f:	data_out=16'h8440;
17'hb920:	data_out=16'h8a00;
17'hb921:	data_out=16'h391;
17'hb922:	data_out=16'h3ed;
17'hb923:	data_out=16'ha00;
17'hb924:	data_out=16'ha00;
17'hb925:	data_out=16'h9d1;
17'hb926:	data_out=16'ha00;
17'hb927:	data_out=16'h8a00;
17'hb928:	data_out=16'h3c6;
17'hb929:	data_out=16'h8f6;
17'hb92a:	data_out=16'h597;
17'hb92b:	data_out=16'h86da;
17'hb92c:	data_out=16'h89ff;
17'hb92d:	data_out=16'h9fa;
17'hb92e:	data_out=16'h801b;
17'hb92f:	data_out=16'h8a00;
17'hb930:	data_out=16'h808b;
17'hb931:	data_out=16'h8a00;
17'hb932:	data_out=16'h89fd;
17'hb933:	data_out=16'h8a00;
17'hb934:	data_out=16'h8a00;
17'hb935:	data_out=16'h89fe;
17'hb936:	data_out=16'h89fc;
17'hb937:	data_out=16'h9b1;
17'hb938:	data_out=16'h8a00;
17'hb939:	data_out=16'h8a00;
17'hb93a:	data_out=16'h9d5;
17'hb93b:	data_out=16'h847d;
17'hb93c:	data_out=16'h113;
17'hb93d:	data_out=16'h8a00;
17'hb93e:	data_out=16'h3c7;
17'hb93f:	data_out=16'h8a00;
17'hb940:	data_out=16'h8a00;
17'hb941:	data_out=16'h809c;
17'hb942:	data_out=16'ha00;
17'hb943:	data_out=16'h89ed;
17'hb944:	data_out=16'h8a00;
17'hb945:	data_out=16'h8a00;
17'hb946:	data_out=16'h9f4;
17'hb947:	data_out=16'h9f5;
17'hb948:	data_out=16'h89fe;
17'hb949:	data_out=16'h9e5;
17'hb94a:	data_out=16'h8314;
17'hb94b:	data_out=16'ha00;
17'hb94c:	data_out=16'h9ef;
17'hb94d:	data_out=16'h80ed;
17'hb94e:	data_out=16'h371;
17'hb94f:	data_out=16'h9fe;
17'hb950:	data_out=16'h8a00;
17'hb951:	data_out=16'h9ca;
17'hb952:	data_out=16'ha00;
17'hb953:	data_out=16'h89ff;
17'hb954:	data_out=16'h8a00;
17'hb955:	data_out=16'h9e6;
17'hb956:	data_out=16'h3c7;
17'hb957:	data_out=16'h8a00;
17'hb958:	data_out=16'h9cd;
17'hb959:	data_out=16'h8a00;
17'hb95a:	data_out=16'h335;
17'hb95b:	data_out=16'h8a00;
17'hb95c:	data_out=16'h8a00;
17'hb95d:	data_out=16'h8a00;
17'hb95e:	data_out=16'h8a00;
17'hb95f:	data_out=16'h8a00;
17'hb960:	data_out=16'ha00;
17'hb961:	data_out=16'h8a00;
17'hb962:	data_out=16'h9c0;
17'hb963:	data_out=16'h89ff;
17'hb964:	data_out=16'h8a00;
17'hb965:	data_out=16'h8a00;
17'hb966:	data_out=16'h2e6;
17'hb967:	data_out=16'h803e;
17'hb968:	data_out=16'h3ea;
17'hb969:	data_out=16'h9e0;
17'hb96a:	data_out=16'h233;
17'hb96b:	data_out=16'h8a00;
17'hb96c:	data_out=16'h8a00;
17'hb96d:	data_out=16'h89ff;
17'hb96e:	data_out=16'h239;
17'hb96f:	data_out=16'h89fd;
17'hb970:	data_out=16'h29a;
17'hb971:	data_out=16'h85a1;
17'hb972:	data_out=16'h8a00;
17'hb973:	data_out=16'h8a00;
17'hb974:	data_out=16'hb4;
17'hb975:	data_out=16'h8a00;
17'hb976:	data_out=16'h9f2;
17'hb977:	data_out=16'h9fc;
17'hb978:	data_out=16'h8a00;
17'hb979:	data_out=16'h87;
17'hb97a:	data_out=16'h89f7;
17'hb97b:	data_out=16'h3cf;
17'hb97c:	data_out=16'h8a00;
17'hb97d:	data_out=16'h8a00;
17'hb97e:	data_out=16'h5c0;
17'hb97f:	data_out=16'h8a00;
17'hb980:	data_out=16'h8a00;
17'hb981:	data_out=16'h8a00;
17'hb982:	data_out=16'h9f2;
17'hb983:	data_out=16'h9fb;
17'hb984:	data_out=16'h8a00;
17'hb985:	data_out=16'h8a00;
17'hb986:	data_out=16'h89fd;
17'hb987:	data_out=16'ha00;
17'hb988:	data_out=16'h4f8;
17'hb989:	data_out=16'ha00;
17'hb98a:	data_out=16'h8a00;
17'hb98b:	data_out=16'ha00;
17'hb98c:	data_out=16'ha00;
17'hb98d:	data_out=16'ha00;
17'hb98e:	data_out=16'h9fb;
17'hb98f:	data_out=16'h9fd;
17'hb990:	data_out=16'h8a00;
17'hb991:	data_out=16'h8a00;
17'hb992:	data_out=16'h9f4;
17'hb993:	data_out=16'ha00;
17'hb994:	data_out=16'h636;
17'hb995:	data_out=16'h8a00;
17'hb996:	data_out=16'h8794;
17'hb997:	data_out=16'h9e2;
17'hb998:	data_out=16'h8037;
17'hb999:	data_out=16'h89e4;
17'hb99a:	data_out=16'h8a00;
17'hb99b:	data_out=16'ha00;
17'hb99c:	data_out=16'h89f9;
17'hb99d:	data_out=16'h8a00;
17'hb99e:	data_out=16'h882e;
17'hb99f:	data_out=16'h543;
17'hb9a0:	data_out=16'h8a00;
17'hb9a1:	data_out=16'h9fb;
17'hb9a2:	data_out=16'h892e;
17'hb9a3:	data_out=16'ha00;
17'hb9a4:	data_out=16'ha00;
17'hb9a5:	data_out=16'h9f1;
17'hb9a6:	data_out=16'ha00;
17'hb9a7:	data_out=16'h89fe;
17'hb9a8:	data_out=16'h9fa;
17'hb9a9:	data_out=16'h9a1;
17'hb9aa:	data_out=16'h9da;
17'hb9ab:	data_out=16'h89ab;
17'hb9ac:	data_out=16'h89fb;
17'hb9ad:	data_out=16'h9fd;
17'hb9ae:	data_out=16'h91d;
17'hb9af:	data_out=16'h8a00;
17'hb9b0:	data_out=16'h3ed;
17'hb9b1:	data_out=16'h8a00;
17'hb9b2:	data_out=16'h8a00;
17'hb9b3:	data_out=16'h89ea;
17'hb9b4:	data_out=16'h8a00;
17'hb9b5:	data_out=16'h89f1;
17'hb9b6:	data_out=16'h89f0;
17'hb9b7:	data_out=16'h9f8;
17'hb9b8:	data_out=16'h8a00;
17'hb9b9:	data_out=16'h89f6;
17'hb9ba:	data_out=16'ha00;
17'hb9bb:	data_out=16'h137;
17'hb9bc:	data_out=16'h8386;
17'hb9bd:	data_out=16'h8a00;
17'hb9be:	data_out=16'h9fa;
17'hb9bf:	data_out=16'h8a00;
17'hb9c0:	data_out=16'h8a00;
17'hb9c1:	data_out=16'h2f9;
17'hb9c2:	data_out=16'ha00;
17'hb9c3:	data_out=16'h8a00;
17'hb9c4:	data_out=16'h8a00;
17'hb9c5:	data_out=16'h8a00;
17'hb9c6:	data_out=16'h9d7;
17'hb9c7:	data_out=16'ha00;
17'hb9c8:	data_out=16'h89ef;
17'hb9c9:	data_out=16'h9fa;
17'hb9ca:	data_out=16'h89f1;
17'hb9cb:	data_out=16'ha00;
17'hb9cc:	data_out=16'h9eb;
17'hb9cd:	data_out=16'h8a00;
17'hb9ce:	data_out=16'h9fb;
17'hb9cf:	data_out=16'ha00;
17'hb9d0:	data_out=16'h8a00;
17'hb9d1:	data_out=16'ha00;
17'hb9d2:	data_out=16'ha00;
17'hb9d3:	data_out=16'h89ff;
17'hb9d4:	data_out=16'h8a00;
17'hb9d5:	data_out=16'ha00;
17'hb9d6:	data_out=16'h9f1;
17'hb9d7:	data_out=16'h54b;
17'hb9d8:	data_out=16'h9ec;
17'hb9d9:	data_out=16'h8a00;
17'hb9da:	data_out=16'h7b9;
17'hb9db:	data_out=16'h8a00;
17'hb9dc:	data_out=16'h8a00;
17'hb9dd:	data_out=16'h8a00;
17'hb9de:	data_out=16'h8a00;
17'hb9df:	data_out=16'h8a00;
17'hb9e0:	data_out=16'ha00;
17'hb9e1:	data_out=16'h8a00;
17'hb9e2:	data_out=16'h9dc;
17'hb9e3:	data_out=16'h89ed;
17'hb9e4:	data_out=16'h8a00;
17'hb9e5:	data_out=16'h8a00;
17'hb9e6:	data_out=16'h9d0;
17'hb9e7:	data_out=16'h7df;
17'hb9e8:	data_out=16'h9fb;
17'hb9e9:	data_out=16'ha00;
17'hb9ea:	data_out=16'h9fb;
17'hb9eb:	data_out=16'h8a00;
17'hb9ec:	data_out=16'h8a00;
17'hb9ed:	data_out=16'h89ee;
17'hb9ee:	data_out=16'h9fb;
17'hb9ef:	data_out=16'h8a00;
17'hb9f0:	data_out=16'h9fb;
17'hb9f1:	data_out=16'h9f7;
17'hb9f2:	data_out=16'h8a00;
17'hb9f3:	data_out=16'h8a00;
17'hb9f4:	data_out=16'h5a2;
17'hb9f5:	data_out=16'h8a00;
17'hb9f6:	data_out=16'ha00;
17'hb9f7:	data_out=16'ha00;
17'hb9f8:	data_out=16'h8a00;
17'hb9f9:	data_out=16'h929;
17'hb9fa:	data_out=16'h8941;
17'hb9fb:	data_out=16'h9fa;
17'hb9fc:	data_out=16'h8a00;
17'hb9fd:	data_out=16'h8a00;
17'hb9fe:	data_out=16'h946;
17'hb9ff:	data_out=16'h8a00;
17'hba00:	data_out=16'h8a00;
17'hba01:	data_out=16'h8a00;
17'hba02:	data_out=16'ha00;
17'hba03:	data_out=16'h9fb;
17'hba04:	data_out=16'h89d1;
17'hba05:	data_out=16'h8a00;
17'hba06:	data_out=16'h84de;
17'hba07:	data_out=16'ha00;
17'hba08:	data_out=16'h8557;
17'hba09:	data_out=16'ha00;
17'hba0a:	data_out=16'h8955;
17'hba0b:	data_out=16'h9b9;
17'hba0c:	data_out=16'ha00;
17'hba0d:	data_out=16'ha00;
17'hba0e:	data_out=16'ha00;
17'hba0f:	data_out=16'ha00;
17'hba10:	data_out=16'h89f6;
17'hba11:	data_out=16'h8a00;
17'hba12:	data_out=16'h188;
17'hba13:	data_out=16'h9ee;
17'hba14:	data_out=16'h95b;
17'hba15:	data_out=16'h89fc;
17'hba16:	data_out=16'h8629;
17'hba17:	data_out=16'h9c4;
17'hba18:	data_out=16'h31a;
17'hba19:	data_out=16'h89d6;
17'hba1a:	data_out=16'h8a00;
17'hba1b:	data_out=16'ha00;
17'hba1c:	data_out=16'h89e9;
17'hba1d:	data_out=16'h8a00;
17'hba1e:	data_out=16'h83cd;
17'hba1f:	data_out=16'h8d7;
17'hba20:	data_out=16'h8a00;
17'hba21:	data_out=16'ha00;
17'hba22:	data_out=16'h89fe;
17'hba23:	data_out=16'ha00;
17'hba24:	data_out=16'ha00;
17'hba25:	data_out=16'ha00;
17'hba26:	data_out=16'ha00;
17'hba27:	data_out=16'h89f9;
17'hba28:	data_out=16'ha00;
17'hba29:	data_out=16'h9b8;
17'hba2a:	data_out=16'h9ff;
17'hba2b:	data_out=16'h89f6;
17'hba2c:	data_out=16'h89c0;
17'hba2d:	data_out=16'h89e2;
17'hba2e:	data_out=16'h8724;
17'hba2f:	data_out=16'h89fe;
17'hba30:	data_out=16'ha00;
17'hba31:	data_out=16'h8a00;
17'hba32:	data_out=16'h89e5;
17'hba33:	data_out=16'h89e7;
17'hba34:	data_out=16'h8a00;
17'hba35:	data_out=16'h8793;
17'hba36:	data_out=16'h89d5;
17'hba37:	data_out=16'ha00;
17'hba38:	data_out=16'h8a00;
17'hba39:	data_out=16'h89f1;
17'hba3a:	data_out=16'ha00;
17'hba3b:	data_out=16'h9ab;
17'hba3c:	data_out=16'h88d5;
17'hba3d:	data_out=16'h8a00;
17'hba3e:	data_out=16'ha00;
17'hba3f:	data_out=16'h8a00;
17'hba40:	data_out=16'h89e4;
17'hba41:	data_out=16'h8179;
17'hba42:	data_out=16'ha00;
17'hba43:	data_out=16'h8a00;
17'hba44:	data_out=16'h89f9;
17'hba45:	data_out=16'h89fb;
17'hba46:	data_out=16'h85bd;
17'hba47:	data_out=16'h9ff;
17'hba48:	data_out=16'h89db;
17'hba49:	data_out=16'ha00;
17'hba4a:	data_out=16'h89ce;
17'hba4b:	data_out=16'h9f3;
17'hba4c:	data_out=16'h9f5;
17'hba4d:	data_out=16'h89ff;
17'hba4e:	data_out=16'h82a9;
17'hba4f:	data_out=16'ha00;
17'hba50:	data_out=16'h89fb;
17'hba51:	data_out=16'ha00;
17'hba52:	data_out=16'ha00;
17'hba53:	data_out=16'h89f6;
17'hba54:	data_out=16'h8a00;
17'hba55:	data_out=16'ha00;
17'hba56:	data_out=16'ha00;
17'hba57:	data_out=16'h9c5;
17'hba58:	data_out=16'h9d9;
17'hba59:	data_out=16'h89ea;
17'hba5a:	data_out=16'h7a4;
17'hba5b:	data_out=16'h89f9;
17'hba5c:	data_out=16'h89ff;
17'hba5d:	data_out=16'h89ff;
17'hba5e:	data_out=16'h89fb;
17'hba5f:	data_out=16'h89ff;
17'hba60:	data_out=16'ha00;
17'hba61:	data_out=16'h89fd;
17'hba62:	data_out=16'h9bc;
17'hba63:	data_out=16'h89eb;
17'hba64:	data_out=16'h8a00;
17'hba65:	data_out=16'h8a00;
17'hba66:	data_out=16'h9fd;
17'hba67:	data_out=16'h9ff;
17'hba68:	data_out=16'ha00;
17'hba69:	data_out=16'h9f0;
17'hba6a:	data_out=16'ha00;
17'hba6b:	data_out=16'h8a00;
17'hba6c:	data_out=16'h8a00;
17'hba6d:	data_out=16'h89eb;
17'hba6e:	data_out=16'ha00;
17'hba6f:	data_out=16'h89fa;
17'hba70:	data_out=16'ha00;
17'hba71:	data_out=16'h9ff;
17'hba72:	data_out=16'h8a00;
17'hba73:	data_out=16'h8a00;
17'hba74:	data_out=16'ha00;
17'hba75:	data_out=16'h8a00;
17'hba76:	data_out=16'h9f9;
17'hba77:	data_out=16'ha00;
17'hba78:	data_out=16'h8a00;
17'hba79:	data_out=16'h1ee;
17'hba7a:	data_out=16'h86fc;
17'hba7b:	data_out=16'ha00;
17'hba7c:	data_out=16'h89fc;
17'hba7d:	data_out=16'h89fa;
17'hba7e:	data_out=16'h9cc;
17'hba7f:	data_out=16'h8a00;
17'hba80:	data_out=16'h89ff;
17'hba81:	data_out=16'h8a00;
17'hba82:	data_out=16'ha00;
17'hba83:	data_out=16'h7f5;
17'hba84:	data_out=16'h8925;
17'hba85:	data_out=16'h8998;
17'hba86:	data_out=16'h839c;
17'hba87:	data_out=16'ha00;
17'hba88:	data_out=16'h82fc;
17'hba89:	data_out=16'ha00;
17'hba8a:	data_out=16'h8863;
17'hba8b:	data_out=16'h623;
17'hba8c:	data_out=16'ha00;
17'hba8d:	data_out=16'ha00;
17'hba8e:	data_out=16'ha00;
17'hba8f:	data_out=16'ha00;
17'hba90:	data_out=16'h89f6;
17'hba91:	data_out=16'h8a00;
17'hba92:	data_out=16'h835d;
17'hba93:	data_out=16'h5e7;
17'hba94:	data_out=16'h738;
17'hba95:	data_out=16'h89b8;
17'hba96:	data_out=16'h8393;
17'hba97:	data_out=16'h6df;
17'hba98:	data_out=16'h9fc;
17'hba99:	data_out=16'h8a00;
17'hba9a:	data_out=16'h89e9;
17'hba9b:	data_out=16'ha00;
17'hba9c:	data_out=16'h89be;
17'hba9d:	data_out=16'h8a00;
17'hba9e:	data_out=16'h803a;
17'hba9f:	data_out=16'h9cf;
17'hbaa0:	data_out=16'h8a00;
17'hbaa1:	data_out=16'ha00;
17'hbaa2:	data_out=16'h89fc;
17'hbaa3:	data_out=16'ha00;
17'hbaa4:	data_out=16'ha00;
17'hbaa5:	data_out=16'ha00;
17'hbaa6:	data_out=16'ha00;
17'hbaa7:	data_out=16'h89e3;
17'hbaa8:	data_out=16'ha00;
17'hbaa9:	data_out=16'h9a2;
17'hbaaa:	data_out=16'h9fe;
17'hbaab:	data_out=16'h8a00;
17'hbaac:	data_out=16'h87cd;
17'hbaad:	data_out=16'h8a00;
17'hbaae:	data_out=16'h8181;
17'hbaaf:	data_out=16'h89fb;
17'hbab0:	data_out=16'ha00;
17'hbab1:	data_out=16'h89c9;
17'hbab2:	data_out=16'h8929;
17'hbab3:	data_out=16'h89e5;
17'hbab4:	data_out=16'h8a00;
17'hbab5:	data_out=16'hf6;
17'hbab6:	data_out=16'h8986;
17'hbab7:	data_out=16'ha00;
17'hbab8:	data_out=16'h8a00;
17'hbab9:	data_out=16'h89ed;
17'hbaba:	data_out=16'h9f7;
17'hbabb:	data_out=16'ha00;
17'hbabc:	data_out=16'h8967;
17'hbabd:	data_out=16'h89cb;
17'hbabe:	data_out=16'ha00;
17'hbabf:	data_out=16'h8996;
17'hbac0:	data_out=16'h895b;
17'hbac1:	data_out=16'ha00;
17'hbac2:	data_out=16'ha00;
17'hbac3:	data_out=16'h8857;
17'hbac4:	data_out=16'h897b;
17'hbac5:	data_out=16'h89a9;
17'hbac6:	data_out=16'h89ec;
17'hbac7:	data_out=16'h9cd;
17'hbac8:	data_out=16'h89d4;
17'hbac9:	data_out=16'ha00;
17'hbaca:	data_out=16'h89c8;
17'hbacb:	data_out=16'h9d1;
17'hbacc:	data_out=16'h9fc;
17'hbacd:	data_out=16'h8a00;
17'hbace:	data_out=16'h631;
17'hbacf:	data_out=16'h9fd;
17'hbad0:	data_out=16'h89e7;
17'hbad1:	data_out=16'ha00;
17'hbad2:	data_out=16'ha00;
17'hbad3:	data_out=16'h89f3;
17'hbad4:	data_out=16'h8a00;
17'hbad5:	data_out=16'ha00;
17'hbad6:	data_out=16'ha00;
17'hbad7:	data_out=16'h9fd;
17'hbad8:	data_out=16'ha00;
17'hbad9:	data_out=16'h8980;
17'hbada:	data_out=16'h4cc;
17'hbadb:	data_out=16'h8980;
17'hbadc:	data_out=16'h89db;
17'hbadd:	data_out=16'h89ae;
17'hbade:	data_out=16'h89b0;
17'hbadf:	data_out=16'h8a00;
17'hbae0:	data_out=16'ha00;
17'hbae1:	data_out=16'h8921;
17'hbae2:	data_out=16'h9d9;
17'hbae3:	data_out=16'h89ea;
17'hbae4:	data_out=16'h8a00;
17'hbae5:	data_out=16'h8a00;
17'hbae6:	data_out=16'h9e4;
17'hbae7:	data_out=16'h9d6;
17'hbae8:	data_out=16'ha00;
17'hbae9:	data_out=16'h9e8;
17'hbaea:	data_out=16'ha00;
17'hbaeb:	data_out=16'h89c4;
17'hbaec:	data_out=16'h89dc;
17'hbaed:	data_out=16'h89ea;
17'hbaee:	data_out=16'ha00;
17'hbaef:	data_out=16'h8993;
17'hbaf0:	data_out=16'ha00;
17'hbaf1:	data_out=16'h9fe;
17'hbaf2:	data_out=16'h89dd;
17'hbaf3:	data_out=16'h89b2;
17'hbaf4:	data_out=16'ha00;
17'hbaf5:	data_out=16'h89a4;
17'hbaf6:	data_out=16'h9de;
17'hbaf7:	data_out=16'ha00;
17'hbaf8:	data_out=16'h8a00;
17'hbaf9:	data_out=16'h9ef;
17'hbafa:	data_out=16'h85db;
17'hbafb:	data_out=16'ha00;
17'hbafc:	data_out=16'h89f2;
17'hbafd:	data_out=16'h488;
17'hbafe:	data_out=16'h9dc;
17'hbaff:	data_out=16'h8a00;
17'hbb00:	data_out=16'h8a00;
17'hbb01:	data_out=16'h8a00;
17'hbb02:	data_out=16'ha00;
17'hbb03:	data_out=16'h8541;
17'hbb04:	data_out=16'h8951;
17'hbb05:	data_out=16'h89a2;
17'hbb06:	data_out=16'h1f7;
17'hbb07:	data_out=16'ha00;
17'hbb08:	data_out=16'h9c7;
17'hbb09:	data_out=16'ha00;
17'hbb0a:	data_out=16'h8952;
17'hbb0b:	data_out=16'h89a2;
17'hbb0c:	data_out=16'ha00;
17'hbb0d:	data_out=16'ha00;
17'hbb0e:	data_out=16'ha00;
17'hbb0f:	data_out=16'ha00;
17'hbb10:	data_out=16'h89f6;
17'hbb11:	data_out=16'h8a00;
17'hbb12:	data_out=16'h8a4;
17'hbb13:	data_out=16'h8863;
17'hbb14:	data_out=16'h83c5;
17'hbb15:	data_out=16'h8906;
17'hbb16:	data_out=16'h860e;
17'hbb17:	data_out=16'h880e;
17'hbb18:	data_out=16'h9fe;
17'hbb19:	data_out=16'h8a00;
17'hbb1a:	data_out=16'h8a00;
17'hbb1b:	data_out=16'ha00;
17'hbb1c:	data_out=16'h89ca;
17'hbb1d:	data_out=16'h8a00;
17'hbb1e:	data_out=16'h8241;
17'hbb1f:	data_out=16'h989;
17'hbb20:	data_out=16'h8a00;
17'hbb21:	data_out=16'ha00;
17'hbb22:	data_out=16'h874c;
17'hbb23:	data_out=16'ha00;
17'hbb24:	data_out=16'ha00;
17'hbb25:	data_out=16'ha00;
17'hbb26:	data_out=16'ha00;
17'hbb27:	data_out=16'h8a00;
17'hbb28:	data_out=16'ha00;
17'hbb29:	data_out=16'h82db;
17'hbb2a:	data_out=16'h9ff;
17'hbb2b:	data_out=16'h8a00;
17'hbb2c:	data_out=16'h879b;
17'hbb2d:	data_out=16'h8a00;
17'hbb2e:	data_out=16'h9b9;
17'hbb2f:	data_out=16'h8a00;
17'hbb30:	data_out=16'h9ff;
17'hbb31:	data_out=16'h8a00;
17'hbb32:	data_out=16'h8760;
17'hbb33:	data_out=16'h89fb;
17'hbb34:	data_out=16'h8a00;
17'hbb35:	data_out=16'h9fb;
17'hbb36:	data_out=16'h84c8;
17'hbb37:	data_out=16'ha00;
17'hbb38:	data_out=16'h8a00;
17'hbb39:	data_out=16'h89fb;
17'hbb3a:	data_out=16'ha00;
17'hbb3b:	data_out=16'ha00;
17'hbb3c:	data_out=16'h8990;
17'hbb3d:	data_out=16'h89ef;
17'hbb3e:	data_out=16'ha00;
17'hbb3f:	data_out=16'h899f;
17'hbb40:	data_out=16'h896a;
17'hbb41:	data_out=16'ha00;
17'hbb42:	data_out=16'ha00;
17'hbb43:	data_out=16'h8a00;
17'hbb44:	data_out=16'h89db;
17'hbb45:	data_out=16'h88f8;
17'hbb46:	data_out=16'h8a00;
17'hbb47:	data_out=16'h9a0;
17'hbb48:	data_out=16'h844e;
17'hbb49:	data_out=16'ha00;
17'hbb4a:	data_out=16'h86b9;
17'hbb4b:	data_out=16'h852;
17'hbb4c:	data_out=16'ha00;
17'hbb4d:	data_out=16'h8a00;
17'hbb4e:	data_out=16'h478;
17'hbb4f:	data_out=16'ha00;
17'hbb50:	data_out=16'h89e8;
17'hbb51:	data_out=16'ha00;
17'hbb52:	data_out=16'ha00;
17'hbb53:	data_out=16'h89ff;
17'hbb54:	data_out=16'h8a00;
17'hbb55:	data_out=16'ha00;
17'hbb56:	data_out=16'ha00;
17'hbb57:	data_out=16'h9ff;
17'hbb58:	data_out=16'ha00;
17'hbb59:	data_out=16'h8999;
17'hbb5a:	data_out=16'h7b2;
17'hbb5b:	data_out=16'h8a00;
17'hbb5c:	data_out=16'h89a2;
17'hbb5d:	data_out=16'h8989;
17'hbb5e:	data_out=16'h88dd;
17'hbb5f:	data_out=16'h8a00;
17'hbb60:	data_out=16'ha00;
17'hbb61:	data_out=16'h8944;
17'hbb62:	data_out=16'h8732;
17'hbb63:	data_out=16'h89fb;
17'hbb64:	data_out=16'h8a00;
17'hbb65:	data_out=16'h8a00;
17'hbb66:	data_out=16'h92f;
17'hbb67:	data_out=16'h8d6;
17'hbb68:	data_out=16'ha00;
17'hbb69:	data_out=16'ha00;
17'hbb6a:	data_out=16'ha00;
17'hbb6b:	data_out=16'h89f7;
17'hbb6c:	data_out=16'h89ee;
17'hbb6d:	data_out=16'h89fc;
17'hbb6e:	data_out=16'ha00;
17'hbb6f:	data_out=16'h89c5;
17'hbb70:	data_out=16'ha00;
17'hbb71:	data_out=16'ha00;
17'hbb72:	data_out=16'h89f8;
17'hbb73:	data_out=16'h89fa;
17'hbb74:	data_out=16'ha00;
17'hbb75:	data_out=16'h8814;
17'hbb76:	data_out=16'h7ec;
17'hbb77:	data_out=16'ha00;
17'hbb78:	data_out=16'h8a00;
17'hbb79:	data_out=16'ha00;
17'hbb7a:	data_out=16'h88a2;
17'hbb7b:	data_out=16'ha00;
17'hbb7c:	data_out=16'h66;
17'hbb7d:	data_out=16'h951;
17'hbb7e:	data_out=16'h9f5;
17'hbb7f:	data_out=16'h8a00;
17'hbb80:	data_out=16'h8a00;
17'hbb81:	data_out=16'h8a00;
17'hbb82:	data_out=16'ha00;
17'hbb83:	data_out=16'h89b1;
17'hbb84:	data_out=16'h87ba;
17'hbb85:	data_out=16'h87f4;
17'hbb86:	data_out=16'h4af;
17'hbb87:	data_out=16'ha00;
17'hbb88:	data_out=16'h9a8;
17'hbb89:	data_out=16'ha00;
17'hbb8a:	data_out=16'h8988;
17'hbb8b:	data_out=16'h8a00;
17'hbb8c:	data_out=16'h9ad;
17'hbb8d:	data_out=16'ha00;
17'hbb8e:	data_out=16'ha00;
17'hbb8f:	data_out=16'ha00;
17'hbb90:	data_out=16'h8a00;
17'hbb91:	data_out=16'h89ff;
17'hbb92:	data_out=16'h8714;
17'hbb93:	data_out=16'h86c5;
17'hbb94:	data_out=16'h89e6;
17'hbb95:	data_out=16'h88c8;
17'hbb96:	data_out=16'h87ec;
17'hbb97:	data_out=16'h89f0;
17'hbb98:	data_out=16'ha00;
17'hbb99:	data_out=16'h8a00;
17'hbb9a:	data_out=16'h89f9;
17'hbb9b:	data_out=16'h8629;
17'hbb9c:	data_out=16'h89c9;
17'hbb9d:	data_out=16'h8a00;
17'hbb9e:	data_out=16'h8957;
17'hbb9f:	data_out=16'h9a0;
17'hbba0:	data_out=16'h8a00;
17'hbba1:	data_out=16'ha00;
17'hbba2:	data_out=16'h89a8;
17'hbba3:	data_out=16'ha00;
17'hbba4:	data_out=16'ha00;
17'hbba5:	data_out=16'ha00;
17'hbba6:	data_out=16'ha00;
17'hbba7:	data_out=16'h8a00;
17'hbba8:	data_out=16'ha00;
17'hbba9:	data_out=16'h8a00;
17'hbbaa:	data_out=16'h925;
17'hbbab:	data_out=16'h8a00;
17'hbbac:	data_out=16'h8904;
17'hbbad:	data_out=16'h8a00;
17'hbbae:	data_out=16'h1e;
17'hbbaf:	data_out=16'h8a00;
17'hbbb0:	data_out=16'h9fd;
17'hbbb1:	data_out=16'h8a00;
17'hbbb2:	data_out=16'h4d4;
17'hbbb3:	data_out=16'h89ff;
17'hbbb4:	data_out=16'h8a00;
17'hbbb5:	data_out=16'h8343;
17'hbbb6:	data_out=16'h865d;
17'hbbb7:	data_out=16'ha00;
17'hbbb8:	data_out=16'h8a00;
17'hbbb9:	data_out=16'h8a00;
17'hbbba:	data_out=16'h569;
17'hbbbb:	data_out=16'ha00;
17'hbbbc:	data_out=16'h8a00;
17'hbbbd:	data_out=16'h89fe;
17'hbbbe:	data_out=16'ha00;
17'hbbbf:	data_out=16'h87c6;
17'hbbc0:	data_out=16'h872e;
17'hbbc1:	data_out=16'h10b;
17'hbbc2:	data_out=16'h87cb;
17'hbbc3:	data_out=16'h8a00;
17'hbbc4:	data_out=16'h89e8;
17'hbbc5:	data_out=16'h88ca;
17'hbbc6:	data_out=16'h8a00;
17'hbbc7:	data_out=16'h719;
17'hbbc8:	data_out=16'h84f4;
17'hbbc9:	data_out=16'h9ff;
17'hbbca:	data_out=16'h341;
17'hbbcb:	data_out=16'h89f2;
17'hbbcc:	data_out=16'ha00;
17'hbbcd:	data_out=16'h8a00;
17'hbbce:	data_out=16'h87a7;
17'hbbcf:	data_out=16'h9ff;
17'hbbd0:	data_out=16'h8a00;
17'hbbd1:	data_out=16'ha00;
17'hbbd2:	data_out=16'ha00;
17'hbbd3:	data_out=16'h8a00;
17'hbbd4:	data_out=16'h8a00;
17'hbbd5:	data_out=16'ha00;
17'hbbd6:	data_out=16'ha00;
17'hbbd7:	data_out=16'ha00;
17'hbbd8:	data_out=16'ha00;
17'hbbd9:	data_out=16'h89a6;
17'hbbda:	data_out=16'h815b;
17'hbbdb:	data_out=16'h8a00;
17'hbbdc:	data_out=16'h889e;
17'hbbdd:	data_out=16'h887d;
17'hbbde:	data_out=16'h8847;
17'hbbdf:	data_out=16'h8a00;
17'hbbe0:	data_out=16'ha00;
17'hbbe1:	data_out=16'h88a8;
17'hbbe2:	data_out=16'h89b5;
17'hbbe3:	data_out=16'h89ff;
17'hbbe4:	data_out=16'h8a00;
17'hbbe5:	data_out=16'h8a00;
17'hbbe6:	data_out=16'h89ff;
17'hbbe7:	data_out=16'h8a00;
17'hbbe8:	data_out=16'ha00;
17'hbbe9:	data_out=16'h9ee;
17'hbbea:	data_out=16'ha00;
17'hbbeb:	data_out=16'h89f3;
17'hbbec:	data_out=16'h89fd;
17'hbbed:	data_out=16'h89ff;
17'hbbee:	data_out=16'ha00;
17'hbbef:	data_out=16'h89de;
17'hbbf0:	data_out=16'ha00;
17'hbbf1:	data_out=16'ha00;
17'hbbf2:	data_out=16'h89d1;
17'hbbf3:	data_out=16'h89e2;
17'hbbf4:	data_out=16'h9fe;
17'hbbf5:	data_out=16'ha00;
17'hbbf6:	data_out=16'h8a00;
17'hbbf7:	data_out=16'h8244;
17'hbbf8:	data_out=16'h8a00;
17'hbbf9:	data_out=16'ha00;
17'hbbfa:	data_out=16'h89fb;
17'hbbfb:	data_out=16'ha00;
17'hbbfc:	data_out=16'h9f3;
17'hbbfd:	data_out=16'h999;
17'hbbfe:	data_out=16'h831b;
17'hbbff:	data_out=16'h8a00;
17'hbc00:	data_out=16'h8a00;
17'hbc01:	data_out=16'h8a00;
17'hbc02:	data_out=16'ha00;
17'hbc03:	data_out=16'h8a00;
17'hbc04:	data_out=16'h519;
17'hbc05:	data_out=16'ha00;
17'hbc06:	data_out=16'h8019;
17'hbc07:	data_out=16'ha00;
17'hbc08:	data_out=16'h89f2;
17'hbc09:	data_out=16'h89ad;
17'hbc0a:	data_out=16'h803b;
17'hbc0b:	data_out=16'h8a00;
17'hbc0c:	data_out=16'h180;
17'hbc0d:	data_out=16'h84c5;
17'hbc0e:	data_out=16'ha00;
17'hbc0f:	data_out=16'h8936;
17'hbc10:	data_out=16'h8a00;
17'hbc11:	data_out=16'h89f0;
17'hbc12:	data_out=16'h8a00;
17'hbc13:	data_out=16'h85f5;
17'hbc14:	data_out=16'h89ff;
17'hbc15:	data_out=16'h89a5;
17'hbc16:	data_out=16'h89bd;
17'hbc17:	data_out=16'h89ff;
17'hbc18:	data_out=16'h8867;
17'hbc19:	data_out=16'h8a00;
17'hbc1a:	data_out=16'h9ff;
17'hbc1b:	data_out=16'h89d3;
17'hbc1c:	data_out=16'h89c6;
17'hbc1d:	data_out=16'h8a00;
17'hbc1e:	data_out=16'h89fe;
17'hbc1f:	data_out=16'h588;
17'hbc20:	data_out=16'h8a00;
17'hbc21:	data_out=16'ha00;
17'hbc22:	data_out=16'h89e3;
17'hbc23:	data_out=16'ha00;
17'hbc24:	data_out=16'ha00;
17'hbc25:	data_out=16'ha00;
17'hbc26:	data_out=16'h80ce;
17'hbc27:	data_out=16'h8a00;
17'hbc28:	data_out=16'ha00;
17'hbc29:	data_out=16'h8a00;
17'hbc2a:	data_out=16'h89eb;
17'hbc2b:	data_out=16'h8a00;
17'hbc2c:	data_out=16'h89cf;
17'hbc2d:	data_out=16'h8a00;
17'hbc2e:	data_out=16'h89fe;
17'hbc2f:	data_out=16'h8a00;
17'hbc30:	data_out=16'ha00;
17'hbc31:	data_out=16'h86cf;
17'hbc32:	data_out=16'ha00;
17'hbc33:	data_out=16'h8a00;
17'hbc34:	data_out=16'h8a00;
17'hbc35:	data_out=16'h89ed;
17'hbc36:	data_out=16'h89f3;
17'hbc37:	data_out=16'h9f8;
17'hbc38:	data_out=16'h81a5;
17'hbc39:	data_out=16'h8a00;
17'hbc3a:	data_out=16'h8a00;
17'hbc3b:	data_out=16'ha00;
17'hbc3c:	data_out=16'h89d0;
17'hbc3d:	data_out=16'h8a00;
17'hbc3e:	data_out=16'ha00;
17'hbc3f:	data_out=16'ha00;
17'hbc40:	data_out=16'h83d7;
17'hbc41:	data_out=16'h8656;
17'hbc42:	data_out=16'h89d1;
17'hbc43:	data_out=16'h8a00;
17'hbc44:	data_out=16'h893f;
17'hbc45:	data_out=16'h89bb;
17'hbc46:	data_out=16'h89f9;
17'hbc47:	data_out=16'h8a00;
17'hbc48:	data_out=16'h89fc;
17'hbc49:	data_out=16'h52f;
17'hbc4a:	data_out=16'h89fe;
17'hbc4b:	data_out=16'h8a00;
17'hbc4c:	data_out=16'h404;
17'hbc4d:	data_out=16'h8a00;
17'hbc4e:	data_out=16'h89da;
17'hbc4f:	data_out=16'h89c8;
17'hbc50:	data_out=16'h8a00;
17'hbc51:	data_out=16'ha00;
17'hbc52:	data_out=16'ha00;
17'hbc53:	data_out=16'h8a00;
17'hbc54:	data_out=16'h8a00;
17'hbc55:	data_out=16'h837;
17'hbc56:	data_out=16'h9fe;
17'hbc57:	data_out=16'h9f2;
17'hbc58:	data_out=16'h9f9;
17'hbc59:	data_out=16'h88ab;
17'hbc5a:	data_out=16'h604;
17'hbc5b:	data_out=16'h84d1;
17'hbc5c:	data_out=16'h34d;
17'hbc5d:	data_out=16'h89c6;
17'hbc5e:	data_out=16'h88f0;
17'hbc5f:	data_out=16'h8a00;
17'hbc60:	data_out=16'h899f;
17'hbc61:	data_out=16'ha00;
17'hbc62:	data_out=16'h8a00;
17'hbc63:	data_out=16'h89ff;
17'hbc64:	data_out=16'h8a00;
17'hbc65:	data_out=16'h89f9;
17'hbc66:	data_out=16'h89ed;
17'hbc67:	data_out=16'h8a00;
17'hbc68:	data_out=16'ha00;
17'hbc69:	data_out=16'h89f9;
17'hbc6a:	data_out=16'ha00;
17'hbc6b:	data_out=16'h89c2;
17'hbc6c:	data_out=16'h89ff;
17'hbc6d:	data_out=16'h89ff;
17'hbc6e:	data_out=16'ha00;
17'hbc6f:	data_out=16'h80bd;
17'hbc70:	data_out=16'ha00;
17'hbc71:	data_out=16'h88c4;
17'hbc72:	data_out=16'h885e;
17'hbc73:	data_out=16'h9f3;
17'hbc74:	data_out=16'ha00;
17'hbc75:	data_out=16'ha00;
17'hbc76:	data_out=16'h8a00;
17'hbc77:	data_out=16'h89f1;
17'hbc78:	data_out=16'h8a00;
17'hbc79:	data_out=16'h818e;
17'hbc7a:	data_out=16'h89ff;
17'hbc7b:	data_out=16'ha00;
17'hbc7c:	data_out=16'h895e;
17'hbc7d:	data_out=16'h8fa;
17'hbc7e:	data_out=16'h89ab;
17'hbc7f:	data_out=16'h89c1;
17'hbc80:	data_out=16'h8a00;
17'hbc81:	data_out=16'h89f8;
17'hbc82:	data_out=16'h9ae;
17'hbc83:	data_out=16'h8a00;
17'hbc84:	data_out=16'h1b2;
17'hbc85:	data_out=16'ha00;
17'hbc86:	data_out=16'h9ee;
17'hbc87:	data_out=16'h85ed;
17'hbc88:	data_out=16'h89ff;
17'hbc89:	data_out=16'h8a00;
17'hbc8a:	data_out=16'h8942;
17'hbc8b:	data_out=16'h8a00;
17'hbc8c:	data_out=16'h8a00;
17'hbc8d:	data_out=16'h88e3;
17'hbc8e:	data_out=16'ha00;
17'hbc8f:	data_out=16'h89f8;
17'hbc90:	data_out=16'h8a00;
17'hbc91:	data_out=16'h89d5;
17'hbc92:	data_out=16'h8a00;
17'hbc93:	data_out=16'h178;
17'hbc94:	data_out=16'h89ee;
17'hbc95:	data_out=16'h8958;
17'hbc96:	data_out=16'h89ce;
17'hbc97:	data_out=16'h89dc;
17'hbc98:	data_out=16'h89fe;
17'hbc99:	data_out=16'h8a00;
17'hbc9a:	data_out=16'ha00;
17'hbc9b:	data_out=16'h82b7;
17'hbc9c:	data_out=16'h9e9;
17'hbc9d:	data_out=16'h8a00;
17'hbc9e:	data_out=16'h89fa;
17'hbc9f:	data_out=16'h964;
17'hbca0:	data_out=16'h89f6;
17'hbca1:	data_out=16'ha00;
17'hbca2:	data_out=16'h89d3;
17'hbca3:	data_out=16'h88f1;
17'hbca4:	data_out=16'h88ff;
17'hbca5:	data_out=16'h8881;
17'hbca6:	data_out=16'h8a00;
17'hbca7:	data_out=16'h8a00;
17'hbca8:	data_out=16'ha00;
17'hbca9:	data_out=16'h8a00;
17'hbcaa:	data_out=16'h89fc;
17'hbcab:	data_out=16'h8a00;
17'hbcac:	data_out=16'h89d2;
17'hbcad:	data_out=16'h8a00;
17'hbcae:	data_out=16'h89fa;
17'hbcaf:	data_out=16'h89fb;
17'hbcb0:	data_out=16'ha00;
17'hbcb1:	data_out=16'h519;
17'hbcb2:	data_out=16'ha00;
17'hbcb3:	data_out=16'h89fe;
17'hbcb4:	data_out=16'h8a00;
17'hbcb5:	data_out=16'h89fe;
17'hbcb6:	data_out=16'h89fa;
17'hbcb7:	data_out=16'h917;
17'hbcb8:	data_out=16'ha00;
17'hbcb9:	data_out=16'h8a00;
17'hbcba:	data_out=16'h8a00;
17'hbcbb:	data_out=16'h9fd;
17'hbcbc:	data_out=16'h9d7;
17'hbcbd:	data_out=16'h89f6;
17'hbcbe:	data_out=16'ha00;
17'hbcbf:	data_out=16'ha00;
17'hbcc0:	data_out=16'h9fa;
17'hbcc1:	data_out=16'h87d5;
17'hbcc2:	data_out=16'h8a00;
17'hbcc3:	data_out=16'hd5;
17'hbcc4:	data_out=16'h2ad;
17'hbcc5:	data_out=16'h895d;
17'hbcc6:	data_out=16'h89fc;
17'hbcc7:	data_out=16'h8a00;
17'hbcc8:	data_out=16'h89fb;
17'hbcc9:	data_out=16'h896c;
17'hbcca:	data_out=16'h8a00;
17'hbccb:	data_out=16'h8a00;
17'hbccc:	data_out=16'h893d;
17'hbccd:	data_out=16'h89fb;
17'hbcce:	data_out=16'h8a00;
17'hbccf:	data_out=16'h8a00;
17'hbcd0:	data_out=16'h89ff;
17'hbcd1:	data_out=16'ha00;
17'hbcd2:	data_out=16'h899f;
17'hbcd3:	data_out=16'h89f3;
17'hbcd4:	data_out=16'h89ff;
17'hbcd5:	data_out=16'h81b;
17'hbcd6:	data_out=16'h8184;
17'hbcd7:	data_out=16'h79a;
17'hbcd8:	data_out=16'ha00;
17'hbcd9:	data_out=16'h8107;
17'hbcda:	data_out=16'h9e0;
17'hbcdb:	data_out=16'h6e6;
17'hbcdc:	data_out=16'ha00;
17'hbcdd:	data_out=16'h89f2;
17'hbcde:	data_out=16'h88ba;
17'hbcdf:	data_out=16'h8a00;
17'hbce0:	data_out=16'h8a00;
17'hbce1:	data_out=16'ha00;
17'hbce2:	data_out=16'h89f7;
17'hbce3:	data_out=16'h89fa;
17'hbce4:	data_out=16'h8a00;
17'hbce5:	data_out=16'h89f3;
17'hbce6:	data_out=16'h89e9;
17'hbce7:	data_out=16'h8a00;
17'hbce8:	data_out=16'ha00;
17'hbce9:	data_out=16'h8a00;
17'hbcea:	data_out=16'ha00;
17'hbceb:	data_out=16'h9ff;
17'hbcec:	data_out=16'h8a00;
17'hbced:	data_out=16'h89fb;
17'hbcee:	data_out=16'ha00;
17'hbcef:	data_out=16'ha00;
17'hbcf0:	data_out=16'ha00;
17'hbcf1:	data_out=16'h89f6;
17'hbcf2:	data_out=16'h9fe;
17'hbcf3:	data_out=16'ha00;
17'hbcf4:	data_out=16'ha00;
17'hbcf5:	data_out=16'ha00;
17'hbcf6:	data_out=16'h8a00;
17'hbcf7:	data_out=16'h89ff;
17'hbcf8:	data_out=16'h9fd;
17'hbcf9:	data_out=16'h89ab;
17'hbcfa:	data_out=16'h89f7;
17'hbcfb:	data_out=16'ha00;
17'hbcfc:	data_out=16'h89ff;
17'hbcfd:	data_out=16'h9e5;
17'hbcfe:	data_out=16'h84a8;
17'hbcff:	data_out=16'ha00;
17'hbd00:	data_out=16'h89fe;
17'hbd01:	data_out=16'h89fc;
17'hbd02:	data_out=16'h86dc;
17'hbd03:	data_out=16'h291;
17'hbd04:	data_out=16'h8a00;
17'hbd05:	data_out=16'ha00;
17'hbd06:	data_out=16'ha00;
17'hbd07:	data_out=16'h8a00;
17'hbd08:	data_out=16'h8a00;
17'hbd09:	data_out=16'h8a00;
17'hbd0a:	data_out=16'h8a00;
17'hbd0b:	data_out=16'h8a00;
17'hbd0c:	data_out=16'h8a00;
17'hbd0d:	data_out=16'h9b2;
17'hbd0e:	data_out=16'ha00;
17'hbd0f:	data_out=16'h8a00;
17'hbd10:	data_out=16'h8a00;
17'hbd11:	data_out=16'h8a00;
17'hbd12:	data_out=16'h8a00;
17'hbd13:	data_out=16'ha00;
17'hbd14:	data_out=16'h9f2;
17'hbd15:	data_out=16'h89d1;
17'hbd16:	data_out=16'h8998;
17'hbd17:	data_out=16'h9f0;
17'hbd18:	data_out=16'h8a00;
17'hbd19:	data_out=16'h8a00;
17'hbd1a:	data_out=16'ha00;
17'hbd1b:	data_out=16'h646;
17'hbd1c:	data_out=16'ha00;
17'hbd1d:	data_out=16'h8a00;
17'hbd1e:	data_out=16'h8994;
17'hbd1f:	data_out=16'h9ff;
17'hbd20:	data_out=16'h899e;
17'hbd21:	data_out=16'ha00;
17'hbd22:	data_out=16'h89c4;
17'hbd23:	data_out=16'h8a00;
17'hbd24:	data_out=16'h8a00;
17'hbd25:	data_out=16'h89fe;
17'hbd26:	data_out=16'h8a00;
17'hbd27:	data_out=16'h8a00;
17'hbd28:	data_out=16'ha00;
17'hbd29:	data_out=16'h8a00;
17'hbd2a:	data_out=16'h89ff;
17'hbd2b:	data_out=16'h8a00;
17'hbd2c:	data_out=16'h8974;
17'hbd2d:	data_out=16'h8a00;
17'hbd2e:	data_out=16'h89c8;
17'hbd2f:	data_out=16'h88f6;
17'hbd30:	data_out=16'h80e;
17'hbd31:	data_out=16'h89e4;
17'hbd32:	data_out=16'h60d;
17'hbd33:	data_out=16'h80b;
17'hbd34:	data_out=16'h8a00;
17'hbd35:	data_out=16'h8a00;
17'hbd36:	data_out=16'h89ff;
17'hbd37:	data_out=16'h832c;
17'hbd38:	data_out=16'ha00;
17'hbd39:	data_out=16'h8621;
17'hbd3a:	data_out=16'h8a00;
17'hbd3b:	data_out=16'h8a00;
17'hbd3c:	data_out=16'h9bd;
17'hbd3d:	data_out=16'h89e8;
17'hbd3e:	data_out=16'ha00;
17'hbd3f:	data_out=16'ha00;
17'hbd40:	data_out=16'h87f6;
17'hbd41:	data_out=16'h885a;
17'hbd42:	data_out=16'h8a00;
17'hbd43:	data_out=16'ha00;
17'hbd44:	data_out=16'h89f4;
17'hbd45:	data_out=16'h89be;
17'hbd46:	data_out=16'h8a00;
17'hbd47:	data_out=16'h8a00;
17'hbd48:	data_out=16'h89ab;
17'hbd49:	data_out=16'h8a00;
17'hbd4a:	data_out=16'h8a00;
17'hbd4b:	data_out=16'h8a00;
17'hbd4c:	data_out=16'h89ff;
17'hbd4d:	data_out=16'h89df;
17'hbd4e:	data_out=16'h8a00;
17'hbd4f:	data_out=16'h8a00;
17'hbd50:	data_out=16'h821;
17'hbd51:	data_out=16'ha00;
17'hbd52:	data_out=16'h8a00;
17'hbd53:	data_out=16'h89d9;
17'hbd54:	data_out=16'h89ec;
17'hbd55:	data_out=16'h845;
17'hbd56:	data_out=16'h8a00;
17'hbd57:	data_out=16'h89f5;
17'hbd58:	data_out=16'ha00;
17'hbd59:	data_out=16'h895f;
17'hbd5a:	data_out=16'ha00;
17'hbd5b:	data_out=16'h89f9;
17'hbd5c:	data_out=16'ha00;
17'hbd5d:	data_out=16'h89af;
17'hbd5e:	data_out=16'h8752;
17'hbd5f:	data_out=16'h8a00;
17'hbd60:	data_out=16'h8a00;
17'hbd61:	data_out=16'h9f1;
17'hbd62:	data_out=16'h8937;
17'hbd63:	data_out=16'h9ff;
17'hbd64:	data_out=16'h8a00;
17'hbd65:	data_out=16'h89ff;
17'hbd66:	data_out=16'h8a00;
17'hbd67:	data_out=16'h8a00;
17'hbd68:	data_out=16'ha00;
17'hbd69:	data_out=16'h8a00;
17'hbd6a:	data_out=16'ha00;
17'hbd6b:	data_out=16'ha00;
17'hbd6c:	data_out=16'h89f3;
17'hbd6d:	data_out=16'h9ff;
17'hbd6e:	data_out=16'ha00;
17'hbd6f:	data_out=16'ha00;
17'hbd70:	data_out=16'ha00;
17'hbd71:	data_out=16'h89ff;
17'hbd72:	data_out=16'h9c1;
17'hbd73:	data_out=16'h9e4;
17'hbd74:	data_out=16'h8f1;
17'hbd75:	data_out=16'ha00;
17'hbd76:	data_out=16'h8a00;
17'hbd77:	data_out=16'h8a00;
17'hbd78:	data_out=16'ha00;
17'hbd79:	data_out=16'h89d9;
17'hbd7a:	data_out=16'h9ff;
17'hbd7b:	data_out=16'ha00;
17'hbd7c:	data_out=16'h8a00;
17'hbd7d:	data_out=16'ha00;
17'hbd7e:	data_out=16'h8127;
17'hbd7f:	data_out=16'ha00;
17'hbd80:	data_out=16'h89ff;
17'hbd81:	data_out=16'h8a00;
17'hbd82:	data_out=16'h8a00;
17'hbd83:	data_out=16'h963;
17'hbd84:	data_out=16'h8a00;
17'hbd85:	data_out=16'h9e8;
17'hbd86:	data_out=16'h9fe;
17'hbd87:	data_out=16'h8a00;
17'hbd88:	data_out=16'h8a00;
17'hbd89:	data_out=16'h8a00;
17'hbd8a:	data_out=16'h8a00;
17'hbd8b:	data_out=16'h8a00;
17'hbd8c:	data_out=16'h8a00;
17'hbd8d:	data_out=16'h98a;
17'hbd8e:	data_out=16'ha00;
17'hbd8f:	data_out=16'h8a00;
17'hbd90:	data_out=16'h8a00;
17'hbd91:	data_out=16'h8a00;
17'hbd92:	data_out=16'h8e2;
17'hbd93:	data_out=16'ha00;
17'hbd94:	data_out=16'h9dc;
17'hbd95:	data_out=16'h89ff;
17'hbd96:	data_out=16'h89fe;
17'hbd97:	data_out=16'h9d8;
17'hbd98:	data_out=16'h8a00;
17'hbd99:	data_out=16'h8a00;
17'hbd9a:	data_out=16'h9d5;
17'hbd9b:	data_out=16'h87f;
17'hbd9c:	data_out=16'h9c6;
17'hbd9d:	data_out=16'h8a00;
17'hbd9e:	data_out=16'h860f;
17'hbd9f:	data_out=16'h9fc;
17'hbda0:	data_out=16'h89f6;
17'hbda1:	data_out=16'ha00;
17'hbda2:	data_out=16'h8897;
17'hbda3:	data_out=16'h8a00;
17'hbda4:	data_out=16'h8a00;
17'hbda5:	data_out=16'h89ff;
17'hbda6:	data_out=16'h8a00;
17'hbda7:	data_out=16'h8a00;
17'hbda8:	data_out=16'ha00;
17'hbda9:	data_out=16'h8a1;
17'hbdaa:	data_out=16'h8a00;
17'hbdab:	data_out=16'h8a00;
17'hbdac:	data_out=16'h89fd;
17'hbdad:	data_out=16'h8a00;
17'hbdae:	data_out=16'h166;
17'hbdaf:	data_out=16'h8979;
17'hbdb0:	data_out=16'h8a00;
17'hbdb1:	data_out=16'h8a00;
17'hbdb2:	data_out=16'h8a00;
17'hbdb3:	data_out=16'ha00;
17'hbdb4:	data_out=16'h8a00;
17'hbdb5:	data_out=16'h8a00;
17'hbdb6:	data_out=16'h8a00;
17'hbdb7:	data_out=16'h8a00;
17'hbdb8:	data_out=16'ha00;
17'hbdb9:	data_out=16'ha00;
17'hbdba:	data_out=16'h8a00;
17'hbdbb:	data_out=16'h8a00;
17'hbdbc:	data_out=16'h94b;
17'hbdbd:	data_out=16'h89fe;
17'hbdbe:	data_out=16'ha00;
17'hbdbf:	data_out=16'h9e8;
17'hbdc0:	data_out=16'h8a00;
17'hbdc1:	data_out=16'h8a00;
17'hbdc2:	data_out=16'h8a00;
17'hbdc3:	data_out=16'ha00;
17'hbdc4:	data_out=16'h8a00;
17'hbdc5:	data_out=16'h89ff;
17'hbdc6:	data_out=16'h8a00;
17'hbdc7:	data_out=16'h8a00;
17'hbdc8:	data_out=16'h81cd;
17'hbdc9:	data_out=16'h8a00;
17'hbdca:	data_out=16'h8a00;
17'hbdcb:	data_out=16'h8a00;
17'hbdcc:	data_out=16'h8a00;
17'hbdcd:	data_out=16'h891b;
17'hbdce:	data_out=16'h8898;
17'hbdcf:	data_out=16'h8a00;
17'hbdd0:	data_out=16'h9b5;
17'hbdd1:	data_out=16'h9f9;
17'hbdd2:	data_out=16'h8a00;
17'hbdd3:	data_out=16'h8a00;
17'hbdd4:	data_out=16'h89fa;
17'hbdd5:	data_out=16'h930;
17'hbdd6:	data_out=16'h8a00;
17'hbdd7:	data_out=16'h8a00;
17'hbdd8:	data_out=16'ha00;
17'hbdd9:	data_out=16'h8a00;
17'hbdda:	data_out=16'h9fe;
17'hbddb:	data_out=16'h8a00;
17'hbddc:	data_out=16'ha00;
17'hbddd:	data_out=16'h89d1;
17'hbdde:	data_out=16'h86f2;
17'hbddf:	data_out=16'h8a00;
17'hbde0:	data_out=16'h8a00;
17'hbde1:	data_out=16'h8a00;
17'hbde2:	data_out=16'h9a8;
17'hbde3:	data_out=16'ha00;
17'hbde4:	data_out=16'h8a00;
17'hbde5:	data_out=16'h8a00;
17'hbde6:	data_out=16'h8a00;
17'hbde7:	data_out=16'h89c3;
17'hbde8:	data_out=16'ha00;
17'hbde9:	data_out=16'h8a00;
17'hbdea:	data_out=16'ha00;
17'hbdeb:	data_out=16'h898d;
17'hbdec:	data_out=16'h89fe;
17'hbded:	data_out=16'ha00;
17'hbdee:	data_out=16'ha00;
17'hbdef:	data_out=16'h9c1;
17'hbdf0:	data_out=16'ha00;
17'hbdf1:	data_out=16'h8a00;
17'hbdf2:	data_out=16'h8946;
17'hbdf3:	data_out=16'h842;
17'hbdf4:	data_out=16'h8a00;
17'hbdf5:	data_out=16'ha00;
17'hbdf6:	data_out=16'h8a00;
17'hbdf7:	data_out=16'h8a00;
17'hbdf8:	data_out=16'ha00;
17'hbdf9:	data_out=16'h89f9;
17'hbdfa:	data_out=16'h9f1;
17'hbdfb:	data_out=16'ha00;
17'hbdfc:	data_out=16'h89ff;
17'hbdfd:	data_out=16'h9ff;
17'hbdfe:	data_out=16'h386;
17'hbdff:	data_out=16'ha00;
17'hbe00:	data_out=16'h8a00;
17'hbe01:	data_out=16'h8a00;
17'hbe02:	data_out=16'h789;
17'hbe03:	data_out=16'h9f1;
17'hbe04:	data_out=16'h8a00;
17'hbe05:	data_out=16'h88e7;
17'hbe06:	data_out=16'h9fe;
17'hbe07:	data_out=16'h8a00;
17'hbe08:	data_out=16'h8a00;
17'hbe09:	data_out=16'h89e0;
17'hbe0a:	data_out=16'h8a00;
17'hbe0b:	data_out=16'h896d;
17'hbe0c:	data_out=16'h8a00;
17'hbe0d:	data_out=16'h9a7;
17'hbe0e:	data_out=16'ha00;
17'hbe0f:	data_out=16'h861d;
17'hbe10:	data_out=16'h896b;
17'hbe11:	data_out=16'h8a00;
17'hbe12:	data_out=16'h9e2;
17'hbe13:	data_out=16'h9fd;
17'hbe14:	data_out=16'h9fe;
17'hbe15:	data_out=16'h8a00;
17'hbe16:	data_out=16'h8a00;
17'hbe17:	data_out=16'ha00;
17'hbe18:	data_out=16'h8a00;
17'hbe19:	data_out=16'h8a00;
17'hbe1a:	data_out=16'h89fc;
17'hbe1b:	data_out=16'h9e2;
17'hbe1c:	data_out=16'ha00;
17'hbe1d:	data_out=16'h8a00;
17'hbe1e:	data_out=16'h9e5;
17'hbe1f:	data_out=16'h9f3;
17'hbe20:	data_out=16'h89ff;
17'hbe21:	data_out=16'ha00;
17'hbe22:	data_out=16'h9f0;
17'hbe23:	data_out=16'h8a00;
17'hbe24:	data_out=16'h8a00;
17'hbe25:	data_out=16'h89ea;
17'hbe26:	data_out=16'h8a00;
17'hbe27:	data_out=16'h8a00;
17'hbe28:	data_out=16'ha00;
17'hbe29:	data_out=16'h9de;
17'hbe2a:	data_out=16'h8a00;
17'hbe2b:	data_out=16'h8980;
17'hbe2c:	data_out=16'h8a00;
17'hbe2d:	data_out=16'h8a00;
17'hbe2e:	data_out=16'h9e8;
17'hbe2f:	data_out=16'h87bb;
17'hbe30:	data_out=16'h8a00;
17'hbe31:	data_out=16'h8a00;
17'hbe32:	data_out=16'h8a00;
17'hbe33:	data_out=16'ha00;
17'hbe34:	data_out=16'h8a00;
17'hbe35:	data_out=16'h8a00;
17'hbe36:	data_out=16'h8a00;
17'hbe37:	data_out=16'h9c5;
17'hbe38:	data_out=16'ha00;
17'hbe39:	data_out=16'ha00;
17'hbe3a:	data_out=16'h8a00;
17'hbe3b:	data_out=16'h8a00;
17'hbe3c:	data_out=16'h98e;
17'hbe3d:	data_out=16'h8a00;
17'hbe3e:	data_out=16'ha00;
17'hbe3f:	data_out=16'h8923;
17'hbe40:	data_out=16'h8a00;
17'hbe41:	data_out=16'h8a00;
17'hbe42:	data_out=16'h8a00;
17'hbe43:	data_out=16'ha00;
17'hbe44:	data_out=16'h8a00;
17'hbe45:	data_out=16'h8a00;
17'hbe46:	data_out=16'h8a00;
17'hbe47:	data_out=16'h8a00;
17'hbe48:	data_out=16'h9f6;
17'hbe49:	data_out=16'h8a00;
17'hbe4a:	data_out=16'h8a00;
17'hbe4b:	data_out=16'h8a00;
17'hbe4c:	data_out=16'h89d6;
17'hbe4d:	data_out=16'h9e3;
17'hbe4e:	data_out=16'h9a6;
17'hbe4f:	data_out=16'h8a00;
17'hbe50:	data_out=16'h9fd;
17'hbe51:	data_out=16'h9d0;
17'hbe52:	data_out=16'h8a00;
17'hbe53:	data_out=16'h89b7;
17'hbe54:	data_out=16'h89ff;
17'hbe55:	data_out=16'h9cf;
17'hbe56:	data_out=16'h8a00;
17'hbe57:	data_out=16'h8a00;
17'hbe58:	data_out=16'ha00;
17'hbe59:	data_out=16'h8a00;
17'hbe5a:	data_out=16'ha00;
17'hbe5b:	data_out=16'h8a00;
17'hbe5c:	data_out=16'ha00;
17'hbe5d:	data_out=16'h8963;
17'hbe5e:	data_out=16'h8515;
17'hbe5f:	data_out=16'h8a00;
17'hbe60:	data_out=16'h8a00;
17'hbe61:	data_out=16'h8a00;
17'hbe62:	data_out=16'h9f6;
17'hbe63:	data_out=16'ha00;
17'hbe64:	data_out=16'h8a00;
17'hbe65:	data_out=16'h8a00;
17'hbe66:	data_out=16'h89db;
17'hbe67:	data_out=16'h82e8;
17'hbe68:	data_out=16'ha00;
17'hbe69:	data_out=16'h8a00;
17'hbe6a:	data_out=16'ha00;
17'hbe6b:	data_out=16'h89e7;
17'hbe6c:	data_out=16'h8a00;
17'hbe6d:	data_out=16'ha00;
17'hbe6e:	data_out=16'ha00;
17'hbe6f:	data_out=16'h9c4;
17'hbe70:	data_out=16'ha00;
17'hbe71:	data_out=16'h8992;
17'hbe72:	data_out=16'h89f0;
17'hbe73:	data_out=16'h89f7;
17'hbe74:	data_out=16'h8a00;
17'hbe75:	data_out=16'h9d6;
17'hbe76:	data_out=16'h89be;
17'hbe77:	data_out=16'h89b5;
17'hbe78:	data_out=16'ha00;
17'hbe79:	data_out=16'h897a;
17'hbe7a:	data_out=16'ha00;
17'hbe7b:	data_out=16'ha00;
17'hbe7c:	data_out=16'h8a00;
17'hbe7d:	data_out=16'h9fa;
17'hbe7e:	data_out=16'h9fe;
17'hbe7f:	data_out=16'h5ee;
17'hbe80:	data_out=16'h8a00;
17'hbe81:	data_out=16'h8a00;
17'hbe82:	data_out=16'h9ef;
17'hbe83:	data_out=16'ha00;
17'hbe84:	data_out=16'h8a00;
17'hbe85:	data_out=16'h89cf;
17'hbe86:	data_out=16'h9fb;
17'hbe87:	data_out=16'h8a00;
17'hbe88:	data_out=16'h877e;
17'hbe89:	data_out=16'h9be;
17'hbe8a:	data_out=16'h8a00;
17'hbe8b:	data_out=16'ha00;
17'hbe8c:	data_out=16'h89b8;
17'hbe8d:	data_out=16'h98;
17'hbe8e:	data_out=16'ha00;
17'hbe8f:	data_out=16'h9e6;
17'hbe90:	data_out=16'h80e0;
17'hbe91:	data_out=16'h89fd;
17'hbe92:	data_out=16'h9e2;
17'hbe93:	data_out=16'h9fe;
17'hbe94:	data_out=16'ha00;
17'hbe95:	data_out=16'h8a00;
17'hbe96:	data_out=16'h89fa;
17'hbe97:	data_out=16'ha00;
17'hbe98:	data_out=16'h89f9;
17'hbe99:	data_out=16'h9e2;
17'hbe9a:	data_out=16'h89cf;
17'hbe9b:	data_out=16'ha00;
17'hbe9c:	data_out=16'h673;
17'hbe9d:	data_out=16'h8a00;
17'hbe9e:	data_out=16'h9fd;
17'hbe9f:	data_out=16'h9ce;
17'hbea0:	data_out=16'h89cb;
17'hbea1:	data_out=16'ha00;
17'hbea2:	data_out=16'h9fd;
17'hbea3:	data_out=16'h8a00;
17'hbea4:	data_out=16'h8a00;
17'hbea5:	data_out=16'h8984;
17'hbea6:	data_out=16'h8883;
17'hbea7:	data_out=16'h89f6;
17'hbea8:	data_out=16'ha00;
17'hbea9:	data_out=16'h9f1;
17'hbeaa:	data_out=16'h87f1;
17'hbeab:	data_out=16'h9ff;
17'hbeac:	data_out=16'h8a00;
17'hbead:	data_out=16'h89db;
17'hbeae:	data_out=16'h9ff;
17'hbeaf:	data_out=16'h86ed;
17'hbeb0:	data_out=16'h8961;
17'hbeb1:	data_out=16'h8a00;
17'hbeb2:	data_out=16'h89cb;
17'hbeb3:	data_out=16'ha00;
17'hbeb4:	data_out=16'h8a00;
17'hbeb5:	data_out=16'h8a00;
17'hbeb6:	data_out=16'h8894;
17'hbeb7:	data_out=16'h9f4;
17'hbeb8:	data_out=16'h899b;
17'hbeb9:	data_out=16'ha00;
17'hbeba:	data_out=16'h89f9;
17'hbebb:	data_out=16'h8a00;
17'hbebc:	data_out=16'h9ed;
17'hbebd:	data_out=16'h8a00;
17'hbebe:	data_out=16'ha00;
17'hbebf:	data_out=16'h89d3;
17'hbec0:	data_out=16'h89ac;
17'hbec1:	data_out=16'h89be;
17'hbec2:	data_out=16'h89f3;
17'hbec3:	data_out=16'ha00;
17'hbec4:	data_out=16'h8a00;
17'hbec5:	data_out=16'h8a00;
17'hbec6:	data_out=16'h9f7;
17'hbec7:	data_out=16'h89ca;
17'hbec8:	data_out=16'h9fe;
17'hbec9:	data_out=16'h89db;
17'hbeca:	data_out=16'h89c1;
17'hbecb:	data_out=16'h89ef;
17'hbecc:	data_out=16'h89a1;
17'hbecd:	data_out=16'h9fb;
17'hbece:	data_out=16'h9f5;
17'hbecf:	data_out=16'h89fe;
17'hbed0:	data_out=16'h86c2;
17'hbed1:	data_out=16'h9df;
17'hbed2:	data_out=16'h8a00;
17'hbed3:	data_out=16'h8740;
17'hbed4:	data_out=16'h896d;
17'hbed5:	data_out=16'h9fc;
17'hbed6:	data_out=16'h89fc;
17'hbed7:	data_out=16'h8518;
17'hbed8:	data_out=16'ha00;
17'hbed9:	data_out=16'h89b0;
17'hbeda:	data_out=16'ha00;
17'hbedb:	data_out=16'h8a00;
17'hbedc:	data_out=16'ha00;
17'hbedd:	data_out=16'h891b;
17'hbede:	data_out=16'h83f5;
17'hbedf:	data_out=16'h89e4;
17'hbee0:	data_out=16'h89f8;
17'hbee1:	data_out=16'h8a00;
17'hbee2:	data_out=16'h9fd;
17'hbee3:	data_out=16'ha00;
17'hbee4:	data_out=16'h8a00;
17'hbee5:	data_out=16'h89b1;
17'hbee6:	data_out=16'h9f6;
17'hbee7:	data_out=16'h76f;
17'hbee8:	data_out=16'ha00;
17'hbee9:	data_out=16'h3f;
17'hbeea:	data_out=16'ha00;
17'hbeeb:	data_out=16'h8971;
17'hbeec:	data_out=16'h8a00;
17'hbeed:	data_out=16'ha00;
17'hbeee:	data_out=16'ha00;
17'hbeef:	data_out=16'h897d;
17'hbef0:	data_out=16'ha00;
17'hbef1:	data_out=16'h9d0;
17'hbef2:	data_out=16'h89db;
17'hbef3:	data_out=16'h89e5;
17'hbef4:	data_out=16'h8a00;
17'hbef5:	data_out=16'h9df;
17'hbef6:	data_out=16'ha00;
17'hbef7:	data_out=16'h9f5;
17'hbef8:	data_out=16'ha00;
17'hbef9:	data_out=16'h25a;
17'hbefa:	data_out=16'ha00;
17'hbefb:	data_out=16'ha00;
17'hbefc:	data_out=16'h89fd;
17'hbefd:	data_out=16'h9f8;
17'hbefe:	data_out=16'h9ff;
17'hbeff:	data_out=16'h89e8;
17'hbf00:	data_out=16'h8a00;
17'hbf01:	data_out=16'h89b6;
17'hbf02:	data_out=16'h9f8;
17'hbf03:	data_out=16'h3d0;
17'hbf04:	data_out=16'h8a00;
17'hbf05:	data_out=16'h89cb;
17'hbf06:	data_out=16'h8070;
17'hbf07:	data_out=16'h993;
17'hbf08:	data_out=16'h3d5;
17'hbf09:	data_out=16'h9f8;
17'hbf0a:	data_out=16'h8994;
17'hbf0b:	data_out=16'ha00;
17'hbf0c:	data_out=16'h9fe;
17'hbf0d:	data_out=16'h89ed;
17'hbf0e:	data_out=16'h9fa;
17'hbf0f:	data_out=16'h9ee;
17'hbf10:	data_out=16'h61c;
17'hbf11:	data_out=16'h893d;
17'hbf12:	data_out=16'h974;
17'hbf13:	data_out=16'h4de;
17'hbf14:	data_out=16'ha00;
17'hbf15:	data_out=16'h8a00;
17'hbf16:	data_out=16'h89eb;
17'hbf17:	data_out=16'ha00;
17'hbf18:	data_out=16'h89fe;
17'hbf19:	data_out=16'ha00;
17'hbf1a:	data_out=16'h89cd;
17'hbf1b:	data_out=16'ha00;
17'hbf1c:	data_out=16'h865b;
17'hbf1d:	data_out=16'h89a9;
17'hbf1e:	data_out=16'h90f;
17'hbf1f:	data_out=16'h9c1;
17'hbf20:	data_out=16'h89b5;
17'hbf21:	data_out=16'h9fb;
17'hbf22:	data_out=16'h9e1;
17'hbf23:	data_out=16'h6c5;
17'hbf24:	data_out=16'h6bc;
17'hbf25:	data_out=16'h9d3;
17'hbf26:	data_out=16'ha00;
17'hbf27:	data_out=16'h8954;
17'hbf28:	data_out=16'h9fe;
17'hbf29:	data_out=16'h9f9;
17'hbf2a:	data_out=16'h839d;
17'hbf2b:	data_out=16'ha00;
17'hbf2c:	data_out=16'h89fa;
17'hbf2d:	data_out=16'h8291;
17'hbf2e:	data_out=16'ha00;
17'hbf2f:	data_out=16'h887d;
17'hbf30:	data_out=16'h38;
17'hbf31:	data_out=16'h89e6;
17'hbf32:	data_out=16'h8981;
17'hbf33:	data_out=16'ha00;
17'hbf34:	data_out=16'h89e9;
17'hbf35:	data_out=16'h892b;
17'hbf36:	data_out=16'ha7;
17'hbf37:	data_out=16'ha00;
17'hbf38:	data_out=16'h89f0;
17'hbf39:	data_out=16'ha00;
17'hbf3a:	data_out=16'h9db;
17'hbf3b:	data_out=16'h89b2;
17'hbf3c:	data_out=16'ha00;
17'hbf3d:	data_out=16'h89d3;
17'hbf3e:	data_out=16'h9fe;
17'hbf3f:	data_out=16'h89cf;
17'hbf40:	data_out=16'h89a6;
17'hbf41:	data_out=16'h680;
17'hbf42:	data_out=16'h8993;
17'hbf43:	data_out=16'h9f7;
17'hbf44:	data_out=16'h89cf;
17'hbf45:	data_out=16'h8a00;
17'hbf46:	data_out=16'ha00;
17'hbf47:	data_out=16'h967;
17'hbf48:	data_out=16'h9df;
17'hbf49:	data_out=16'h9e4;
17'hbf4a:	data_out=16'h833c;
17'hbf4b:	data_out=16'h89ae;
17'hbf4c:	data_out=16'h896f;
17'hbf4d:	data_out=16'h9e7;
17'hbf4e:	data_out=16'ha00;
17'hbf4f:	data_out=16'h8748;
17'hbf50:	data_out=16'h894a;
17'hbf51:	data_out=16'h9dd;
17'hbf52:	data_out=16'h87bb;
17'hbf53:	data_out=16'h56c;
17'hbf54:	data_out=16'h8967;
17'hbf55:	data_out=16'ha00;
17'hbf56:	data_out=16'h9f6;
17'hbf57:	data_out=16'h9a2;
17'hbf58:	data_out=16'ha00;
17'hbf59:	data_out=16'h89ac;
17'hbf5a:	data_out=16'ha00;
17'hbf5b:	data_out=16'h898b;
17'hbf5c:	data_out=16'h8536;
17'hbf5d:	data_out=16'h897b;
17'hbf5e:	data_out=16'h8686;
17'hbf5f:	data_out=16'h89ee;
17'hbf60:	data_out=16'h9e5;
17'hbf61:	data_out=16'h89ae;
17'hbf62:	data_out=16'ha00;
17'hbf63:	data_out=16'ha00;
17'hbf64:	data_out=16'h8a00;
17'hbf65:	data_out=16'h84fa;
17'hbf66:	data_out=16'ha00;
17'hbf67:	data_out=16'h9f2;
17'hbf68:	data_out=16'h9fc;
17'hbf69:	data_out=16'h9f4;
17'hbf6a:	data_out=16'h9f9;
17'hbf6b:	data_out=16'h8979;
17'hbf6c:	data_out=16'h8a00;
17'hbf6d:	data_out=16'ha00;
17'hbf6e:	data_out=16'h9f9;
17'hbf6f:	data_out=16'h89a4;
17'hbf70:	data_out=16'h9f9;
17'hbf71:	data_out=16'h50f;
17'hbf72:	data_out=16'h89e2;
17'hbf73:	data_out=16'h89bb;
17'hbf74:	data_out=16'h807e;
17'hbf75:	data_out=16'h8856;
17'hbf76:	data_out=16'ha00;
17'hbf77:	data_out=16'h9f9;
17'hbf78:	data_out=16'h9e5;
17'hbf79:	data_out=16'h9f2;
17'hbf7a:	data_out=16'ha00;
17'hbf7b:	data_out=16'h9fe;
17'hbf7c:	data_out=16'h8a00;
17'hbf7d:	data_out=16'h5ce;
17'hbf7e:	data_out=16'h56b;
17'hbf7f:	data_out=16'h8a00;
17'hbf80:	data_out=16'h8a00;
17'hbf81:	data_out=16'h8a00;
17'hbf82:	data_out=16'h8219;
17'hbf83:	data_out=16'h86ef;
17'hbf84:	data_out=16'h8a00;
17'hbf85:	data_out=16'h8a00;
17'hbf86:	data_out=16'h89e4;
17'hbf87:	data_out=16'h9f4;
17'hbf88:	data_out=16'h8352;
17'hbf89:	data_out=16'h9fd;
17'hbf8a:	data_out=16'h89ff;
17'hbf8b:	data_out=16'ha00;
17'hbf8c:	data_out=16'h9f8;
17'hbf8d:	data_out=16'h89ff;
17'hbf8e:	data_out=16'h8177;
17'hbf8f:	data_out=16'h8861;
17'hbf90:	data_out=16'h9e5;
17'hbf91:	data_out=16'h89fd;
17'hbf92:	data_out=16'h89b7;
17'hbf93:	data_out=16'h8775;
17'hbf94:	data_out=16'h826c;
17'hbf95:	data_out=16'h8a00;
17'hbf96:	data_out=16'h8a00;
17'hbf97:	data_out=16'h854e;
17'hbf98:	data_out=16'h89ff;
17'hbf99:	data_out=16'ha00;
17'hbf9a:	data_out=16'h8a00;
17'hbf9b:	data_out=16'h378;
17'hbf9c:	data_out=16'h89b4;
17'hbf9d:	data_out=16'h89ee;
17'hbf9e:	data_out=16'h882f;
17'hbf9f:	data_out=16'h89f6;
17'hbfa0:	data_out=16'h89fb;
17'hbfa1:	data_out=16'h8060;
17'hbfa2:	data_out=16'h9eb;
17'hbfa3:	data_out=16'ha00;
17'hbfa4:	data_out=16'ha00;
17'hbfa5:	data_out=16'h9d7;
17'hbfa6:	data_out=16'ha00;
17'hbfa7:	data_out=16'h89d0;
17'hbfa8:	data_out=16'h21d;
17'hbfa9:	data_out=16'ha00;
17'hbfaa:	data_out=16'h8887;
17'hbfab:	data_out=16'ha00;
17'hbfac:	data_out=16'h8a00;
17'hbfad:	data_out=16'h9f5;
17'hbfae:	data_out=16'h8639;
17'hbfaf:	data_out=16'h89a2;
17'hbfb0:	data_out=16'h83ac;
17'hbfb1:	data_out=16'h8a00;
17'hbfb2:	data_out=16'h89e3;
17'hbfb3:	data_out=16'h842c;
17'hbfb4:	data_out=16'h89f4;
17'hbfb5:	data_out=16'h89eb;
17'hbfb6:	data_out=16'h83d0;
17'hbfb7:	data_out=16'h93b;
17'hbfb8:	data_out=16'h8a00;
17'hbfb9:	data_out=16'h8629;
17'hbfba:	data_out=16'h9fe;
17'hbfbb:	data_out=16'h89ec;
17'hbfbc:	data_out=16'h5dc;
17'hbfbd:	data_out=16'h89f6;
17'hbfbe:	data_out=16'h228;
17'hbfbf:	data_out=16'h8a00;
17'hbfc0:	data_out=16'h8a00;
17'hbfc1:	data_out=16'h8984;
17'hbfc2:	data_out=16'h8824;
17'hbfc3:	data_out=16'h4ef;
17'hbfc4:	data_out=16'h8a00;
17'hbfc5:	data_out=16'h8a00;
17'hbfc6:	data_out=16'ha00;
17'hbfc7:	data_out=16'h9bd;
17'hbfc8:	data_out=16'h88cf;
17'hbfc9:	data_out=16'h9e1;
17'hbfca:	data_out=16'h843d;
17'hbfcb:	data_out=16'h89a2;
17'hbfcc:	data_out=16'hd4;
17'hbfcd:	data_out=16'h9f8;
17'hbfce:	data_out=16'ha00;
17'hbfcf:	data_out=16'h9f5;
17'hbfd0:	data_out=16'h89df;
17'hbfd1:	data_out=16'h89f4;
17'hbfd2:	data_out=16'h9d7;
17'hbfd3:	data_out=16'h862d;
17'hbfd4:	data_out=16'h89bb;
17'hbfd5:	data_out=16'h3c6;
17'hbfd6:	data_out=16'h278;
17'hbfd7:	data_out=16'h84e5;
17'hbfd8:	data_out=16'h8751;
17'hbfd9:	data_out=16'h89fd;
17'hbfda:	data_out=16'h969;
17'hbfdb:	data_out=16'h89fa;
17'hbfdc:	data_out=16'h89b9;
17'hbfdd:	data_out=16'h89d8;
17'hbfde:	data_out=16'h89a1;
17'hbfdf:	data_out=16'h89f8;
17'hbfe0:	data_out=16'h9ec;
17'hbfe1:	data_out=16'h8a00;
17'hbfe2:	data_out=16'h85cb;
17'hbfe3:	data_out=16'h84c0;
17'hbfe4:	data_out=16'h89ff;
17'hbfe5:	data_out=16'h8820;
17'hbfe6:	data_out=16'ha00;
17'hbfe7:	data_out=16'ha00;
17'hbfe8:	data_out=16'h97;
17'hbfe9:	data_out=16'h9f9;
17'hbfea:	data_out=16'h820b;
17'hbfeb:	data_out=16'h8a00;
17'hbfec:	data_out=16'h8a00;
17'hbfed:	data_out=16'h84ac;
17'hbfee:	data_out=16'h8209;
17'hbfef:	data_out=16'h8a00;
17'hbff0:	data_out=16'h81bc;
17'hbff1:	data_out=16'h89b8;
17'hbff2:	data_out=16'h8a00;
17'hbff3:	data_out=16'h8a00;
17'hbff4:	data_out=16'h83a4;
17'hbff5:	data_out=16'h89fe;
17'hbff6:	data_out=16'ha00;
17'hbff7:	data_out=16'h14d;
17'hbff8:	data_out=16'h100;
17'hbff9:	data_out=16'h825b;
17'hbffa:	data_out=16'h843e;
17'hbffb:	data_out=16'h22b;
17'hbffc:	data_out=16'h8a00;
17'hbffd:	data_out=16'h89f8;
17'hbffe:	data_out=16'h835f;
17'hbfff:	data_out=16'h8a00;
17'hc000:	data_out=16'h89ff;
17'hc001:	data_out=16'h8a00;
17'hc002:	data_out=16'h89b7;
17'hc003:	data_out=16'h87b3;
17'hc004:	data_out=16'h8a00;
17'hc005:	data_out=16'h8a00;
17'hc006:	data_out=16'h8a00;
17'hc007:	data_out=16'h9fa;
17'hc008:	data_out=16'h89a6;
17'hc009:	data_out=16'ha00;
17'hc00a:	data_out=16'h8a00;
17'hc00b:	data_out=16'ha00;
17'hc00c:	data_out=16'h9f9;
17'hc00d:	data_out=16'h89fe;
17'hc00e:	data_out=16'h89e7;
17'hc00f:	data_out=16'h88e2;
17'hc010:	data_out=16'h9ab;
17'hc011:	data_out=16'h8a00;
17'hc012:	data_out=16'h89f4;
17'hc013:	data_out=16'h84cc;
17'hc014:	data_out=16'h8913;
17'hc015:	data_out=16'h8a00;
17'hc016:	data_out=16'h8a00;
17'hc017:	data_out=16'h8895;
17'hc018:	data_out=16'h89ff;
17'hc019:	data_out=16'ha00;
17'hc01a:	data_out=16'h8a00;
17'hc01b:	data_out=16'h8647;
17'hc01c:	data_out=16'h89fb;
17'hc01d:	data_out=16'h89ea;
17'hc01e:	data_out=16'h89f2;
17'hc01f:	data_out=16'h89fc;
17'hc020:	data_out=16'h89ff;
17'hc021:	data_out=16'h89f5;
17'hc022:	data_out=16'h9ed;
17'hc023:	data_out=16'ha00;
17'hc024:	data_out=16'ha00;
17'hc025:	data_out=16'h9be;
17'hc026:	data_out=16'ha00;
17'hc027:	data_out=16'h8a00;
17'hc028:	data_out=16'h89fe;
17'hc029:	data_out=16'ha00;
17'hc02a:	data_out=16'h841b;
17'hc02b:	data_out=16'ha00;
17'hc02c:	data_out=16'h8a00;
17'hc02d:	data_out=16'ha00;
17'hc02e:	data_out=16'h8785;
17'hc02f:	data_out=16'h89fd;
17'hc030:	data_out=16'h89b7;
17'hc031:	data_out=16'h8a00;
17'hc032:	data_out=16'h89ff;
17'hc033:	data_out=16'h89f3;
17'hc034:	data_out=16'h89ce;
17'hc035:	data_out=16'h8a00;
17'hc036:	data_out=16'h87e0;
17'hc037:	data_out=16'h887b;
17'hc038:	data_out=16'h8a00;
17'hc039:	data_out=16'h89f2;
17'hc03a:	data_out=16'h9f5;
17'hc03b:	data_out=16'h8a00;
17'hc03c:	data_out=16'h808e;
17'hc03d:	data_out=16'h89f8;
17'hc03e:	data_out=16'h89fe;
17'hc03f:	data_out=16'h8a00;
17'hc040:	data_out=16'h8a00;
17'hc041:	data_out=16'h8a00;
17'hc042:	data_out=16'h9fa;
17'hc043:	data_out=16'h89ec;
17'hc044:	data_out=16'h8a00;
17'hc045:	data_out=16'h8a00;
17'hc046:	data_out=16'ha00;
17'hc047:	data_out=16'h9fa;
17'hc048:	data_out=16'h89fa;
17'hc049:	data_out=16'h9d0;
17'hc04a:	data_out=16'h89de;
17'hc04b:	data_out=16'h9f2;
17'hc04c:	data_out=16'h9f0;
17'hc04d:	data_out=16'h9ee;
17'hc04e:	data_out=16'h8064;
17'hc04f:	data_out=16'ha00;
17'hc050:	data_out=16'h8a00;
17'hc051:	data_out=16'h89fb;
17'hc052:	data_out=16'ha00;
17'hc053:	data_out=16'h89fc;
17'hc054:	data_out=16'h89f6;
17'hc055:	data_out=16'h88a1;
17'hc056:	data_out=16'h890f;
17'hc057:	data_out=16'h89ee;
17'hc058:	data_out=16'h89f6;
17'hc059:	data_out=16'h89fb;
17'hc05a:	data_out=16'h893f;
17'hc05b:	data_out=16'h8a00;
17'hc05c:	data_out=16'h8a00;
17'hc05d:	data_out=16'h89f9;
17'hc05e:	data_out=16'h89fd;
17'hc05f:	data_out=16'h89fd;
17'hc060:	data_out=16'h9fc;
17'hc061:	data_out=16'h8a00;
17'hc062:	data_out=16'h8332;
17'hc063:	data_out=16'h89f5;
17'hc064:	data_out=16'h84a6;
17'hc065:	data_out=16'h89e9;
17'hc066:	data_out=16'ha00;
17'hc067:	data_out=16'ha00;
17'hc068:	data_out=16'h89f8;
17'hc069:	data_out=16'h80f6;
17'hc06a:	data_out=16'h89d6;
17'hc06b:	data_out=16'h8a00;
17'hc06c:	data_out=16'h8a00;
17'hc06d:	data_out=16'h89f4;
17'hc06e:	data_out=16'h89d6;
17'hc06f:	data_out=16'h8a00;
17'hc070:	data_out=16'h89e0;
17'hc071:	data_out=16'h89f8;
17'hc072:	data_out=16'h8a00;
17'hc073:	data_out=16'h8a00;
17'hc074:	data_out=16'h89ac;
17'hc075:	data_out=16'h8a00;
17'hc076:	data_out=16'ha00;
17'hc077:	data_out=16'h881a;
17'hc078:	data_out=16'h8931;
17'hc079:	data_out=16'h89dd;
17'hc07a:	data_out=16'h89e1;
17'hc07b:	data_out=16'h89fe;
17'hc07c:	data_out=16'h8a00;
17'hc07d:	data_out=16'h8a00;
17'hc07e:	data_out=16'h185;
17'hc07f:	data_out=16'h8a00;
17'hc080:	data_out=16'h8a00;
17'hc081:	data_out=16'h8a00;
17'hc082:	data_out=16'h8a00;
17'hc083:	data_out=16'h881c;
17'hc084:	data_out=16'h8a00;
17'hc085:	data_out=16'h8a00;
17'hc086:	data_out=16'h678;
17'hc087:	data_out=16'ha00;
17'hc088:	data_out=16'h8a00;
17'hc089:	data_out=16'ha00;
17'hc08a:	data_out=16'h89fe;
17'hc08b:	data_out=16'ha00;
17'hc08c:	data_out=16'ha00;
17'hc08d:	data_out=16'h8a00;
17'hc08e:	data_out=16'h8a00;
17'hc08f:	data_out=16'h89e2;
17'hc090:	data_out=16'h995;
17'hc091:	data_out=16'h8a00;
17'hc092:	data_out=16'h8a00;
17'hc093:	data_out=16'h622;
17'hc094:	data_out=16'h89fa;
17'hc095:	data_out=16'h8a00;
17'hc096:	data_out=16'h8a00;
17'hc097:	data_out=16'h8930;
17'hc098:	data_out=16'h8a00;
17'hc099:	data_out=16'ha00;
17'hc09a:	data_out=16'h8a00;
17'hc09b:	data_out=16'h89fc;
17'hc09c:	data_out=16'h8a00;
17'hc09d:	data_out=16'h89d4;
17'hc09e:	data_out=16'h89fd;
17'hc09f:	data_out=16'h8a00;
17'hc0a0:	data_out=16'h8a00;
17'hc0a1:	data_out=16'h8a00;
17'hc0a2:	data_out=16'h9f3;
17'hc0a3:	data_out=16'ha00;
17'hc0a4:	data_out=16'ha00;
17'hc0a5:	data_out=16'h9b1;
17'hc0a6:	data_out=16'ha00;
17'hc0a7:	data_out=16'h8a00;
17'hc0a8:	data_out=16'h8a00;
17'hc0a9:	data_out=16'h9f5;
17'hc0aa:	data_out=16'h838a;
17'hc0ab:	data_out=16'h9f8;
17'hc0ac:	data_out=16'h8a00;
17'hc0ad:	data_out=16'ha00;
17'hc0ae:	data_out=16'h84d7;
17'hc0af:	data_out=16'h8a00;
17'hc0b0:	data_out=16'h89d0;
17'hc0b1:	data_out=16'h8a00;
17'hc0b2:	data_out=16'h89e0;
17'hc0b3:	data_out=16'h8a00;
17'hc0b4:	data_out=16'h89bf;
17'hc0b5:	data_out=16'h8a00;
17'hc0b6:	data_out=16'h89ff;
17'hc0b7:	data_out=16'h8a00;
17'hc0b8:	data_out=16'h8a00;
17'hc0b9:	data_out=16'h8a00;
17'hc0ba:	data_out=16'ha00;
17'hc0bb:	data_out=16'h8a00;
17'hc0bc:	data_out=16'h8755;
17'hc0bd:	data_out=16'h8a00;
17'hc0be:	data_out=16'h8a00;
17'hc0bf:	data_out=16'h8a00;
17'hc0c0:	data_out=16'h89ff;
17'hc0c1:	data_out=16'h8a00;
17'hc0c2:	data_out=16'ha00;
17'hc0c3:	data_out=16'h89d7;
17'hc0c4:	data_out=16'h8a00;
17'hc0c5:	data_out=16'h8a00;
17'hc0c6:	data_out=16'h5d;
17'hc0c7:	data_out=16'ha00;
17'hc0c8:	data_out=16'h2be;
17'hc0c9:	data_out=16'h9d0;
17'hc0ca:	data_out=16'h8847;
17'hc0cb:	data_out=16'ha00;
17'hc0cc:	data_out=16'ha00;
17'hc0cd:	data_out=16'h9f0;
17'hc0ce:	data_out=16'h87d6;
17'hc0cf:	data_out=16'ha00;
17'hc0d0:	data_out=16'h89fc;
17'hc0d1:	data_out=16'h8a00;
17'hc0d2:	data_out=16'ha00;
17'hc0d3:	data_out=16'h8a00;
17'hc0d4:	data_out=16'h8a00;
17'hc0d5:	data_out=16'h89d7;
17'hc0d6:	data_out=16'h8a00;
17'hc0d7:	data_out=16'h8a00;
17'hc0d8:	data_out=16'h8a00;
17'hc0d9:	data_out=16'h89fa;
17'hc0da:	data_out=16'h8a00;
17'hc0db:	data_out=16'h8a00;
17'hc0dc:	data_out=16'h8a00;
17'hc0dd:	data_out=16'h89ff;
17'hc0de:	data_out=16'h89ff;
17'hc0df:	data_out=16'h8a00;
17'hc0e0:	data_out=16'ha00;
17'hc0e1:	data_out=16'h8a00;
17'hc0e2:	data_out=16'ha00;
17'hc0e3:	data_out=16'h8a00;
17'hc0e4:	data_out=16'h80fd;
17'hc0e5:	data_out=16'h89df;
17'hc0e6:	data_out=16'ha00;
17'hc0e7:	data_out=16'ha00;
17'hc0e8:	data_out=16'h8a00;
17'hc0e9:	data_out=16'h89f8;
17'hc0ea:	data_out=16'h8a00;
17'hc0eb:	data_out=16'h8a00;
17'hc0ec:	data_out=16'h8a00;
17'hc0ed:	data_out=16'h8a00;
17'hc0ee:	data_out=16'h8a00;
17'hc0ef:	data_out=16'h8a00;
17'hc0f0:	data_out=16'h8a00;
17'hc0f1:	data_out=16'h89ff;
17'hc0f2:	data_out=16'h8a00;
17'hc0f3:	data_out=16'h8a00;
17'hc0f4:	data_out=16'h89da;
17'hc0f5:	data_out=16'h8a00;
17'hc0f6:	data_out=16'ha00;
17'hc0f7:	data_out=16'h82ef;
17'hc0f8:	data_out=16'h9f3;
17'hc0f9:	data_out=16'h8a00;
17'hc0fa:	data_out=16'h89ff;
17'hc0fb:	data_out=16'h8a00;
17'hc0fc:	data_out=16'h8a00;
17'hc0fd:	data_out=16'h8a00;
17'hc0fe:	data_out=16'h9e7;
17'hc0ff:	data_out=16'h8a00;
17'hc100:	data_out=16'h8a00;
17'hc101:	data_out=16'h8a00;
17'hc102:	data_out=16'h8a00;
17'hc103:	data_out=16'h8802;
17'hc104:	data_out=16'h8a00;
17'hc105:	data_out=16'h8a00;
17'hc106:	data_out=16'h91e;
17'hc107:	data_out=16'ha00;
17'hc108:	data_out=16'h8a00;
17'hc109:	data_out=16'ha00;
17'hc10a:	data_out=16'h89ee;
17'hc10b:	data_out=16'ha00;
17'hc10c:	data_out=16'ha00;
17'hc10d:	data_out=16'h8a00;
17'hc10e:	data_out=16'h8a00;
17'hc10f:	data_out=16'h89da;
17'hc110:	data_out=16'h89d8;
17'hc111:	data_out=16'h8a00;
17'hc112:	data_out=16'h8a00;
17'hc113:	data_out=16'h9fd;
17'hc114:	data_out=16'h89fd;
17'hc115:	data_out=16'h8a00;
17'hc116:	data_out=16'h8a00;
17'hc117:	data_out=16'h8391;
17'hc118:	data_out=16'h8a00;
17'hc119:	data_out=16'ha00;
17'hc11a:	data_out=16'h8a00;
17'hc11b:	data_out=16'h89ff;
17'hc11c:	data_out=16'h8a00;
17'hc11d:	data_out=16'h89c1;
17'hc11e:	data_out=16'h8a00;
17'hc11f:	data_out=16'h8a00;
17'hc120:	data_out=16'h8a00;
17'hc121:	data_out=16'h8a00;
17'hc122:	data_out=16'ha00;
17'hc123:	data_out=16'ha00;
17'hc124:	data_out=16'h9ff;
17'hc125:	data_out=16'h855;
17'hc126:	data_out=16'ha00;
17'hc127:	data_out=16'h8a00;
17'hc128:	data_out=16'h8a00;
17'hc129:	data_out=16'h9fe;
17'hc12a:	data_out=16'h7ad;
17'hc12b:	data_out=16'h9f5;
17'hc12c:	data_out=16'h8a00;
17'hc12d:	data_out=16'ha00;
17'hc12e:	data_out=16'h594;
17'hc12f:	data_out=16'h8a00;
17'hc130:	data_out=16'h891;
17'hc131:	data_out=16'h8a00;
17'hc132:	data_out=16'h7f6;
17'hc133:	data_out=16'h8a00;
17'hc134:	data_out=16'h9ca;
17'hc135:	data_out=16'h8a00;
17'hc136:	data_out=16'h8a00;
17'hc137:	data_out=16'h8a00;
17'hc138:	data_out=16'h8a00;
17'hc139:	data_out=16'h8a00;
17'hc13a:	data_out=16'ha00;
17'hc13b:	data_out=16'h89ff;
17'hc13c:	data_out=16'h844e;
17'hc13d:	data_out=16'h8a00;
17'hc13e:	data_out=16'h8a00;
17'hc13f:	data_out=16'h8a00;
17'hc140:	data_out=16'h89fe;
17'hc141:	data_out=16'h8a00;
17'hc142:	data_out=16'ha00;
17'hc143:	data_out=16'h1a6;
17'hc144:	data_out=16'h8a00;
17'hc145:	data_out=16'h8a00;
17'hc146:	data_out=16'h80e7;
17'hc147:	data_out=16'ha00;
17'hc148:	data_out=16'h9e1;
17'hc149:	data_out=16'h81b;
17'hc14a:	data_out=16'h901;
17'hc14b:	data_out=16'ha00;
17'hc14c:	data_out=16'ha00;
17'hc14d:	data_out=16'h958;
17'hc14e:	data_out=16'h88c0;
17'hc14f:	data_out=16'ha00;
17'hc150:	data_out=16'h89ff;
17'hc151:	data_out=16'h8a00;
17'hc152:	data_out=16'ha00;
17'hc153:	data_out=16'h8a00;
17'hc154:	data_out=16'h8a00;
17'hc155:	data_out=16'h88fb;
17'hc156:	data_out=16'h8a00;
17'hc157:	data_out=16'h8a00;
17'hc158:	data_out=16'h8a00;
17'hc159:	data_out=16'h8a00;
17'hc15a:	data_out=16'h8a00;
17'hc15b:	data_out=16'h8a00;
17'hc15c:	data_out=16'h8a00;
17'hc15d:	data_out=16'h8a00;
17'hc15e:	data_out=16'h8a00;
17'hc15f:	data_out=16'h8a00;
17'hc160:	data_out=16'ha00;
17'hc161:	data_out=16'h8a00;
17'hc162:	data_out=16'ha00;
17'hc163:	data_out=16'h8a00;
17'hc164:	data_out=16'h9d2;
17'hc165:	data_out=16'h9bf;
17'hc166:	data_out=16'h9f6;
17'hc167:	data_out=16'ha00;
17'hc168:	data_out=16'h8a00;
17'hc169:	data_out=16'h89fb;
17'hc16a:	data_out=16'h8a00;
17'hc16b:	data_out=16'h8a00;
17'hc16c:	data_out=16'h8a00;
17'hc16d:	data_out=16'h8a00;
17'hc16e:	data_out=16'h8a00;
17'hc16f:	data_out=16'h6c2;
17'hc170:	data_out=16'h8a00;
17'hc171:	data_out=16'h89e8;
17'hc172:	data_out=16'h8a00;
17'hc173:	data_out=16'h8a00;
17'hc174:	data_out=16'h87d;
17'hc175:	data_out=16'h8a00;
17'hc176:	data_out=16'ha00;
17'hc177:	data_out=16'h81b7;
17'hc178:	data_out=16'h9fe;
17'hc179:	data_out=16'h8a00;
17'hc17a:	data_out=16'h8a00;
17'hc17b:	data_out=16'h8a00;
17'hc17c:	data_out=16'h8a00;
17'hc17d:	data_out=16'h8a00;
17'hc17e:	data_out=16'h9dc;
17'hc17f:	data_out=16'h8a00;
17'hc180:	data_out=16'h8a00;
17'hc181:	data_out=16'h8a00;
17'hc182:	data_out=16'h8a00;
17'hc183:	data_out=16'h896d;
17'hc184:	data_out=16'h89ff;
17'hc185:	data_out=16'h8a00;
17'hc186:	data_out=16'ha00;
17'hc187:	data_out=16'ha00;
17'hc188:	data_out=16'h8a00;
17'hc189:	data_out=16'ha00;
17'hc18a:	data_out=16'h820d;
17'hc18b:	data_out=16'ha00;
17'hc18c:	data_out=16'ha00;
17'hc18d:	data_out=16'h8a00;
17'hc18e:	data_out=16'h8a00;
17'hc18f:	data_out=16'h89ef;
17'hc190:	data_out=16'h89d6;
17'hc191:	data_out=16'h8a00;
17'hc192:	data_out=16'h8a00;
17'hc193:	data_out=16'h9b1;
17'hc194:	data_out=16'h89f7;
17'hc195:	data_out=16'h8a00;
17'hc196:	data_out=16'h89ff;
17'hc197:	data_out=16'h8218;
17'hc198:	data_out=16'h8a00;
17'hc199:	data_out=16'ha00;
17'hc19a:	data_out=16'h89f5;
17'hc19b:	data_out=16'h8a00;
17'hc19c:	data_out=16'h8a00;
17'hc19d:	data_out=16'h89d6;
17'hc19e:	data_out=16'h8a00;
17'hc19f:	data_out=16'h89ec;
17'hc1a0:	data_out=16'h8a00;
17'hc1a1:	data_out=16'h8a00;
17'hc1a2:	data_out=16'ha00;
17'hc1a3:	data_out=16'h965;
17'hc1a4:	data_out=16'h945;
17'hc1a5:	data_out=16'h9b8;
17'hc1a6:	data_out=16'h9fb;
17'hc1a7:	data_out=16'h8a00;
17'hc1a8:	data_out=16'h8a00;
17'hc1a9:	data_out=16'h84fd;
17'hc1aa:	data_out=16'h4d8;
17'hc1ab:	data_out=16'h9e6;
17'hc1ac:	data_out=16'h8a00;
17'hc1ad:	data_out=16'ha00;
17'hc1ae:	data_out=16'h814;
17'hc1af:	data_out=16'h8a00;
17'hc1b0:	data_out=16'ha00;
17'hc1b1:	data_out=16'h8a00;
17'hc1b2:	data_out=16'ha00;
17'hc1b3:	data_out=16'h8a00;
17'hc1b4:	data_out=16'h30;
17'hc1b5:	data_out=16'h8a00;
17'hc1b6:	data_out=16'h8a00;
17'hc1b7:	data_out=16'h8a00;
17'hc1b8:	data_out=16'h8a00;
17'hc1b9:	data_out=16'h8a00;
17'hc1ba:	data_out=16'ha00;
17'hc1bb:	data_out=16'h9d3;
17'hc1bc:	data_out=16'h88ab;
17'hc1bd:	data_out=16'h8a00;
17'hc1be:	data_out=16'h8a00;
17'hc1bf:	data_out=16'h8a00;
17'hc1c0:	data_out=16'h801;
17'hc1c1:	data_out=16'h8a00;
17'hc1c2:	data_out=16'ha00;
17'hc1c3:	data_out=16'h964;
17'hc1c4:	data_out=16'h8a00;
17'hc1c5:	data_out=16'h8a00;
17'hc1c6:	data_out=16'h8a00;
17'hc1c7:	data_out=16'ha00;
17'hc1c8:	data_out=16'ha00;
17'hc1c9:	data_out=16'h943;
17'hc1ca:	data_out=16'h9f1;
17'hc1cb:	data_out=16'ha00;
17'hc1cc:	data_out=16'ha00;
17'hc1cd:	data_out=16'h93e;
17'hc1ce:	data_out=16'h842e;
17'hc1cf:	data_out=16'ha00;
17'hc1d0:	data_out=16'h89c0;
17'hc1d1:	data_out=16'h8a00;
17'hc1d2:	data_out=16'ha00;
17'hc1d3:	data_out=16'h8a00;
17'hc1d4:	data_out=16'h8a00;
17'hc1d5:	data_out=16'h8961;
17'hc1d6:	data_out=16'h8a00;
17'hc1d7:	data_out=16'h8a00;
17'hc1d8:	data_out=16'h8a00;
17'hc1d9:	data_out=16'h89c0;
17'hc1da:	data_out=16'h8a00;
17'hc1db:	data_out=16'h8a00;
17'hc1dc:	data_out=16'h8a00;
17'hc1dd:	data_out=16'h8a00;
17'hc1de:	data_out=16'h89ef;
17'hc1df:	data_out=16'h8a00;
17'hc1e0:	data_out=16'ha00;
17'hc1e1:	data_out=16'h8a00;
17'hc1e2:	data_out=16'ha00;
17'hc1e3:	data_out=16'h8a00;
17'hc1e4:	data_out=16'h960;
17'hc1e5:	data_out=16'ha00;
17'hc1e6:	data_out=16'h9ff;
17'hc1e7:	data_out=16'ha00;
17'hc1e8:	data_out=16'h8a00;
17'hc1e9:	data_out=16'h8a00;
17'hc1ea:	data_out=16'h8a00;
17'hc1eb:	data_out=16'h8a00;
17'hc1ec:	data_out=16'h8a00;
17'hc1ed:	data_out=16'h8a00;
17'hc1ee:	data_out=16'h8a00;
17'hc1ef:	data_out=16'ha00;
17'hc1f0:	data_out=16'h8a00;
17'hc1f1:	data_out=16'h89ed;
17'hc1f2:	data_out=16'h89f6;
17'hc1f3:	data_out=16'h89d6;
17'hc1f4:	data_out=16'h9ff;
17'hc1f5:	data_out=16'h8a00;
17'hc1f6:	data_out=16'ha00;
17'hc1f7:	data_out=16'he6;
17'hc1f8:	data_out=16'ha00;
17'hc1f9:	data_out=16'h8a00;
17'hc1fa:	data_out=16'h8a00;
17'hc1fb:	data_out=16'h8a00;
17'hc1fc:	data_out=16'h8a00;
17'hc1fd:	data_out=16'h8a00;
17'hc1fe:	data_out=16'h9fd;
17'hc1ff:	data_out=16'h8a00;
17'hc200:	data_out=16'h8a00;
17'hc201:	data_out=16'h8a00;
17'hc202:	data_out=16'h8a00;
17'hc203:	data_out=16'h89f8;
17'hc204:	data_out=16'h956;
17'hc205:	data_out=16'h8a00;
17'hc206:	data_out=16'ha00;
17'hc207:	data_out=16'ha00;
17'hc208:	data_out=16'h8a00;
17'hc209:	data_out=16'ha00;
17'hc20a:	data_out=16'h8298;
17'hc20b:	data_out=16'ha00;
17'hc20c:	data_out=16'ha00;
17'hc20d:	data_out=16'h8a00;
17'hc20e:	data_out=16'h8a00;
17'hc20f:	data_out=16'h89fa;
17'hc210:	data_out=16'h89c0;
17'hc211:	data_out=16'h50f;
17'hc212:	data_out=16'h82bd;
17'hc213:	data_out=16'h26a;
17'hc214:	data_out=16'h89fb;
17'hc215:	data_out=16'h8a00;
17'hc216:	data_out=16'h8a00;
17'hc217:	data_out=16'h89f1;
17'hc218:	data_out=16'h8a00;
17'hc219:	data_out=16'ha00;
17'hc21a:	data_out=16'h8e9;
17'hc21b:	data_out=16'h8a00;
17'hc21c:	data_out=16'h8a00;
17'hc21d:	data_out=16'h88ee;
17'hc21e:	data_out=16'h8a00;
17'hc21f:	data_out=16'h89ea;
17'hc220:	data_out=16'h8a00;
17'hc221:	data_out=16'h8a00;
17'hc222:	data_out=16'ha00;
17'hc223:	data_out=16'h84ce;
17'hc224:	data_out=16'h84f3;
17'hc225:	data_out=16'h9b2;
17'hc226:	data_out=16'h80e5;
17'hc227:	data_out=16'h89ff;
17'hc228:	data_out=16'h8a00;
17'hc229:	data_out=16'h8a00;
17'hc22a:	data_out=16'h88cf;
17'hc22b:	data_out=16'h9ff;
17'hc22c:	data_out=16'h8a00;
17'hc22d:	data_out=16'ha00;
17'hc22e:	data_out=16'h8503;
17'hc22f:	data_out=16'h89fd;
17'hc230:	data_out=16'h9fe;
17'hc231:	data_out=16'h8a00;
17'hc232:	data_out=16'h9ff;
17'hc233:	data_out=16'h8a00;
17'hc234:	data_out=16'h2cf;
17'hc235:	data_out=16'h8a00;
17'hc236:	data_out=16'h8a00;
17'hc237:	data_out=16'h8a00;
17'hc238:	data_out=16'h80dd;
17'hc239:	data_out=16'h8a00;
17'hc23a:	data_out=16'ha00;
17'hc23b:	data_out=16'h8456;
17'hc23c:	data_out=16'h8a00;
17'hc23d:	data_out=16'h8a00;
17'hc23e:	data_out=16'h8a00;
17'hc23f:	data_out=16'h8a00;
17'hc240:	data_out=16'ha00;
17'hc241:	data_out=16'h8a00;
17'hc242:	data_out=16'ha00;
17'hc243:	data_out=16'h67b;
17'hc244:	data_out=16'h8a00;
17'hc245:	data_out=16'h8a00;
17'hc246:	data_out=16'h8a00;
17'hc247:	data_out=16'ha00;
17'hc248:	data_out=16'ha00;
17'hc249:	data_out=16'h91d;
17'hc24a:	data_out=16'ha00;
17'hc24b:	data_out=16'ha00;
17'hc24c:	data_out=16'ha00;
17'hc24d:	data_out=16'ha00;
17'hc24e:	data_out=16'h8a00;
17'hc24f:	data_out=16'ha00;
17'hc250:	data_out=16'h89a7;
17'hc251:	data_out=16'h8a00;
17'hc252:	data_out=16'h833d;
17'hc253:	data_out=16'h8a00;
17'hc254:	data_out=16'h8a00;
17'hc255:	data_out=16'h89fe;
17'hc256:	data_out=16'h8a00;
17'hc257:	data_out=16'h8a00;
17'hc258:	data_out=16'h8a00;
17'hc259:	data_out=16'ha00;
17'hc25a:	data_out=16'h8a00;
17'hc25b:	data_out=16'h89ff;
17'hc25c:	data_out=16'h8a00;
17'hc25d:	data_out=16'h89f8;
17'hc25e:	data_out=16'h89ec;
17'hc25f:	data_out=16'h89fe;
17'hc260:	data_out=16'h9e9;
17'hc261:	data_out=16'h8a00;
17'hc262:	data_out=16'h827f;
17'hc263:	data_out=16'h8a00;
17'hc264:	data_out=16'h77c;
17'hc265:	data_out=16'ha00;
17'hc266:	data_out=16'ha00;
17'hc267:	data_out=16'ha00;
17'hc268:	data_out=16'h8a00;
17'hc269:	data_out=16'h8a00;
17'hc26a:	data_out=16'h8a00;
17'hc26b:	data_out=16'h89f2;
17'hc26c:	data_out=16'h8a00;
17'hc26d:	data_out=16'h8a00;
17'hc26e:	data_out=16'h8a00;
17'hc26f:	data_out=16'h9ff;
17'hc270:	data_out=16'h8a00;
17'hc271:	data_out=16'h89f6;
17'hc272:	data_out=16'h89da;
17'hc273:	data_out=16'h8606;
17'hc274:	data_out=16'h9f1;
17'hc275:	data_out=16'h8a00;
17'hc276:	data_out=16'ha00;
17'hc277:	data_out=16'h86f4;
17'hc278:	data_out=16'ha00;
17'hc279:	data_out=16'h8a00;
17'hc27a:	data_out=16'h89fd;
17'hc27b:	data_out=16'h8a00;
17'hc27c:	data_out=16'h8a00;
17'hc27d:	data_out=16'h8a00;
17'hc27e:	data_out=16'ha00;
17'hc27f:	data_out=16'h8a00;
17'hc280:	data_out=16'h9f4;
17'hc281:	data_out=16'h281;
17'hc282:	data_out=16'h8a00;
17'hc283:	data_out=16'h8a00;
17'hc284:	data_out=16'ha00;
17'hc285:	data_out=16'h89fb;
17'hc286:	data_out=16'h89b1;
17'hc287:	data_out=16'h8a00;
17'hc288:	data_out=16'h8a00;
17'hc289:	data_out=16'h26;
17'hc28a:	data_out=16'h128;
17'hc28b:	data_out=16'h899d;
17'hc28c:	data_out=16'h8a00;
17'hc28d:	data_out=16'h8a00;
17'hc28e:	data_out=16'h84e5;
17'hc28f:	data_out=16'h8a00;
17'hc290:	data_out=16'h89e9;
17'hc291:	data_out=16'ha00;
17'hc292:	data_out=16'h8a00;
17'hc293:	data_out=16'h89ff;
17'hc294:	data_out=16'h8a00;
17'hc295:	data_out=16'h8560;
17'hc296:	data_out=16'h8a00;
17'hc297:	data_out=16'h8a00;
17'hc298:	data_out=16'h89a4;
17'hc299:	data_out=16'ha00;
17'hc29a:	data_out=16'h77f;
17'hc29b:	data_out=16'h8a00;
17'hc29c:	data_out=16'h810b;
17'hc29d:	data_out=16'h19;
17'hc29e:	data_out=16'h8a00;
17'hc29f:	data_out=16'h89f6;
17'hc2a0:	data_out=16'h9fe;
17'hc2a1:	data_out=16'h84fa;
17'hc2a2:	data_out=16'ha00;
17'hc2a3:	data_out=16'h8a00;
17'hc2a4:	data_out=16'h8a00;
17'hc2a5:	data_out=16'h15c;
17'hc2a6:	data_out=16'h8a00;
17'hc2a7:	data_out=16'h8139;
17'hc2a8:	data_out=16'h854b;
17'hc2a9:	data_out=16'h8a00;
17'hc2aa:	data_out=16'h8a00;
17'hc2ab:	data_out=16'ha00;
17'hc2ac:	data_out=16'h8a00;
17'hc2ad:	data_out=16'h63e;
17'hc2ae:	data_out=16'h89fd;
17'hc2af:	data_out=16'h840b;
17'hc2b0:	data_out=16'h8a00;
17'hc2b1:	data_out=16'h9ce;
17'hc2b2:	data_out=16'h89f8;
17'hc2b3:	data_out=16'h89fe;
17'hc2b4:	data_out=16'ha00;
17'hc2b5:	data_out=16'h89fa;
17'hc2b6:	data_out=16'h8a00;
17'hc2b7:	data_out=16'h8a00;
17'hc2b8:	data_out=16'ha00;
17'hc2b9:	data_out=16'h89fe;
17'hc2ba:	data_out=16'h52e;
17'hc2bb:	data_out=16'h8a00;
17'hc2bc:	data_out=16'h8a00;
17'hc2bd:	data_out=16'h9fb;
17'hc2be:	data_out=16'h8551;
17'hc2bf:	data_out=16'h89fb;
17'hc2c0:	data_out=16'h429;
17'hc2c1:	data_out=16'h8a00;
17'hc2c2:	data_out=16'h705;
17'hc2c3:	data_out=16'h89ff;
17'hc2c4:	data_out=16'h86f4;
17'hc2c5:	data_out=16'h861f;
17'hc2c6:	data_out=16'h8a00;
17'hc2c7:	data_out=16'h3f;
17'hc2c8:	data_out=16'h8845;
17'hc2c9:	data_out=16'h1;
17'hc2ca:	data_out=16'h89be;
17'hc2cb:	data_out=16'h86ea;
17'hc2cc:	data_out=16'h532;
17'hc2cd:	data_out=16'ha00;
17'hc2ce:	data_out=16'h8a00;
17'hc2cf:	data_out=16'h5d4;
17'hc2d0:	data_out=16'h8872;
17'hc2d1:	data_out=16'h8a00;
17'hc2d2:	data_out=16'h8900;
17'hc2d3:	data_out=16'h89fc;
17'hc2d4:	data_out=16'h7cc;
17'hc2d5:	data_out=16'h8a00;
17'hc2d6:	data_out=16'h86d3;
17'hc2d7:	data_out=16'h8051;
17'hc2d8:	data_out=16'h8a00;
17'hc2d9:	data_out=16'h9c9;
17'hc2da:	data_out=16'h8a00;
17'hc2db:	data_out=16'h82ec;
17'hc2dc:	data_out=16'h8633;
17'hc2dd:	data_out=16'h89fa;
17'hc2de:	data_out=16'h8534;
17'hc2df:	data_out=16'h803a;
17'hc2e0:	data_out=16'h8a00;
17'hc2e1:	data_out=16'h84d0;
17'hc2e2:	data_out=16'h8a00;
17'hc2e3:	data_out=16'h89ff;
17'hc2e4:	data_out=16'ha00;
17'hc2e5:	data_out=16'ha00;
17'hc2e6:	data_out=16'h9fc;
17'hc2e7:	data_out=16'h82ff;
17'hc2e8:	data_out=16'h850f;
17'hc2e9:	data_out=16'h8a00;
17'hc2ea:	data_out=16'h84d6;
17'hc2eb:	data_out=16'h9fe;
17'hc2ec:	data_out=16'h80e0;
17'hc2ed:	data_out=16'h89ff;
17'hc2ee:	data_out=16'h84d7;
17'hc2ef:	data_out=16'h89fd;
17'hc2f0:	data_out=16'h84e3;
17'hc2f1:	data_out=16'h8a00;
17'hc2f2:	data_out=16'h896;
17'hc2f3:	data_out=16'ha00;
17'hc2f4:	data_out=16'h8a00;
17'hc2f5:	data_out=16'h8a00;
17'hc2f6:	data_out=16'ha00;
17'hc2f7:	data_out=16'h89fe;
17'hc2f8:	data_out=16'h8951;
17'hc2f9:	data_out=16'h8a00;
17'hc2fa:	data_out=16'h8a00;
17'hc2fb:	data_out=16'h8554;
17'hc2fc:	data_out=16'h842b;
17'hc2fd:	data_out=16'h895c;
17'hc2fe:	data_out=16'h84fd;
17'hc2ff:	data_out=16'h2;
17'hc300:	data_out=16'ha00;
17'hc301:	data_out=16'h7bb;
17'hc302:	data_out=16'h8a00;
17'hc303:	data_out=16'h8237;
17'hc304:	data_out=16'h70d;
17'hc305:	data_out=16'h32a;
17'hc306:	data_out=16'h8246;
17'hc307:	data_out=16'h88c8;
17'hc308:	data_out=16'h8a00;
17'hc309:	data_out=16'h3b6;
17'hc30a:	data_out=16'h605;
17'hc30b:	data_out=16'h89f6;
17'hc30c:	data_out=16'h8a00;
17'hc30d:	data_out=16'h8a00;
17'hc30e:	data_out=16'h8167;
17'hc30f:	data_out=16'h8a00;
17'hc310:	data_out=16'h825e;
17'hc311:	data_out=16'ha00;
17'hc312:	data_out=16'h88fb;
17'hc313:	data_out=16'h8997;
17'hc314:	data_out=16'h80ab;
17'hc315:	data_out=16'h31e;
17'hc316:	data_out=16'h873f;
17'hc317:	data_out=16'h87f9;
17'hc318:	data_out=16'h8168;
17'hc319:	data_out=16'h706;
17'hc31a:	data_out=16'h24a;
17'hc31b:	data_out=16'h8a00;
17'hc31c:	data_out=16'h975;
17'hc31d:	data_out=16'h9ff;
17'hc31e:	data_out=16'h8250;
17'hc31f:	data_out=16'h2ac;
17'hc320:	data_out=16'ha00;
17'hc321:	data_out=16'h8181;
17'hc322:	data_out=16'h5e9;
17'hc323:	data_out=16'h8553;
17'hc324:	data_out=16'h8551;
17'hc325:	data_out=16'h8332;
17'hc326:	data_out=16'h8a00;
17'hc327:	data_out=16'ha00;
17'hc328:	data_out=16'h81a9;
17'hc329:	data_out=16'h855b;
17'hc32a:	data_out=16'h8a00;
17'hc32b:	data_out=16'ha00;
17'hc32c:	data_out=16'h83f3;
17'hc32d:	data_out=16'h8296;
17'hc32e:	data_out=16'h8a00;
17'hc32f:	data_out=16'h415;
17'hc330:	data_out=16'h8a00;
17'hc331:	data_out=16'h9ff;
17'hc332:	data_out=16'h8a00;
17'hc333:	data_out=16'h40d;
17'hc334:	data_out=16'ha00;
17'hc335:	data_out=16'h879f;
17'hc336:	data_out=16'h8a00;
17'hc337:	data_out=16'h8a00;
17'hc338:	data_out=16'ha00;
17'hc339:	data_out=16'h497;
17'hc33a:	data_out=16'h218;
17'hc33b:	data_out=16'h846b;
17'hc33c:	data_out=16'h8a00;
17'hc33d:	data_out=16'ha00;
17'hc33e:	data_out=16'h81ab;
17'hc33f:	data_out=16'h343;
17'hc340:	data_out=16'h1f;
17'hc341:	data_out=16'h8a00;
17'hc342:	data_out=16'h8a00;
17'hc343:	data_out=16'h8394;
17'hc344:	data_out=16'h811;
17'hc345:	data_out=16'h2d3;
17'hc346:	data_out=16'h8669;
17'hc347:	data_out=16'h8124;
17'hc348:	data_out=16'h8585;
17'hc349:	data_out=16'h8339;
17'hc34a:	data_out=16'h89fe;
17'hc34b:	data_out=16'h8a00;
17'hc34c:	data_out=16'h8556;
17'hc34d:	data_out=16'h672;
17'hc34e:	data_out=16'h8a00;
17'hc34f:	data_out=16'h8336;
17'hc350:	data_out=16'h814c;
17'hc351:	data_out=16'h8a00;
17'hc352:	data_out=16'h8486;
17'hc353:	data_out=16'h3f8;
17'hc354:	data_out=16'ha00;
17'hc355:	data_out=16'h8a00;
17'hc356:	data_out=16'h1b9;
17'hc357:	data_out=16'h407;
17'hc358:	data_out=16'h8a00;
17'hc359:	data_out=16'h389;
17'hc35a:	data_out=16'h8a00;
17'hc35b:	data_out=16'ha00;
17'hc35c:	data_out=16'h5d2;
17'hc35d:	data_out=16'h8623;
17'hc35e:	data_out=16'h231;
17'hc35f:	data_out=16'h129;
17'hc360:	data_out=16'h8a00;
17'hc361:	data_out=16'h9cb;
17'hc362:	data_out=16'h8a00;
17'hc363:	data_out=16'h322;
17'hc364:	data_out=16'ha00;
17'hc365:	data_out=16'h297;
17'hc366:	data_out=16'h55d;
17'hc367:	data_out=16'h8313;
17'hc368:	data_out=16'h818e;
17'hc369:	data_out=16'h8a00;
17'hc36a:	data_out=16'h815c;
17'hc36b:	data_out=16'ha00;
17'hc36c:	data_out=16'h16;
17'hc36d:	data_out=16'h385;
17'hc36e:	data_out=16'h815c;
17'hc36f:	data_out=16'h88e1;
17'hc370:	data_out=16'h8162;
17'hc371:	data_out=16'h8a00;
17'hc372:	data_out=16'h92b;
17'hc373:	data_out=16'ha00;
17'hc374:	data_out=16'h8a00;
17'hc375:	data_out=16'h8a00;
17'hc376:	data_out=16'ha00;
17'hc377:	data_out=16'h84f6;
17'hc378:	data_out=16'h830c;
17'hc379:	data_out=16'h8a00;
17'hc37a:	data_out=16'h45;
17'hc37b:	data_out=16'h81ad;
17'hc37c:	data_out=16'h4a;
17'hc37d:	data_out=16'h80d1;
17'hc37e:	data_out=16'h275;
17'hc37f:	data_out=16'h4ab;
17'hc380:	data_out=16'h646;
17'hc381:	data_out=16'h25b;
17'hc382:	data_out=16'h84a2;
17'hc383:	data_out=16'h2d;
17'hc384:	data_out=16'h361;
17'hc385:	data_out=16'h214;
17'hc386:	data_out=16'h80f8;
17'hc387:	data_out=16'h81ec;
17'hc388:	data_out=16'h8421;
17'hc389:	data_out=16'h1a6;
17'hc38a:	data_out=16'h13f;
17'hc38b:	data_out=16'h84c0;
17'hc38c:	data_out=16'h87fb;
17'hc38d:	data_out=16'h8288;
17'hc38e:	data_out=16'h8088;
17'hc38f:	data_out=16'h83c9;
17'hc390:	data_out=16'h805c;
17'hc391:	data_out=16'h4c8;
17'hc392:	data_out=16'h8423;
17'hc393:	data_out=16'h80da;
17'hc394:	data_out=16'h810b;
17'hc395:	data_out=16'h1f7;
17'hc396:	data_out=16'h8070;
17'hc397:	data_out=16'h82d4;
17'hc398:	data_out=16'h80a8;
17'hc399:	data_out=16'h2cb;
17'hc39a:	data_out=16'h22f;
17'hc39b:	data_out=16'h81cd;
17'hc39c:	data_out=16'h5c3;
17'hc39d:	data_out=16'h29f;
17'hc39e:	data_out=16'h807a;
17'hc39f:	data_out=16'h35;
17'hc3a0:	data_out=16'h7fc;
17'hc3a1:	data_out=16'h809d;
17'hc3a2:	data_out=16'h196;
17'hc3a3:	data_out=16'h81d6;
17'hc3a4:	data_out=16'h81d5;
17'hc3a5:	data_out=16'h8114;
17'hc3a6:	data_out=16'h82d3;
17'hc3a7:	data_out=16'h341;
17'hc3a8:	data_out=16'h80a4;
17'hc3a9:	data_out=16'h8176;
17'hc3aa:	data_out=16'h8637;
17'hc3ab:	data_out=16'ha00;
17'hc3ac:	data_out=16'h8035;
17'hc3ad:	data_out=16'h816c;
17'hc3ae:	data_out=16'h856f;
17'hc3af:	data_out=16'h243;
17'hc3b0:	data_out=16'h8321;
17'hc3b1:	data_out=16'h655;
17'hc3b2:	data_out=16'h829d;
17'hc3b3:	data_out=16'h30;
17'hc3b4:	data_out=16'h6ec;
17'hc3b5:	data_out=16'h81fe;
17'hc3b6:	data_out=16'h8355;
17'hc3b7:	data_out=16'h84a7;
17'hc3b8:	data_out=16'ha00;
17'hc3b9:	data_out=16'h183;
17'hc3ba:	data_out=16'h80d3;
17'hc3bb:	data_out=16'h106;
17'hc3bc:	data_out=16'h8548;
17'hc3bd:	data_out=16'h9ea;
17'hc3be:	data_out=16'h809c;
17'hc3bf:	data_out=16'h25a;
17'hc3c0:	data_out=16'hdf;
17'hc3c1:	data_out=16'h8510;
17'hc3c2:	data_out=16'h8291;
17'hc3c3:	data_out=16'h80f5;
17'hc3c4:	data_out=16'h34b;
17'hc3c5:	data_out=16'h1e8;
17'hc3c6:	data_out=16'h8354;
17'hc3c7:	data_out=16'h8154;
17'hc3c8:	data_out=16'h82a9;
17'hc3c9:	data_out=16'h80cb;
17'hc3ca:	data_out=16'h8303;
17'hc3cb:	data_out=16'h87ca;
17'hc3cc:	data_out=16'h81fe;
17'hc3cd:	data_out=16'h2e0;
17'hc3ce:	data_out=16'h8479;
17'hc3cf:	data_out=16'h81a5;
17'hc3d0:	data_out=16'h50;
17'hc3d1:	data_out=16'h82e6;
17'hc3d2:	data_out=16'h81c2;
17'hc3d3:	data_out=16'h12d;
17'hc3d4:	data_out=16'h406;
17'hc3d5:	data_out=16'h85f7;
17'hc3d6:	data_out=16'h804b;
17'hc3d7:	data_out=16'h3a;
17'hc3d8:	data_out=16'h85c6;
17'hc3d9:	data_out=16'h113;
17'hc3da:	data_out=16'h8423;
17'hc3db:	data_out=16'h2e6;
17'hc3dc:	data_out=16'h240;
17'hc3dd:	data_out=16'h81a3;
17'hc3de:	data_out=16'h100;
17'hc3df:	data_out=16'h8025;
17'hc3e0:	data_out=16'h82df;
17'hc3e1:	data_out=16'h4ac;
17'hc3e2:	data_out=16'h85c9;
17'hc3e3:	data_out=16'h8007;
17'hc3e4:	data_out=16'h916;
17'hc3e5:	data_out=16'h241;
17'hc3e6:	data_out=16'h27c;
17'hc3e7:	data_out=16'h81a2;
17'hc3e8:	data_out=16'h8094;
17'hc3e9:	data_out=16'h8609;
17'hc3ea:	data_out=16'h808f;
17'hc3eb:	data_out=16'h61f;
17'hc3ec:	data_out=16'h80a9;
17'hc3ed:	data_out=16'h13;
17'hc3ee:	data_out=16'h8091;
17'hc3ef:	data_out=16'h80b7;
17'hc3f0:	data_out=16'h8093;
17'hc3f1:	data_out=16'h852d;
17'hc3f2:	data_out=16'h34c;
17'hc3f3:	data_out=16'h5cf;
17'hc3f4:	data_out=16'h8359;
17'hc3f5:	data_out=16'h8368;
17'hc3f6:	data_out=16'h49e;
17'hc3f7:	data_out=16'h8085;
17'hc3f8:	data_out=16'h81;
17'hc3f9:	data_out=16'h873a;
17'hc3fa:	data_out=16'h80c4;
17'hc3fb:	data_out=16'h80a6;
17'hc3fc:	data_out=16'h80fa;
17'hc3fd:	data_out=16'h80b8;
17'hc3fe:	data_out=16'h22d;
17'hc3ff:	data_out=16'h146;
17'hc400:	data_out=16'h802b;
17'hc401:	data_out=16'h3a;
17'hc402:	data_out=16'h8006;
17'hc403:	data_out=16'hf;
17'hc404:	data_out=16'h29;
17'hc405:	data_out=16'h8000;
17'hc406:	data_out=16'h1b;
17'hc407:	data_out=16'h801a;
17'hc408:	data_out=16'h8027;
17'hc409:	data_out=16'h8011;
17'hc40a:	data_out=16'h4;
17'hc40b:	data_out=16'h801b;
17'hc40c:	data_out=16'h8027;
17'hc40d:	data_out=16'h801f;
17'hc40e:	data_out=16'h800c;
17'hc40f:	data_out=16'h8010;
17'hc410:	data_out=16'h8037;
17'hc411:	data_out=16'h8015;
17'hc412:	data_out=16'h803a;
17'hc413:	data_out=16'h8013;
17'hc414:	data_out=16'h8059;
17'hc415:	data_out=16'h8014;
17'hc416:	data_out=16'h800e;
17'hc417:	data_out=16'h8051;
17'hc418:	data_out=16'h11;
17'hc419:	data_out=16'h8048;
17'hc41a:	data_out=16'h2b;
17'hc41b:	data_out=16'h802d;
17'hc41c:	data_out=16'h8026;
17'hc41d:	data_out=16'h8003;
17'hc41e:	data_out=16'h803f;
17'hc41f:	data_out=16'h1a;
17'hc420:	data_out=16'h8003;
17'hc421:	data_out=16'h8009;
17'hc422:	data_out=16'h8049;
17'hc423:	data_out=16'h6f;
17'hc424:	data_out=16'h7a;
17'hc425:	data_out=16'h801e;
17'hc426:	data_out=16'h8026;
17'hc427:	data_out=16'h8017;
17'hc428:	data_out=16'h1;
17'hc429:	data_out=16'h802f;
17'hc42a:	data_out=16'h8025;
17'hc42b:	data_out=16'h8021;
17'hc42c:	data_out=16'h8003;
17'hc42d:	data_out=16'h5;
17'hc42e:	data_out=16'h803e;
17'hc42f:	data_out=16'h1d;
17'hc430:	data_out=16'h8032;
17'hc431:	data_out=16'h8028;
17'hc432:	data_out=16'h8037;
17'hc433:	data_out=16'h805a;
17'hc434:	data_out=16'h8011;
17'hc435:	data_out=16'ha;
17'hc436:	data_out=16'h44;
17'hc437:	data_out=16'h801e;
17'hc438:	data_out=16'h66;
17'hc439:	data_out=16'h8033;
17'hc43a:	data_out=16'h26;
17'hc43b:	data_out=16'h6;
17'hc43c:	data_out=16'h8027;
17'hc43d:	data_out=16'h8002;
17'hc43e:	data_out=16'h8005;
17'hc43f:	data_out=16'h12;
17'hc440:	data_out=16'h5e;
17'hc441:	data_out=16'h8023;
17'hc442:	data_out=16'h15;
17'hc443:	data_out=16'h1c;
17'hc444:	data_out=16'h8005;
17'hc445:	data_out=16'h1e;
17'hc446:	data_out=16'h8047;
17'hc447:	data_out=16'h48;
17'hc448:	data_out=16'h8058;
17'hc449:	data_out=16'h8007;
17'hc44a:	data_out=16'h3;
17'hc44b:	data_out=16'h12;
17'hc44c:	data_out=16'h8000;
17'hc44d:	data_out=16'h8029;
17'hc44e:	data_out=16'h8026;
17'hc44f:	data_out=16'h4;
17'hc450:	data_out=16'h64;
17'hc451:	data_out=16'h8005;
17'hc452:	data_out=16'h61;
17'hc453:	data_out=16'h803a;
17'hc454:	data_out=16'h19;
17'hc455:	data_out=16'h3;
17'hc456:	data_out=16'h8032;
17'hc457:	data_out=16'h10;
17'hc458:	data_out=16'h801d;
17'hc459:	data_out=16'h14;
17'hc45a:	data_out=16'h8027;
17'hc45b:	data_out=16'h47;
17'hc45c:	data_out=16'hd;
17'hc45d:	data_out=16'h801c;
17'hc45e:	data_out=16'h7;
17'hc45f:	data_out=16'h8008;
17'hc460:	data_out=16'h8020;
17'hc461:	data_out=16'h16;
17'hc462:	data_out=16'h8010;
17'hc463:	data_out=16'h8052;
17'hc464:	data_out=16'h8033;
17'hc465:	data_out=16'h8002;
17'hc466:	data_out=16'h804c;
17'hc467:	data_out=16'h804f;
17'hc468:	data_out=16'h2;
17'hc469:	data_out=16'hb;
17'hc46a:	data_out=16'h8005;
17'hc46b:	data_out=16'h8012;
17'hc46c:	data_out=16'h0;
17'hc46d:	data_out=16'h8057;
17'hc46e:	data_out=16'h800b;
17'hc46f:	data_out=16'h8016;
17'hc470:	data_out=16'h800c;
17'hc471:	data_out=16'h801d;
17'hc472:	data_out=16'h803d;
17'hc473:	data_out=16'h8001;
17'hc474:	data_out=16'h803b;
17'hc475:	data_out=16'h8011;
17'hc476:	data_out=16'h8039;
17'hc477:	data_out=16'h29;
17'hc478:	data_out=16'h801a;
17'hc479:	data_out=16'h8016;
17'hc47a:	data_out=16'h805a;
17'hc47b:	data_out=16'h800b;
17'hc47c:	data_out=16'he;
17'hc47d:	data_out=16'h28;
17'hc47e:	data_out=16'h8024;
17'hc47f:	data_out=16'h7;
17'hc480:	data_out=16'h807c;
17'hc481:	data_out=16'h10a;
17'hc482:	data_out=16'h66;
17'hc483:	data_out=16'h806f;
17'hc484:	data_out=16'h82f0;
17'hc485:	data_out=16'h81b6;
17'hc486:	data_out=16'h823d;
17'hc487:	data_out=16'h81de;
17'hc488:	data_out=16'h8005;
17'hc489:	data_out=16'h81f0;
17'hc48a:	data_out=16'h80d7;
17'hc48b:	data_out=16'h1c;
17'hc48c:	data_out=16'h813d;
17'hc48d:	data_out=16'h8012;
17'hc48e:	data_out=16'h807c;
17'hc48f:	data_out=16'h804a;
17'hc490:	data_out=16'h8062;
17'hc491:	data_out=16'h829c;
17'hc492:	data_out=16'h136;
17'hc493:	data_out=16'h814d;
17'hc494:	data_out=16'h17a;
17'hc495:	data_out=16'h8180;
17'hc496:	data_out=16'h81d3;
17'hc497:	data_out=16'h224;
17'hc498:	data_out=16'h80b3;
17'hc499:	data_out=16'h8112;
17'hc49a:	data_out=16'h8311;
17'hc49b:	data_out=16'h282;
17'hc49c:	data_out=16'h810e;
17'hc49d:	data_out=16'hf9;
17'hc49e:	data_out=16'h1a9;
17'hc49f:	data_out=16'h82d9;
17'hc4a0:	data_out=16'h213;
17'hc4a1:	data_out=16'h807f;
17'hc4a2:	data_out=16'h92;
17'hc4a3:	data_out=16'h8157;
17'hc4a4:	data_out=16'h8166;
17'hc4a5:	data_out=16'h818f;
17'hc4a6:	data_out=16'h81c1;
17'hc4a7:	data_out=16'h158;
17'hc4a8:	data_out=16'h8082;
17'hc4a9:	data_out=16'h41;
17'hc4aa:	data_out=16'h7a;
17'hc4ab:	data_out=16'h13;
17'hc4ac:	data_out=16'h8197;
17'hc4ad:	data_out=16'hd8;
17'hc4ae:	data_out=16'h95;
17'hc4af:	data_out=16'h249;
17'hc4b0:	data_out=16'h8300;
17'hc4b1:	data_out=16'h80be;
17'hc4b2:	data_out=16'h830c;
17'hc4b3:	data_out=16'h171;
17'hc4b4:	data_out=16'h80a7;
17'hc4b5:	data_out=16'h827a;
17'hc4b6:	data_out=16'h192;
17'hc4b7:	data_out=16'h98;
17'hc4b8:	data_out=16'h81ba;
17'hc4b9:	data_out=16'h6b;
17'hc4ba:	data_out=16'h800e;
17'hc4bb:	data_out=16'h8266;
17'hc4bc:	data_out=16'h1b3;
17'hc4bd:	data_out=16'h8252;
17'hc4be:	data_out=16'h8083;
17'hc4bf:	data_out=16'h8258;
17'hc4c0:	data_out=16'h82f4;
17'hc4c1:	data_out=16'h172;
17'hc4c2:	data_out=16'ha1;
17'hc4c3:	data_out=16'h8269;
17'hc4c4:	data_out=16'h8268;
17'hc4c5:	data_out=16'h81e5;
17'hc4c6:	data_out=16'h194;
17'hc4c7:	data_out=16'h812e;
17'hc4c8:	data_out=16'ha6;
17'hc4c9:	data_out=16'h81cc;
17'hc4ca:	data_out=16'h8119;
17'hc4cb:	data_out=16'hc9;
17'hc4cc:	data_out=16'h8092;
17'hc4cd:	data_out=16'hd1;
17'hc4ce:	data_out=16'h20;
17'hc4cf:	data_out=16'h8151;
17'hc4d0:	data_out=16'h82c3;
17'hc4d1:	data_out=16'h81af;
17'hc4d2:	data_out=16'h81a1;
17'hc4d3:	data_out=16'h405;
17'hc4d4:	data_out=16'h1be;
17'hc4d5:	data_out=16'h22;
17'hc4d6:	data_out=16'h81e7;
17'hc4d7:	data_out=16'h8268;
17'hc4d8:	data_out=16'h89;
17'hc4d9:	data_out=16'h831e;
17'hc4da:	data_out=16'h310;
17'hc4db:	data_out=16'h82a0;
17'hc4dc:	data_out=16'hca;
17'hc4dd:	data_out=16'h9e;
17'hc4de:	data_out=16'h1dc;
17'hc4df:	data_out=16'h9d;
17'hc4e0:	data_out=16'h81d3;
17'hc4e1:	data_out=16'h8306;
17'hc4e2:	data_out=16'hf5;
17'hc4e3:	data_out=16'h17b;
17'hc4e4:	data_out=16'h8195;
17'hc4e5:	data_out=16'h8176;
17'hc4e6:	data_out=16'h8134;
17'hc4e7:	data_out=16'h16;
17'hc4e8:	data_out=16'h8081;
17'hc4e9:	data_out=16'h36;
17'hc4ea:	data_out=16'h8087;
17'hc4eb:	data_out=16'h82f8;
17'hc4ec:	data_out=16'h21c;
17'hc4ed:	data_out=16'h17c;
17'hc4ee:	data_out=16'h8083;
17'hc4ef:	data_out=16'h8157;
17'hc4f0:	data_out=16'h8082;
17'hc4f1:	data_out=16'h8028;
17'hc4f2:	data_out=16'h8310;
17'hc4f3:	data_out=16'h8295;
17'hc4f4:	data_out=16'h8302;
17'hc4f5:	data_out=16'h8177;
17'hc4f6:	data_out=16'h8087;
17'hc4f7:	data_out=16'h83bf;
17'hc4f8:	data_out=16'h828d;
17'hc4f9:	data_out=16'h5e;
17'hc4fa:	data_out=16'h195;
17'hc4fb:	data_out=16'h8084;
17'hc4fc:	data_out=16'h8;
17'hc4fd:	data_out=16'h8252;
17'hc4fe:	data_out=16'h8250;
17'hc4ff:	data_out=16'h838f;
17'hc500:	data_out=16'h55e;
17'hc501:	data_out=16'h8f4;
17'hc502:	data_out=16'h261;
17'hc503:	data_out=16'h2ad;
17'hc504:	data_out=16'h869c;
17'hc505:	data_out=16'h837f;
17'hc506:	data_out=16'h8822;
17'hc507:	data_out=16'h81d2;
17'hc508:	data_out=16'h238;
17'hc509:	data_out=16'h82d2;
17'hc50a:	data_out=16'h1d9;
17'hc50b:	data_out=16'h11;
17'hc50c:	data_out=16'h8372;
17'hc50d:	data_out=16'h22c;
17'hc50e:	data_out=16'h8172;
17'hc50f:	data_out=16'h27c;
17'hc510:	data_out=16'h281;
17'hc511:	data_out=16'h85fe;
17'hc512:	data_out=16'h643;
17'hc513:	data_out=16'h800a;
17'hc514:	data_out=16'h34f;
17'hc515:	data_out=16'h820c;
17'hc516:	data_out=16'h813a;
17'hc517:	data_out=16'h56a;
17'hc518:	data_out=16'h80b4;
17'hc519:	data_out=16'h8237;
17'hc51a:	data_out=16'h871a;
17'hc51b:	data_out=16'h9d0;
17'hc51c:	data_out=16'h8371;
17'hc51d:	data_out=16'h71f;
17'hc51e:	data_out=16'h620;
17'hc51f:	data_out=16'h88d6;
17'hc520:	data_out=16'ha00;
17'hc521:	data_out=16'h8172;
17'hc522:	data_out=16'h590;
17'hc523:	data_out=16'h8355;
17'hc524:	data_out=16'h8355;
17'hc525:	data_out=16'h80b9;
17'hc526:	data_out=16'h842d;
17'hc527:	data_out=16'h819;
17'hc528:	data_out=16'h8168;
17'hc529:	data_out=16'h4b0;
17'hc52a:	data_out=16'h60c;
17'hc52b:	data_out=16'hf0;
17'hc52c:	data_out=16'h81dd;
17'hc52d:	data_out=16'h770;
17'hc52e:	data_out=16'h65e;
17'hc52f:	data_out=16'ha00;
17'hc530:	data_out=16'h869a;
17'hc531:	data_out=16'h1af;
17'hc532:	data_out=16'h8665;
17'hc533:	data_out=16'h3b9;
17'hc534:	data_out=16'h61;
17'hc535:	data_out=16'h86fa;
17'hc536:	data_out=16'h712;
17'hc537:	data_out=16'h25f;
17'hc538:	data_out=16'h824c;
17'hc539:	data_out=16'h465;
17'hc53a:	data_out=16'h6af;
17'hc53b:	data_out=16'h85c4;
17'hc53c:	data_out=16'h6dd;
17'hc53d:	data_out=16'h81ba;
17'hc53e:	data_out=16'h816f;
17'hc53f:	data_out=16'h851c;
17'hc540:	data_out=16'h8670;
17'hc541:	data_out=16'h2be;
17'hc542:	data_out=16'h655;
17'hc543:	data_out=16'h89e2;
17'hc544:	data_out=16'h851b;
17'hc545:	data_out=16'h82b7;
17'hc546:	data_out=16'h420;
17'hc547:	data_out=16'h4d;
17'hc548:	data_out=16'h687;
17'hc549:	data_out=16'h818a;
17'hc54a:	data_out=16'h2d;
17'hc54b:	data_out=16'h629;
17'hc54c:	data_out=16'h37f;
17'hc54d:	data_out=16'h679;
17'hc54e:	data_out=16'h5f8;
17'hc54f:	data_out=16'hf0;
17'hc550:	data_out=16'h86c9;
17'hc551:	data_out=16'h86f2;
17'hc552:	data_out=16'h84cb;
17'hc553:	data_out=16'ha00;
17'hc554:	data_out=16'ha00;
17'hc555:	data_out=16'h81c9;
17'hc556:	data_out=16'h8490;
17'hc557:	data_out=16'h845b;
17'hc558:	data_out=16'h800f;
17'hc559:	data_out=16'h84e7;
17'hc55a:	data_out=16'h9e7;
17'hc55b:	data_out=16'h885f;
17'hc55c:	data_out=16'h503;
17'hc55d:	data_out=16'h917;
17'hc55e:	data_out=16'ha00;
17'hc55f:	data_out=16'h523;
17'hc560:	data_out=16'h8350;
17'hc561:	data_out=16'h8743;
17'hc562:	data_out=16'h208;
17'hc563:	data_out=16'h3e5;
17'hc564:	data_out=16'h8255;
17'hc565:	data_out=16'h80bb;
17'hc566:	data_out=16'h8374;
17'hc567:	data_out=16'h2a2;
17'hc568:	data_out=16'h8166;
17'hc569:	data_out=16'h2ee;
17'hc56a:	data_out=16'h8180;
17'hc56b:	data_out=16'h8667;
17'hc56c:	data_out=16'ha00;
17'hc56d:	data_out=16'h400;
17'hc56e:	data_out=16'h8174;
17'hc56f:	data_out=16'h808b;
17'hc570:	data_out=16'h8173;
17'hc571:	data_out=16'h111;
17'hc572:	data_out=16'h8620;
17'hc573:	data_out=16'h8508;
17'hc574:	data_out=16'h86ab;
17'hc575:	data_out=16'h866d;
17'hc576:	data_out=16'h8169;
17'hc577:	data_out=16'h8903;
17'hc578:	data_out=16'h89a8;
17'hc579:	data_out=16'h616;
17'hc57a:	data_out=16'h3c8;
17'hc57b:	data_out=16'h8166;
17'hc57c:	data_out=16'he0;
17'hc57d:	data_out=16'h89a9;
17'hc57e:	data_out=16'h8584;
17'hc57f:	data_out=16'h86c3;
17'hc580:	data_out=16'h6d7;
17'hc581:	data_out=16'h9ff;
17'hc582:	data_out=16'h800;
17'hc583:	data_out=16'h504;
17'hc584:	data_out=16'h89fb;
17'hc585:	data_out=16'h89f4;
17'hc586:	data_out=16'h89fa;
17'hc587:	data_out=16'h89fe;
17'hc588:	data_out=16'h870;
17'hc589:	data_out=16'h8170;
17'hc58a:	data_out=16'h8a00;
17'hc58b:	data_out=16'h689;
17'hc58c:	data_out=16'h8a00;
17'hc58d:	data_out=16'h9e7;
17'hc58e:	data_out=16'h826b;
17'hc58f:	data_out=16'h8f5;
17'hc590:	data_out=16'h9eb;
17'hc591:	data_out=16'h89f5;
17'hc592:	data_out=16'ha00;
17'hc593:	data_out=16'h47d;
17'hc594:	data_out=16'h9fe;
17'hc595:	data_out=16'h8694;
17'hc596:	data_out=16'h87c6;
17'hc597:	data_out=16'h9fc;
17'hc598:	data_out=16'h37a;
17'hc599:	data_out=16'h89fd;
17'hc59a:	data_out=16'h89f5;
17'hc59b:	data_out=16'h9ff;
17'hc59c:	data_out=16'h8706;
17'hc59d:	data_out=16'h24c;
17'hc59e:	data_out=16'h9fe;
17'hc59f:	data_out=16'h89f8;
17'hc5a0:	data_out=16'h9ff;
17'hc5a1:	data_out=16'h826a;
17'hc5a2:	data_out=16'h9dd;
17'hc5a3:	data_out=16'h8a00;
17'hc5a4:	data_out=16'h8a00;
17'hc5a5:	data_out=16'h8291;
17'hc5a6:	data_out=16'h8a00;
17'hc5a7:	data_out=16'h77c;
17'hc5a8:	data_out=16'h8277;
17'hc5a9:	data_out=16'h9a2;
17'hc5aa:	data_out=16'h9f4;
17'hc5ab:	data_out=16'h21;
17'hc5ac:	data_out=16'h890f;
17'hc5ad:	data_out=16'h9fe;
17'hc5ae:	data_out=16'h9d8;
17'hc5af:	data_out=16'ha00;
17'hc5b0:	data_out=16'h89fc;
17'hc5b1:	data_out=16'h89fa;
17'hc5b2:	data_out=16'h8a00;
17'hc5b3:	data_out=16'ha00;
17'hc5b4:	data_out=16'h832f;
17'hc5b5:	data_out=16'h89ff;
17'hc5b6:	data_out=16'h9ff;
17'hc5b7:	data_out=16'h7e2;
17'hc5b8:	data_out=16'h82fa;
17'hc5b9:	data_out=16'ha00;
17'hc5ba:	data_out=16'h8f3;
17'hc5bb:	data_out=16'h8a00;
17'hc5bc:	data_out=16'h9fb;
17'hc5bd:	data_out=16'h86fa;
17'hc5be:	data_out=16'h8279;
17'hc5bf:	data_out=16'h89f4;
17'hc5c0:	data_out=16'h89fe;
17'hc5c1:	data_out=16'h9f5;
17'hc5c2:	data_out=16'h318;
17'hc5c3:	data_out=16'h89fd;
17'hc5c4:	data_out=16'h89f3;
17'hc5c5:	data_out=16'h86d0;
17'hc5c6:	data_out=16'h975;
17'hc5c7:	data_out=16'h8548;
17'hc5c8:	data_out=16'ha00;
17'hc5c9:	data_out=16'h8504;
17'hc5ca:	data_out=16'h8657;
17'hc5cb:	data_out=16'h857d;
17'hc5cc:	data_out=16'h11c;
17'hc5cd:	data_out=16'h9ff;
17'hc5ce:	data_out=16'ha00;
17'hc5cf:	data_out=16'h83c0;
17'hc5d0:	data_out=16'h893d;
17'hc5d1:	data_out=16'h870d;
17'hc5d2:	data_out=16'h8a00;
17'hc5d3:	data_out=16'h9ff;
17'hc5d4:	data_out=16'ha00;
17'hc5d5:	data_out=16'h9f6;
17'hc5d6:	data_out=16'h8961;
17'hc5d7:	data_out=16'h87c8;
17'hc5d8:	data_out=16'h9fb;
17'hc5d9:	data_out=16'h89fe;
17'hc5da:	data_out=16'ha00;
17'hc5db:	data_out=16'h89f4;
17'hc5dc:	data_out=16'h763;
17'hc5dd:	data_out=16'h9ff;
17'hc5de:	data_out=16'ha00;
17'hc5df:	data_out=16'ha00;
17'hc5e0:	data_out=16'h8a00;
17'hc5e1:	data_out=16'h89fb;
17'hc5e2:	data_out=16'h9f8;
17'hc5e3:	data_out=16'ha00;
17'hc5e4:	data_out=16'h8492;
17'hc5e5:	data_out=16'h89fc;
17'hc5e6:	data_out=16'h89fb;
17'hc5e7:	data_out=16'h205;
17'hc5e8:	data_out=16'h826e;
17'hc5e9:	data_out=16'h59d;
17'hc5ea:	data_out=16'h826d;
17'hc5eb:	data_out=16'h89f2;
17'hc5ec:	data_out=16'h9fd;
17'hc5ed:	data_out=16'ha00;
17'hc5ee:	data_out=16'h826d;
17'hc5ef:	data_out=16'h89fb;
17'hc5f0:	data_out=16'h826c;
17'hc5f1:	data_out=16'h112;
17'hc5f2:	data_out=16'h89fd;
17'hc5f3:	data_out=16'h89fd;
17'hc5f4:	data_out=16'h89f9;
17'hc5f5:	data_out=16'h89e6;
17'hc5f6:	data_out=16'h897f;
17'hc5f7:	data_out=16'h886c;
17'hc5f8:	data_out=16'h89fa;
17'hc5f9:	data_out=16'h9f7;
17'hc5fa:	data_out=16'ha00;
17'hc5fb:	data_out=16'h8279;
17'hc5fc:	data_out=16'h553;
17'hc5fd:	data_out=16'h89f0;
17'hc5fe:	data_out=16'h83c6;
17'hc5ff:	data_out=16'h89a2;
17'hc600:	data_out=16'h89d3;
17'hc601:	data_out=16'h89fc;
17'hc602:	data_out=16'h9f7;
17'hc603:	data_out=16'h530;
17'hc604:	data_out=16'h8a00;
17'hc605:	data_out=16'h8a00;
17'hc606:	data_out=16'h86d3;
17'hc607:	data_out=16'h85d1;
17'hc608:	data_out=16'ha00;
17'hc609:	data_out=16'h9cb;
17'hc60a:	data_out=16'h8a00;
17'hc60b:	data_out=16'ha00;
17'hc60c:	data_out=16'h2d9;
17'hc60d:	data_out=16'h9fa;
17'hc60e:	data_out=16'hbc;
17'hc60f:	data_out=16'h9f3;
17'hc610:	data_out=16'h976;
17'hc611:	data_out=16'h89fd;
17'hc612:	data_out=16'ha00;
17'hc613:	data_out=16'ha00;
17'hc614:	data_out=16'h9fb;
17'hc615:	data_out=16'h8a00;
17'hc616:	data_out=16'h8a00;
17'hc617:	data_out=16'h9fd;
17'hc618:	data_out=16'ha00;
17'hc619:	data_out=16'h89d0;
17'hc61a:	data_out=16'h8a00;
17'hc61b:	data_out=16'ha00;
17'hc61c:	data_out=16'h8799;
17'hc61d:	data_out=16'h89f9;
17'hc61e:	data_out=16'h9fa;
17'hc61f:	data_out=16'h2aa;
17'hc620:	data_out=16'h89f6;
17'hc621:	data_out=16'hf2;
17'hc622:	data_out=16'h7b6;
17'hc623:	data_out=16'h80ef;
17'hc624:	data_out=16'h80ed;
17'hc625:	data_out=16'h5ba;
17'hc626:	data_out=16'h9fe;
17'hc627:	data_out=16'h89f3;
17'hc628:	data_out=16'h144;
17'hc629:	data_out=16'h9fc;
17'hc62a:	data_out=16'h98b;
17'hc62b:	data_out=16'h9ff;
17'hc62c:	data_out=16'h8a00;
17'hc62d:	data_out=16'h2d;
17'hc62e:	data_out=16'h934;
17'hc62f:	data_out=16'h89f5;
17'hc630:	data_out=16'h89fc;
17'hc631:	data_out=16'h8a00;
17'hc632:	data_out=16'h8a00;
17'hc633:	data_out=16'h9ff;
17'hc634:	data_out=16'h89f6;
17'hc635:	data_out=16'h8a00;
17'hc636:	data_out=16'ha00;
17'hc637:	data_out=16'h9f2;
17'hc638:	data_out=16'h89f9;
17'hc639:	data_out=16'ha00;
17'hc63a:	data_out=16'h8ea;
17'hc63b:	data_out=16'h89fb;
17'hc63c:	data_out=16'h9ea;
17'hc63d:	data_out=16'h89fc;
17'hc63e:	data_out=16'h146;
17'hc63f:	data_out=16'h8a00;
17'hc640:	data_out=16'h8a00;
17'hc641:	data_out=16'h9fc;
17'hc642:	data_out=16'h4b9;
17'hc643:	data_out=16'h8449;
17'hc644:	data_out=16'h89fe;
17'hc645:	data_out=16'h8a00;
17'hc646:	data_out=16'h9f2;
17'hc647:	data_out=16'h9ed;
17'hc648:	data_out=16'h9f5;
17'hc649:	data_out=16'h2b2;
17'hc64a:	data_out=16'h89eb;
17'hc64b:	data_out=16'h27b;
17'hc64c:	data_out=16'h262;
17'hc64d:	data_out=16'h949;
17'hc64e:	data_out=16'ha00;
17'hc64f:	data_out=16'h309;
17'hc650:	data_out=16'h8a00;
17'hc651:	data_out=16'h9ed;
17'hc652:	data_out=16'h82ec;
17'hc653:	data_out=16'h8267;
17'hc654:	data_out=16'h89ed;
17'hc655:	data_out=16'h9f0;
17'hc656:	data_out=16'h682;
17'hc657:	data_out=16'h315;
17'hc658:	data_out=16'h9fa;
17'hc659:	data_out=16'h8a00;
17'hc65a:	data_out=16'ha00;
17'hc65b:	data_out=16'h8a00;
17'hc65c:	data_out=16'h89cc;
17'hc65d:	data_out=16'h89fc;
17'hc65e:	data_out=16'h89f6;
17'hc65f:	data_out=16'h3f9;
17'hc660:	data_out=16'ha00;
17'hc661:	data_out=16'h8a00;
17'hc662:	data_out=16'h9f9;
17'hc663:	data_out=16'h9ff;
17'hc664:	data_out=16'h8807;
17'hc665:	data_out=16'h8a00;
17'hc666:	data_out=16'h8990;
17'hc667:	data_out=16'h89b;
17'hc668:	data_out=16'h11d;
17'hc669:	data_out=16'ha00;
17'hc66a:	data_out=16'h9a;
17'hc66b:	data_out=16'h8a00;
17'hc66c:	data_out=16'h89ea;
17'hc66d:	data_out=16'h9ff;
17'hc66e:	data_out=16'h9a;
17'hc66f:	data_out=16'h8a00;
17'hc670:	data_out=16'hac;
17'hc671:	data_out=16'h9ea;
17'hc672:	data_out=16'h8a00;
17'hc673:	data_out=16'h8a00;
17'hc674:	data_out=16'h89f8;
17'hc675:	data_out=16'h8a00;
17'hc676:	data_out=16'h8665;
17'hc677:	data_out=16'h571;
17'hc678:	data_out=16'h8a00;
17'hc679:	data_out=16'ha00;
17'hc67a:	data_out=16'h9fd;
17'hc67b:	data_out=16'h147;
17'hc67c:	data_out=16'h4db;
17'hc67d:	data_out=16'h89ff;
17'hc67e:	data_out=16'h897;
17'hc67f:	data_out=16'h8a00;
17'hc680:	data_out=16'h8a00;
17'hc681:	data_out=16'h8a00;
17'hc682:	data_out=16'h89e5;
17'hc683:	data_out=16'h8198;
17'hc684:	data_out=16'h8a00;
17'hc685:	data_out=16'h8a00;
17'hc686:	data_out=16'h77a;
17'hc687:	data_out=16'ha00;
17'hc688:	data_out=16'h959;
17'hc689:	data_out=16'h9fe;
17'hc68a:	data_out=16'h8a00;
17'hc68b:	data_out=16'ha00;
17'hc68c:	data_out=16'ha00;
17'hc68d:	data_out=16'h9fa;
17'hc68e:	data_out=16'h8775;
17'hc68f:	data_out=16'h8ad;
17'hc690:	data_out=16'h3c7;
17'hc691:	data_out=16'h8a00;
17'hc692:	data_out=16'h93c;
17'hc693:	data_out=16'h9fd;
17'hc694:	data_out=16'h8669;
17'hc695:	data_out=16'h8a00;
17'hc696:	data_out=16'h8a00;
17'hc697:	data_out=16'h9cb;
17'hc698:	data_out=16'h8597;
17'hc699:	data_out=16'h894f;
17'hc69a:	data_out=16'h8a00;
17'hc69b:	data_out=16'h2ed;
17'hc69c:	data_out=16'h8a00;
17'hc69d:	data_out=16'h8a00;
17'hc69e:	data_out=16'h8a00;
17'hc69f:	data_out=16'h84a4;
17'hc6a0:	data_out=16'h8a00;
17'hc6a1:	data_out=16'h869f;
17'hc6a2:	data_out=16'h305;
17'hc6a3:	data_out=16'ha00;
17'hc6a4:	data_out=16'ha00;
17'hc6a5:	data_out=16'h93a;
17'hc6a6:	data_out=16'ha00;
17'hc6a7:	data_out=16'h8a00;
17'hc6a8:	data_out=16'h8605;
17'hc6a9:	data_out=16'hd1;
17'hc6aa:	data_out=16'h7f7;
17'hc6ab:	data_out=16'h1d6;
17'hc6ac:	data_out=16'h8a00;
17'hc6ad:	data_out=16'ha00;
17'hc6ae:	data_out=16'h7c4;
17'hc6af:	data_out=16'h8a00;
17'hc6b0:	data_out=16'h87de;
17'hc6b1:	data_out=16'h8a00;
17'hc6b2:	data_out=16'h89f3;
17'hc6b3:	data_out=16'h8a00;
17'hc6b4:	data_out=16'h8a00;
17'hc6b5:	data_out=16'h8a00;
17'hc6b6:	data_out=16'h8a00;
17'hc6b7:	data_out=16'h803c;
17'hc6b8:	data_out=16'h8a00;
17'hc6b9:	data_out=16'h8a00;
17'hc6ba:	data_out=16'h9e2;
17'hc6bb:	data_out=16'h86d2;
17'hc6bc:	data_out=16'h87c6;
17'hc6bd:	data_out=16'h8a00;
17'hc6be:	data_out=16'h8602;
17'hc6bf:	data_out=16'h8a00;
17'hc6c0:	data_out=16'h8a00;
17'hc6c1:	data_out=16'h9a8;
17'hc6c2:	data_out=16'ha00;
17'hc6c3:	data_out=16'h8139;
17'hc6c4:	data_out=16'h8a00;
17'hc6c5:	data_out=16'h8a00;
17'hc6c6:	data_out=16'h838c;
17'hc6c7:	data_out=16'h9f0;
17'hc6c8:	data_out=16'h31d;
17'hc6c9:	data_out=16'h9da;
17'hc6ca:	data_out=16'h967;
17'hc6cb:	data_out=16'ha00;
17'hc6cc:	data_out=16'h9ef;
17'hc6cd:	data_out=16'h25d;
17'hc6ce:	data_out=16'hb1;
17'hc6cf:	data_out=16'ha00;
17'hc6d0:	data_out=16'h8a00;
17'hc6d1:	data_out=16'h97f;
17'hc6d2:	data_out=16'ha00;
17'hc6d3:	data_out=16'h8a00;
17'hc6d4:	data_out=16'h8a00;
17'hc6d5:	data_out=16'h9d3;
17'hc6d6:	data_out=16'h89ef;
17'hc6d7:	data_out=16'h8a00;
17'hc6d8:	data_out=16'h817;
17'hc6d9:	data_out=16'h8a00;
17'hc6da:	data_out=16'h4e9;
17'hc6db:	data_out=16'h8a00;
17'hc6dc:	data_out=16'h8a00;
17'hc6dd:	data_out=16'h8a00;
17'hc6de:	data_out=16'h8a00;
17'hc6df:	data_out=16'h8a00;
17'hc6e0:	data_out=16'ha00;
17'hc6e1:	data_out=16'h8a00;
17'hc6e2:	data_out=16'h9e2;
17'hc6e3:	data_out=16'h8a00;
17'hc6e4:	data_out=16'h89fd;
17'hc6e5:	data_out=16'h8a00;
17'hc6e6:	data_out=16'h80e0;
17'hc6e7:	data_out=16'h848a;
17'hc6e8:	data_out=16'h863d;
17'hc6e9:	data_out=16'h9eb;
17'hc6ea:	data_out=16'h884b;
17'hc6eb:	data_out=16'h8a00;
17'hc6ec:	data_out=16'h8a00;
17'hc6ed:	data_out=16'h8a00;
17'hc6ee:	data_out=16'h8844;
17'hc6ef:	data_out=16'h89ec;
17'hc6f0:	data_out=16'h87c4;
17'hc6f1:	data_out=16'h207;
17'hc6f2:	data_out=16'h8a00;
17'hc6f3:	data_out=16'h8a00;
17'hc6f4:	data_out=16'h8714;
17'hc6f5:	data_out=16'h8a00;
17'hc6f6:	data_out=16'h6c3;
17'hc6f7:	data_out=16'h9f6;
17'hc6f8:	data_out=16'h8a00;
17'hc6f9:	data_out=16'h40f;
17'hc6fa:	data_out=16'h8a00;
17'hc6fb:	data_out=16'h85fd;
17'hc6fc:	data_out=16'h8a00;
17'hc6fd:	data_out=16'h8a00;
17'hc6fe:	data_out=16'h721;
17'hc6ff:	data_out=16'h8a00;
17'hc700:	data_out=16'h8a00;
17'hc701:	data_out=16'h8a00;
17'hc702:	data_out=16'h89d4;
17'hc703:	data_out=16'h6ee;
17'hc704:	data_out=16'h8a00;
17'hc705:	data_out=16'h8a00;
17'hc706:	data_out=16'h9c1;
17'hc707:	data_out=16'ha00;
17'hc708:	data_out=16'h855d;
17'hc709:	data_out=16'ha00;
17'hc70a:	data_out=16'h8a00;
17'hc70b:	data_out=16'ha00;
17'hc70c:	data_out=16'ha00;
17'hc70d:	data_out=16'h9f0;
17'hc70e:	data_out=16'h8a00;
17'hc70f:	data_out=16'h98c;
17'hc710:	data_out=16'h3a2;
17'hc711:	data_out=16'h8a00;
17'hc712:	data_out=16'h70a;
17'hc713:	data_out=16'ha00;
17'hc714:	data_out=16'h414;
17'hc715:	data_out=16'h8a00;
17'hc716:	data_out=16'h89ff;
17'hc717:	data_out=16'h9ca;
17'hc718:	data_out=16'h8507;
17'hc719:	data_out=16'ha00;
17'hc71a:	data_out=16'h8a00;
17'hc71b:	data_out=16'h93b;
17'hc71c:	data_out=16'h8a00;
17'hc71d:	data_out=16'h8a00;
17'hc71e:	data_out=16'h89fe;
17'hc71f:	data_out=16'h745;
17'hc720:	data_out=16'h8a00;
17'hc721:	data_out=16'h8a00;
17'hc722:	data_out=16'h343;
17'hc723:	data_out=16'ha00;
17'hc724:	data_out=16'ha00;
17'hc725:	data_out=16'h9f0;
17'hc726:	data_out=16'ha00;
17'hc727:	data_out=16'h8a00;
17'hc728:	data_out=16'h8a00;
17'hc729:	data_out=16'h8299;
17'hc72a:	data_out=16'h4ab;
17'hc72b:	data_out=16'h803b;
17'hc72c:	data_out=16'h89ff;
17'hc72d:	data_out=16'ha00;
17'hc72e:	data_out=16'h8163;
17'hc72f:	data_out=16'h8a00;
17'hc730:	data_out=16'h839d;
17'hc731:	data_out=16'h8a00;
17'hc732:	data_out=16'h8a00;
17'hc733:	data_out=16'h89ff;
17'hc734:	data_out=16'h8a00;
17'hc735:	data_out=16'h89fd;
17'hc736:	data_out=16'h89ff;
17'hc737:	data_out=16'h83b4;
17'hc738:	data_out=16'h8a00;
17'hc739:	data_out=16'h8a00;
17'hc73a:	data_out=16'ha00;
17'hc73b:	data_out=16'h204;
17'hc73c:	data_out=16'h8a00;
17'hc73d:	data_out=16'h8a00;
17'hc73e:	data_out=16'h8a00;
17'hc73f:	data_out=16'h8a00;
17'hc740:	data_out=16'h8a00;
17'hc741:	data_out=16'h875c;
17'hc742:	data_out=16'ha00;
17'hc743:	data_out=16'h6d0;
17'hc744:	data_out=16'h8a00;
17'hc745:	data_out=16'h8a00;
17'hc746:	data_out=16'h89d4;
17'hc747:	data_out=16'ha00;
17'hc748:	data_out=16'h8cb;
17'hc749:	data_out=16'h9fe;
17'hc74a:	data_out=16'h249;
17'hc74b:	data_out=16'ha00;
17'hc74c:	data_out=16'h9f3;
17'hc74d:	data_out=16'h8327;
17'hc74e:	data_out=16'h8242;
17'hc74f:	data_out=16'ha00;
17'hc750:	data_out=16'h8a00;
17'hc751:	data_out=16'h9d3;
17'hc752:	data_out=16'ha00;
17'hc753:	data_out=16'h8a00;
17'hc754:	data_out=16'h8a00;
17'hc755:	data_out=16'h9f0;
17'hc756:	data_out=16'h9cf;
17'hc757:	data_out=16'h8a00;
17'hc758:	data_out=16'h89d7;
17'hc759:	data_out=16'h8a00;
17'hc75a:	data_out=16'h13f;
17'hc75b:	data_out=16'h8a00;
17'hc75c:	data_out=16'h8a00;
17'hc75d:	data_out=16'h8a00;
17'hc75e:	data_out=16'h8a00;
17'hc75f:	data_out=16'h8a00;
17'hc760:	data_out=16'ha00;
17'hc761:	data_out=16'h8a00;
17'hc762:	data_out=16'h9e8;
17'hc763:	data_out=16'h89ff;
17'hc764:	data_out=16'h8a00;
17'hc765:	data_out=16'h8a00;
17'hc766:	data_out=16'ha00;
17'hc767:	data_out=16'h9da;
17'hc768:	data_out=16'h8a00;
17'hc769:	data_out=16'h9dd;
17'hc76a:	data_out=16'h8a00;
17'hc76b:	data_out=16'h8a00;
17'hc76c:	data_out=16'h8a00;
17'hc76d:	data_out=16'h89ff;
17'hc76e:	data_out=16'h8a00;
17'hc76f:	data_out=16'h8a00;
17'hc770:	data_out=16'h8a00;
17'hc771:	data_out=16'h308;
17'hc772:	data_out=16'h8a00;
17'hc773:	data_out=16'h8a00;
17'hc774:	data_out=16'h82d3;
17'hc775:	data_out=16'h8a00;
17'hc776:	data_out=16'ha00;
17'hc777:	data_out=16'ha00;
17'hc778:	data_out=16'h8a00;
17'hc779:	data_out=16'h8769;
17'hc77a:	data_out=16'h88f5;
17'hc77b:	data_out=16'h8a00;
17'hc77c:	data_out=16'h8a00;
17'hc77d:	data_out=16'h8a00;
17'hc77e:	data_out=16'h9b4;
17'hc77f:	data_out=16'h8a00;
17'hc780:	data_out=16'h8a00;
17'hc781:	data_out=16'h8a00;
17'hc782:	data_out=16'h85f6;
17'hc783:	data_out=16'h4c5;
17'hc784:	data_out=16'h89fc;
17'hc785:	data_out=16'h8a00;
17'hc786:	data_out=16'h9c2;
17'hc787:	data_out=16'ha00;
17'hc788:	data_out=16'h89fb;
17'hc789:	data_out=16'ha00;
17'hc78a:	data_out=16'h8a00;
17'hc78b:	data_out=16'ha00;
17'hc78c:	data_out=16'ha00;
17'hc78d:	data_out=16'h9dd;
17'hc78e:	data_out=16'h89ff;
17'hc78f:	data_out=16'h9e4;
17'hc790:	data_out=16'h856a;
17'hc791:	data_out=16'h8a00;
17'hc792:	data_out=16'h8a8;
17'hc793:	data_out=16'h9d9;
17'hc794:	data_out=16'h9b9;
17'hc795:	data_out=16'h8a00;
17'hc796:	data_out=16'h88a1;
17'hc797:	data_out=16'h9b7;
17'hc798:	data_out=16'h81a1;
17'hc799:	data_out=16'h320;
17'hc79a:	data_out=16'h8a00;
17'hc79b:	data_out=16'h9f4;
17'hc79c:	data_out=16'h8a00;
17'hc79d:	data_out=16'h8a00;
17'hc79e:	data_out=16'h8569;
17'hc79f:	data_out=16'h918;
17'hc7a0:	data_out=16'h8a00;
17'hc7a1:	data_out=16'h89ff;
17'hc7a2:	data_out=16'h89ff;
17'hc7a3:	data_out=16'ha00;
17'hc7a4:	data_out=16'ha00;
17'hc7a5:	data_out=16'h9e8;
17'hc7a6:	data_out=16'ha00;
17'hc7a7:	data_out=16'h8a00;
17'hc7a8:	data_out=16'h89fb;
17'hc7a9:	data_out=16'h89db;
17'hc7aa:	data_out=16'h787;
17'hc7ab:	data_out=16'hd3;
17'hc7ac:	data_out=16'h89fd;
17'hc7ad:	data_out=16'h9eb;
17'hc7ae:	data_out=16'h308;
17'hc7af:	data_out=16'h8a00;
17'hc7b0:	data_out=16'h8019;
17'hc7b1:	data_out=16'h8a00;
17'hc7b2:	data_out=16'h8a00;
17'hc7b3:	data_out=16'h89f7;
17'hc7b4:	data_out=16'h8a00;
17'hc7b5:	data_out=16'h8132;
17'hc7b6:	data_out=16'h89fc;
17'hc7b7:	data_out=16'h33c;
17'hc7b8:	data_out=16'h8a00;
17'hc7b9:	data_out=16'h89f9;
17'hc7ba:	data_out=16'ha00;
17'hc7bb:	data_out=16'h9ee;
17'hc7bc:	data_out=16'h89ff;
17'hc7bd:	data_out=16'h8a00;
17'hc7be:	data_out=16'h89fa;
17'hc7bf:	data_out=16'h8a00;
17'hc7c0:	data_out=16'h8a00;
17'hc7c1:	data_out=16'h89f2;
17'hc7c2:	data_out=16'ha00;
17'hc7c3:	data_out=16'h83d2;
17'hc7c4:	data_out=16'h8a00;
17'hc7c5:	data_out=16'h8a00;
17'hc7c6:	data_out=16'h8a00;
17'hc7c7:	data_out=16'ha00;
17'hc7c8:	data_out=16'h84f;
17'hc7c9:	data_out=16'h9ff;
17'hc7ca:	data_out=16'h80a2;
17'hc7cb:	data_out=16'ha00;
17'hc7cc:	data_out=16'h9d1;
17'hc7cd:	data_out=16'h8a00;
17'hc7ce:	data_out=16'h87ea;
17'hc7cf:	data_out=16'ha00;
17'hc7d0:	data_out=16'h8a00;
17'hc7d1:	data_out=16'h9d7;
17'hc7d2:	data_out=16'ha00;
17'hc7d3:	data_out=16'h8a00;
17'hc7d4:	data_out=16'h8a00;
17'hc7d5:	data_out=16'ha00;
17'hc7d6:	data_out=16'h9e6;
17'hc7d7:	data_out=16'h7f5;
17'hc7d8:	data_out=16'h89aa;
17'hc7d9:	data_out=16'h8a00;
17'hc7da:	data_out=16'h80c2;
17'hc7db:	data_out=16'h8a00;
17'hc7dc:	data_out=16'h8a00;
17'hc7dd:	data_out=16'h8a00;
17'hc7de:	data_out=16'h8a00;
17'hc7df:	data_out=16'h8a00;
17'hc7e0:	data_out=16'ha00;
17'hc7e1:	data_out=16'h8a00;
17'hc7e2:	data_out=16'h9cc;
17'hc7e3:	data_out=16'h89f9;
17'hc7e4:	data_out=16'h8a00;
17'hc7e5:	data_out=16'h8a00;
17'hc7e6:	data_out=16'ha00;
17'hc7e7:	data_out=16'ha00;
17'hc7e8:	data_out=16'h89e5;
17'hc7e9:	data_out=16'h9de;
17'hc7ea:	data_out=16'h89ff;
17'hc7eb:	data_out=16'h8a00;
17'hc7ec:	data_out=16'h8a00;
17'hc7ed:	data_out=16'h89f9;
17'hc7ee:	data_out=16'h89ff;
17'hc7ef:	data_out=16'h8a00;
17'hc7f0:	data_out=16'h89ff;
17'hc7f1:	data_out=16'h9dd;
17'hc7f2:	data_out=16'h8a00;
17'hc7f3:	data_out=16'h8a00;
17'hc7f4:	data_out=16'h61;
17'hc7f5:	data_out=16'h8a00;
17'hc7f6:	data_out=16'ha00;
17'hc7f7:	data_out=16'h9e2;
17'hc7f8:	data_out=16'h8a00;
17'hc7f9:	data_out=16'h89fb;
17'hc7fa:	data_out=16'h850a;
17'hc7fb:	data_out=16'h89f9;
17'hc7fc:	data_out=16'h8a00;
17'hc7fd:	data_out=16'h83b1;
17'hc7fe:	data_out=16'h9e4;
17'hc7ff:	data_out=16'h8a00;
17'hc800:	data_out=16'h89fe;
17'hc801:	data_out=16'h8a00;
17'hc802:	data_out=16'h9ff;
17'hc803:	data_out=16'h632;
17'hc804:	data_out=16'h89a8;
17'hc805:	data_out=16'h8a00;
17'hc806:	data_out=16'h9a0;
17'hc807:	data_out=16'ha00;
17'hc808:	data_out=16'h89ca;
17'hc809:	data_out=16'ha00;
17'hc80a:	data_out=16'h8995;
17'hc80b:	data_out=16'h9eb;
17'hc80c:	data_out=16'ha00;
17'hc80d:	data_out=16'h9fd;
17'hc80e:	data_out=16'h9ff;
17'hc80f:	data_out=16'h9ff;
17'hc810:	data_out=16'h89f5;
17'hc811:	data_out=16'h8a00;
17'hc812:	data_out=16'h9f3;
17'hc813:	data_out=16'h9c6;
17'hc814:	data_out=16'h9d7;
17'hc815:	data_out=16'h89f5;
17'hc816:	data_out=16'h8232;
17'hc817:	data_out=16'h9d1;
17'hc818:	data_out=16'h6c1;
17'hc819:	data_out=16'h89d7;
17'hc81a:	data_out=16'h8a00;
17'hc81b:	data_out=16'ha00;
17'hc81c:	data_out=16'h89f7;
17'hc81d:	data_out=16'h8a00;
17'hc81e:	data_out=16'h2fd;
17'hc81f:	data_out=16'h9bd;
17'hc820:	data_out=16'h8a00;
17'hc821:	data_out=16'h9ff;
17'hc822:	data_out=16'h8a00;
17'hc823:	data_out=16'ha00;
17'hc824:	data_out=16'ha00;
17'hc825:	data_out=16'h9e8;
17'hc826:	data_out=16'ha00;
17'hc827:	data_out=16'h89c4;
17'hc828:	data_out=16'h9ff;
17'hc829:	data_out=16'h8701;
17'hc82a:	data_out=16'h5cb;
17'hc82b:	data_out=16'h89e4;
17'hc82c:	data_out=16'h8554;
17'hc82d:	data_out=16'h831d;
17'hc82e:	data_out=16'h275;
17'hc82f:	data_out=16'h89fe;
17'hc830:	data_out=16'h992;
17'hc831:	data_out=16'h89d5;
17'hc832:	data_out=16'h89ec;
17'hc833:	data_out=16'h860c;
17'hc834:	data_out=16'h8a00;
17'hc835:	data_out=16'ha00;
17'hc836:	data_out=16'h89d8;
17'hc837:	data_out=16'ha00;
17'hc838:	data_out=16'h8a00;
17'hc839:	data_out=16'h895c;
17'hc83a:	data_out=16'h9ff;
17'hc83b:	data_out=16'ha00;
17'hc83c:	data_out=16'h8a00;
17'hc83d:	data_out=16'h8a00;
17'hc83e:	data_out=16'h9ff;
17'hc83f:	data_out=16'h8a00;
17'hc840:	data_out=16'h89ed;
17'hc841:	data_out=16'h87a5;
17'hc842:	data_out=16'h9ee;
17'hc843:	data_out=16'h859c;
17'hc844:	data_out=16'h898e;
17'hc845:	data_out=16'h89f4;
17'hc846:	data_out=16'h8a00;
17'hc847:	data_out=16'ha00;
17'hc848:	data_out=16'h85b;
17'hc849:	data_out=16'ha00;
17'hc84a:	data_out=16'h8494;
17'hc84b:	data_out=16'h9db;
17'hc84c:	data_out=16'h9ce;
17'hc84d:	data_out=16'h8a00;
17'hc84e:	data_out=16'h86a2;
17'hc84f:	data_out=16'h9fe;
17'hc850:	data_out=16'h89f6;
17'hc851:	data_out=16'ha00;
17'hc852:	data_out=16'ha00;
17'hc853:	data_out=16'h89f1;
17'hc854:	data_out=16'h8a00;
17'hc855:	data_out=16'ha00;
17'hc856:	data_out=16'ha00;
17'hc857:	data_out=16'h9c7;
17'hc858:	data_out=16'h9d3;
17'hc859:	data_out=16'h89f4;
17'hc85a:	data_out=16'h1fe;
17'hc85b:	data_out=16'h89a2;
17'hc85c:	data_out=16'h8a00;
17'hc85d:	data_out=16'h8a00;
17'hc85e:	data_out=16'h89fd;
17'hc85f:	data_out=16'h8a00;
17'hc860:	data_out=16'h9ff;
17'hc861:	data_out=16'h89f3;
17'hc862:	data_out=16'h9ce;
17'hc863:	data_out=16'h8839;
17'hc864:	data_out=16'h8a00;
17'hc865:	data_out=16'h8a00;
17'hc866:	data_out=16'ha00;
17'hc867:	data_out=16'ha00;
17'hc868:	data_out=16'h9ff;
17'hc869:	data_out=16'h9cd;
17'hc86a:	data_out=16'h9ff;
17'hc86b:	data_out=16'h89ff;
17'hc86c:	data_out=16'h8a00;
17'hc86d:	data_out=16'h886d;
17'hc86e:	data_out=16'h9ff;
17'hc86f:	data_out=16'h89f8;
17'hc870:	data_out=16'h9ff;
17'hc871:	data_out=16'h9fa;
17'hc872:	data_out=16'h8a00;
17'hc873:	data_out=16'h8a00;
17'hc874:	data_out=16'ha00;
17'hc875:	data_out=16'h8a00;
17'hc876:	data_out=16'ha00;
17'hc877:	data_out=16'h9cb;
17'hc878:	data_out=16'h8a00;
17'hc879:	data_out=16'h89a7;
17'hc87a:	data_out=16'h159;
17'hc87b:	data_out=16'h9ff;
17'hc87c:	data_out=16'h89f1;
17'hc87d:	data_out=16'h8e2;
17'hc87e:	data_out=16'h9c9;
17'hc87f:	data_out=16'h8a00;
17'hc880:	data_out=16'h8a00;
17'hc881:	data_out=16'h8a00;
17'hc882:	data_out=16'ha00;
17'hc883:	data_out=16'hd6;
17'hc884:	data_out=16'h88c0;
17'hc885:	data_out=16'h8946;
17'hc886:	data_out=16'h9af;
17'hc887:	data_out=16'ha00;
17'hc888:	data_out=16'h86b3;
17'hc889:	data_out=16'ha00;
17'hc88a:	data_out=16'h897a;
17'hc88b:	data_out=16'h9e8;
17'hc88c:	data_out=16'ha00;
17'hc88d:	data_out=16'ha00;
17'hc88e:	data_out=16'ha00;
17'hc88f:	data_out=16'h9ff;
17'hc890:	data_out=16'h89f5;
17'hc891:	data_out=16'h89ee;
17'hc892:	data_out=16'h816b;
17'hc893:	data_out=16'h5cf;
17'hc894:	data_out=16'h9ff;
17'hc895:	data_out=16'h89b7;
17'hc896:	data_out=16'h807e;
17'hc897:	data_out=16'h658;
17'hc898:	data_out=16'h9ff;
17'hc899:	data_out=16'h89ff;
17'hc89a:	data_out=16'h8981;
17'hc89b:	data_out=16'ha00;
17'hc89c:	data_out=16'h89cf;
17'hc89d:	data_out=16'h8a00;
17'hc89e:	data_out=16'h236;
17'hc89f:	data_out=16'h9e9;
17'hc8a0:	data_out=16'h89f6;
17'hc8a1:	data_out=16'ha00;
17'hc8a2:	data_out=16'h8a00;
17'hc8a3:	data_out=16'ha00;
17'hc8a4:	data_out=16'ha00;
17'hc8a5:	data_out=16'ha00;
17'hc8a6:	data_out=16'ha00;
17'hc8a7:	data_out=16'h8951;
17'hc8a8:	data_out=16'ha00;
17'hc8a9:	data_out=16'h8a00;
17'hc8aa:	data_out=16'h8267;
17'hc8ab:	data_out=16'h89f9;
17'hc8ac:	data_out=16'h8464;
17'hc8ad:	data_out=16'h8a00;
17'hc8ae:	data_out=16'h82cc;
17'hc8af:	data_out=16'h89c4;
17'hc8b0:	data_out=16'ha00;
17'hc8b1:	data_out=16'h896c;
17'hc8b2:	data_out=16'h8941;
17'hc8b3:	data_out=16'h8595;
17'hc8b4:	data_out=16'h8a00;
17'hc8b5:	data_out=16'ha00;
17'hc8b6:	data_out=16'h8976;
17'hc8b7:	data_out=16'ha00;
17'hc8b8:	data_out=16'h8a00;
17'hc8b9:	data_out=16'h88f4;
17'hc8ba:	data_out=16'h9f2;
17'hc8bb:	data_out=16'ha00;
17'hc8bc:	data_out=16'h89f1;
17'hc8bd:	data_out=16'h89bc;
17'hc8be:	data_out=16'ha00;
17'hc8bf:	data_out=16'h8946;
17'hc8c0:	data_out=16'h894f;
17'hc8c1:	data_out=16'h609;
17'hc8c2:	data_out=16'h9cb;
17'hc8c3:	data_out=16'h846e;
17'hc8c4:	data_out=16'h6b1;
17'hc8c5:	data_out=16'h89ae;
17'hc8c6:	data_out=16'h8a00;
17'hc8c7:	data_out=16'h9c6;
17'hc8c8:	data_out=16'h8870;
17'hc8c9:	data_out=16'ha00;
17'hc8ca:	data_out=16'h82e2;
17'hc8cb:	data_out=16'h9b6;
17'hc8cc:	data_out=16'h9ce;
17'hc8cd:	data_out=16'h8a00;
17'hc8ce:	data_out=16'h8983;
17'hc8cf:	data_out=16'h9e1;
17'hc8d0:	data_out=16'h89bd;
17'hc8d1:	data_out=16'ha00;
17'hc8d2:	data_out=16'ha00;
17'hc8d3:	data_out=16'h898c;
17'hc8d4:	data_out=16'h89f3;
17'hc8d5:	data_out=16'ha00;
17'hc8d6:	data_out=16'ha00;
17'hc8d7:	data_out=16'h9ce;
17'hc8d8:	data_out=16'ha00;
17'hc8d9:	data_out=16'h89b7;
17'hc8da:	data_out=16'h1a2;
17'hc8db:	data_out=16'h88ea;
17'hc8dc:	data_out=16'h89a8;
17'hc8dd:	data_out=16'h89ba;
17'hc8de:	data_out=16'h898b;
17'hc8df:	data_out=16'h8a00;
17'hc8e0:	data_out=16'h9f4;
17'hc8e1:	data_out=16'h8934;
17'hc8e2:	data_out=16'h79d;
17'hc8e3:	data_out=16'h87ce;
17'hc8e4:	data_out=16'h8a00;
17'hc8e5:	data_out=16'h8a00;
17'hc8e6:	data_out=16'ha00;
17'hc8e7:	data_out=16'h9e6;
17'hc8e8:	data_out=16'ha00;
17'hc8e9:	data_out=16'h9b9;
17'hc8ea:	data_out=16'ha00;
17'hc8eb:	data_out=16'h8975;
17'hc8ec:	data_out=16'h8a00;
17'hc8ed:	data_out=16'h8811;
17'hc8ee:	data_out=16'ha00;
17'hc8ef:	data_out=16'h8962;
17'hc8f0:	data_out=16'ha00;
17'hc8f1:	data_out=16'h9fb;
17'hc8f2:	data_out=16'h89fa;
17'hc8f3:	data_out=16'h89dc;
17'hc8f4:	data_out=16'ha00;
17'hc8f5:	data_out=16'h89a3;
17'hc8f6:	data_out=16'ha00;
17'hc8f7:	data_out=16'h9f7;
17'hc8f8:	data_out=16'h8a00;
17'hc8f9:	data_out=16'h81a5;
17'hc8fa:	data_out=16'h8b;
17'hc8fb:	data_out=16'ha00;
17'hc8fc:	data_out=16'h89de;
17'hc8fd:	data_out=16'h9ff;
17'hc8fe:	data_out=16'h9de;
17'hc8ff:	data_out=16'h8a00;
17'hc900:	data_out=16'h8a00;
17'hc901:	data_out=16'h8a00;
17'hc902:	data_out=16'ha00;
17'hc903:	data_out=16'h88c0;
17'hc904:	data_out=16'h865a;
17'hc905:	data_out=16'h894d;
17'hc906:	data_out=16'h9b1;
17'hc907:	data_out=16'ha00;
17'hc908:	data_out=16'h830b;
17'hc909:	data_out=16'ha00;
17'hc90a:	data_out=16'h8a00;
17'hc90b:	data_out=16'h982;
17'hc90c:	data_out=16'ha00;
17'hc90d:	data_out=16'h622;
17'hc90e:	data_out=16'ha00;
17'hc90f:	data_out=16'h9fb;
17'hc910:	data_out=16'h89e8;
17'hc911:	data_out=16'h87b7;
17'hc912:	data_out=16'h874f;
17'hc913:	data_out=16'h89bb;
17'hc914:	data_out=16'h8873;
17'hc915:	data_out=16'h895e;
17'hc916:	data_out=16'h886e;
17'hc917:	data_out=16'h8939;
17'hc918:	data_out=16'h9fd;
17'hc919:	data_out=16'h8a00;
17'hc91a:	data_out=16'h89c5;
17'hc91b:	data_out=16'h3bd;
17'hc91c:	data_out=16'h89c5;
17'hc91d:	data_out=16'h8a00;
17'hc91e:	data_out=16'h86f2;
17'hc91f:	data_out=16'h9ba;
17'hc920:	data_out=16'h89fe;
17'hc921:	data_out=16'ha00;
17'hc922:	data_out=16'h8532;
17'hc923:	data_out=16'ha00;
17'hc924:	data_out=16'ha00;
17'hc925:	data_out=16'ha00;
17'hc926:	data_out=16'ha00;
17'hc927:	data_out=16'h89e9;
17'hc928:	data_out=16'ha00;
17'hc929:	data_out=16'h89ff;
17'hc92a:	data_out=16'h12e;
17'hc92b:	data_out=16'h8a00;
17'hc92c:	data_out=16'h8909;
17'hc92d:	data_out=16'h8a00;
17'hc92e:	data_out=16'h8605;
17'hc92f:	data_out=16'h89f5;
17'hc930:	data_out=16'ha00;
17'hc931:	data_out=16'h89ff;
17'hc932:	data_out=16'h195;
17'hc933:	data_out=16'h89eb;
17'hc934:	data_out=16'h8a00;
17'hc935:	data_out=16'h9ff;
17'hc936:	data_out=16'h87b4;
17'hc937:	data_out=16'h9fc;
17'hc938:	data_out=16'h8a00;
17'hc939:	data_out=16'h89f3;
17'hc93a:	data_out=16'h9ff;
17'hc93b:	data_out=16'ha00;
17'hc93c:	data_out=16'h89ff;
17'hc93d:	data_out=16'h89f0;
17'hc93e:	data_out=16'ha00;
17'hc93f:	data_out=16'h8943;
17'hc940:	data_out=16'h8955;
17'hc941:	data_out=16'h8236;
17'hc942:	data_out=16'ha00;
17'hc943:	data_out=16'h8a00;
17'hc944:	data_out=16'h1de;
17'hc945:	data_out=16'h895c;
17'hc946:	data_out=16'h8a00;
17'hc947:	data_out=16'h996;
17'hc948:	data_out=16'h88ba;
17'hc949:	data_out=16'ha00;
17'hc94a:	data_out=16'h13a;
17'hc94b:	data_out=16'h9e8;
17'hc94c:	data_out=16'h9fb;
17'hc94d:	data_out=16'h89e2;
17'hc94e:	data_out=16'h899d;
17'hc94f:	data_out=16'h9fe;
17'hc950:	data_out=16'h89e6;
17'hc951:	data_out=16'ha00;
17'hc952:	data_out=16'ha00;
17'hc953:	data_out=16'h89f3;
17'hc954:	data_out=16'h8a00;
17'hc955:	data_out=16'ha00;
17'hc956:	data_out=16'ha00;
17'hc957:	data_out=16'h9fe;
17'hc958:	data_out=16'ha00;
17'hc959:	data_out=16'h89d1;
17'hc95a:	data_out=16'h87ba;
17'hc95b:	data_out=16'h89c6;
17'hc95c:	data_out=16'h89c0;
17'hc95d:	data_out=16'h89b0;
17'hc95e:	data_out=16'h891c;
17'hc95f:	data_out=16'h8a00;
17'hc960:	data_out=16'h9fa;
17'hc961:	data_out=16'h890a;
17'hc962:	data_out=16'h883d;
17'hc963:	data_out=16'h89ec;
17'hc964:	data_out=16'h8a00;
17'hc965:	data_out=16'h89fe;
17'hc966:	data_out=16'h9fd;
17'hc967:	data_out=16'h8086;
17'hc968:	data_out=16'ha00;
17'hc969:	data_out=16'h9d6;
17'hc96a:	data_out=16'ha00;
17'hc96b:	data_out=16'h89f1;
17'hc96c:	data_out=16'h8a00;
17'hc96d:	data_out=16'h89ee;
17'hc96e:	data_out=16'ha00;
17'hc96f:	data_out=16'h89b6;
17'hc970:	data_out=16'ha00;
17'hc971:	data_out=16'h4f6;
17'hc972:	data_out=16'h8a00;
17'hc973:	data_out=16'h8a00;
17'hc974:	data_out=16'ha00;
17'hc975:	data_out=16'h8850;
17'hc976:	data_out=16'h8a1;
17'hc977:	data_out=16'ha00;
17'hc978:	data_out=16'h8a00;
17'hc979:	data_out=16'h779;
17'hc97a:	data_out=16'h8946;
17'hc97b:	data_out=16'ha00;
17'hc97c:	data_out=16'h895d;
17'hc97d:	data_out=16'h9f2;
17'hc97e:	data_out=16'h9ff;
17'hc97f:	data_out=16'h8a00;
17'hc980:	data_out=16'h8a00;
17'hc981:	data_out=16'h8a00;
17'hc982:	data_out=16'h70a;
17'hc983:	data_out=16'h89c2;
17'hc984:	data_out=16'h8133;
17'hc985:	data_out=16'h87ec;
17'hc986:	data_out=16'h9d6;
17'hc987:	data_out=16'ha00;
17'hc988:	data_out=16'h89c4;
17'hc989:	data_out=16'h9ff;
17'hc98a:	data_out=16'h8a00;
17'hc98b:	data_out=16'h89e5;
17'hc98c:	data_out=16'h9d3;
17'hc98d:	data_out=16'h87e3;
17'hc98e:	data_out=16'ha00;
17'hc98f:	data_out=16'h830c;
17'hc990:	data_out=16'h89e6;
17'hc991:	data_out=16'h8372;
17'hc992:	data_out=16'h89fc;
17'hc993:	data_out=16'h89cf;
17'hc994:	data_out=16'h89e0;
17'hc995:	data_out=16'h89ee;
17'hc996:	data_out=16'h89e7;
17'hc997:	data_out=16'h89e4;
17'hc998:	data_out=16'h87ab;
17'hc999:	data_out=16'h8a00;
17'hc99a:	data_out=16'h89bc;
17'hc99b:	data_out=16'h897e;
17'hc99c:	data_out=16'h89c8;
17'hc99d:	data_out=16'h8a00;
17'hc99e:	data_out=16'h89ee;
17'hc99f:	data_out=16'h9c9;
17'hc9a0:	data_out=16'h89ff;
17'hc9a1:	data_out=16'ha00;
17'hc9a2:	data_out=16'h86c2;
17'hc9a3:	data_out=16'ha00;
17'hc9a4:	data_out=16'ha00;
17'hc9a5:	data_out=16'ha00;
17'hc9a6:	data_out=16'h9fe;
17'hc9a7:	data_out=16'h89fa;
17'hc9a8:	data_out=16'ha00;
17'hc9a9:	data_out=16'h8a00;
17'hc9aa:	data_out=16'h879b;
17'hc9ab:	data_out=16'h8a00;
17'hc9ac:	data_out=16'h89f0;
17'hc9ad:	data_out=16'h8a00;
17'hc9ae:	data_out=16'h89de;
17'hc9af:	data_out=16'h89ff;
17'hc9b0:	data_out=16'h9ff;
17'hc9b1:	data_out=16'h89ff;
17'hc9b2:	data_out=16'h41a;
17'hc9b3:	data_out=16'h89fd;
17'hc9b4:	data_out=16'h8a00;
17'hc9b5:	data_out=16'h895b;
17'hc9b6:	data_out=16'h89d1;
17'hc9b7:	data_out=16'h9f;
17'hc9b8:	data_out=16'h8a00;
17'hc9b9:	data_out=16'h89fe;
17'hc9ba:	data_out=16'h97;
17'hc9bb:	data_out=16'ha00;
17'hc9bc:	data_out=16'h8a00;
17'hc9bd:	data_out=16'h89f1;
17'hc9be:	data_out=16'ha00;
17'hc9bf:	data_out=16'h87d4;
17'hc9c0:	data_out=16'h8821;
17'hc9c1:	data_out=16'h88c9;
17'hc9c2:	data_out=16'h88f9;
17'hc9c3:	data_out=16'h8888;
17'hc9c4:	data_out=16'h8913;
17'hc9c5:	data_out=16'h89ef;
17'hc9c6:	data_out=16'h8a00;
17'hc9c7:	data_out=16'h89fd;
17'hc9c8:	data_out=16'h89d7;
17'hc9c9:	data_out=16'ha00;
17'hc9ca:	data_out=16'h89ed;
17'hc9cb:	data_out=16'h898f;
17'hc9cc:	data_out=16'h9ff;
17'hc9cd:	data_out=16'h8996;
17'hc9ce:	data_out=16'h89e0;
17'hc9cf:	data_out=16'h9fe;
17'hc9d0:	data_out=16'h89fa;
17'hc9d1:	data_out=16'ha00;
17'hc9d2:	data_out=16'ha00;
17'hc9d3:	data_out=16'h89ff;
17'hc9d4:	data_out=16'h8a00;
17'hc9d5:	data_out=16'h81d5;
17'hc9d6:	data_out=16'h9fe;
17'hc9d7:	data_out=16'h9fe;
17'hc9d8:	data_out=16'h8432;
17'hc9d9:	data_out=16'h8994;
17'hc9da:	data_out=16'h89d5;
17'hc9db:	data_out=16'h89ec;
17'hc9dc:	data_out=16'h89d5;
17'hc9dd:	data_out=16'h89ca;
17'hc9de:	data_out=16'h88e9;
17'hc9df:	data_out=16'h8a00;
17'hc9e0:	data_out=16'h8b7;
17'hc9e1:	data_out=16'h8515;
17'hc9e2:	data_out=16'h89c2;
17'hc9e3:	data_out=16'h89fd;
17'hc9e4:	data_out=16'h8a00;
17'hc9e5:	data_out=16'h8a00;
17'hc9e6:	data_out=16'h9f1;
17'hc9e7:	data_out=16'h8a00;
17'hc9e8:	data_out=16'ha00;
17'hc9e9:	data_out=16'h89c6;
17'hc9ea:	data_out=16'ha00;
17'hc9eb:	data_out=16'h89f2;
17'hc9ec:	data_out=16'h8a00;
17'hc9ed:	data_out=16'h89fe;
17'hc9ee:	data_out=16'ha00;
17'hc9ef:	data_out=16'h89ec;
17'hc9f0:	data_out=16'ha00;
17'hc9f1:	data_out=16'h87f5;
17'hc9f2:	data_out=16'h8a00;
17'hc9f3:	data_out=16'h8a00;
17'hc9f4:	data_out=16'h9ff;
17'hc9f5:	data_out=16'ha00;
17'hc9f6:	data_out=16'h879d;
17'hc9f7:	data_out=16'h865c;
17'hc9f8:	data_out=16'h8a00;
17'hc9f9:	data_out=16'h8939;
17'hc9fa:	data_out=16'h89f5;
17'hc9fb:	data_out=16'ha00;
17'hc9fc:	data_out=16'h8969;
17'hc9fd:	data_out=16'h9d6;
17'hc9fe:	data_out=16'h9ff;
17'hc9ff:	data_out=16'h89fc;
17'hca00:	data_out=16'h8a00;
17'hca01:	data_out=16'h8a00;
17'hca02:	data_out=16'h80f0;
17'hca03:	data_out=16'h89f4;
17'hca04:	data_out=16'h881;
17'hca05:	data_out=16'ha00;
17'hca06:	data_out=16'h9d8;
17'hca07:	data_out=16'h97c;
17'hca08:	data_out=16'h8a00;
17'hca09:	data_out=16'h89b9;
17'hca0a:	data_out=16'h89f7;
17'hca0b:	data_out=16'h8a00;
17'hca0c:	data_out=16'h8a00;
17'hca0d:	data_out=16'h89f0;
17'hca0e:	data_out=16'ha00;
17'hca0f:	data_out=16'h89fa;
17'hca10:	data_out=16'h89ff;
17'hca11:	data_out=16'h564;
17'hca12:	data_out=16'h8a00;
17'hca13:	data_out=16'h89bc;
17'hca14:	data_out=16'h89e1;
17'hca15:	data_out=16'h89e6;
17'hca16:	data_out=16'h89fc;
17'hca17:	data_out=16'h89db;
17'hca18:	data_out=16'h89fc;
17'hca19:	data_out=16'h89fe;
17'hca1a:	data_out=16'ha00;
17'hca1b:	data_out=16'h89e4;
17'hca1c:	data_out=16'h8507;
17'hca1d:	data_out=16'h8a00;
17'hca1e:	data_out=16'h89fb;
17'hca1f:	data_out=16'h99d;
17'hca20:	data_out=16'h89f3;
17'hca21:	data_out=16'ha00;
17'hca22:	data_out=16'h88d7;
17'hca23:	data_out=16'ha00;
17'hca24:	data_out=16'ha00;
17'hca25:	data_out=16'ha00;
17'hca26:	data_out=16'h89e6;
17'hca27:	data_out=16'h89fd;
17'hca28:	data_out=16'ha00;
17'hca29:	data_out=16'h8a00;
17'hca2a:	data_out=16'h89fb;
17'hca2b:	data_out=16'h8a00;
17'hca2c:	data_out=16'h89fb;
17'hca2d:	data_out=16'h8a00;
17'hca2e:	data_out=16'h89ff;
17'hca2f:	data_out=16'h89fe;
17'hca30:	data_out=16'ha00;
17'hca31:	data_out=16'h89a5;
17'hca32:	data_out=16'ha00;
17'hca33:	data_out=16'h89fe;
17'hca34:	data_out=16'h8a00;
17'hca35:	data_out=16'h89f0;
17'hca36:	data_out=16'h89fb;
17'hca37:	data_out=16'h86ad;
17'hca38:	data_out=16'h9f9;
17'hca39:	data_out=16'h89ff;
17'hca3a:	data_out=16'h8a00;
17'hca3b:	data_out=16'ha00;
17'hca3c:	data_out=16'h89d6;
17'hca3d:	data_out=16'h89ec;
17'hca3e:	data_out=16'ha00;
17'hca3f:	data_out=16'ha00;
17'hca40:	data_out=16'h9eb;
17'hca41:	data_out=16'h89a5;
17'hca42:	data_out=16'h89e7;
17'hca43:	data_out=16'h950;
17'hca44:	data_out=16'h232;
17'hca45:	data_out=16'h89f5;
17'hca46:	data_out=16'h8a00;
17'hca47:	data_out=16'h8a00;
17'hca48:	data_out=16'h8a00;
17'hca49:	data_out=16'h9fb;
17'hca4a:	data_out=16'h8a00;
17'hca4b:	data_out=16'h8a00;
17'hca4c:	data_out=16'h246;
17'hca4d:	data_out=16'h8957;
17'hca4e:	data_out=16'h8a00;
17'hca4f:	data_out=16'h89ca;
17'hca50:	data_out=16'h89f7;
17'hca51:	data_out=16'h9e3;
17'hca52:	data_out=16'h9f6;
17'hca53:	data_out=16'h89fa;
17'hca54:	data_out=16'h89ff;
17'hca55:	data_out=16'h8984;
17'hca56:	data_out=16'h860d;
17'hca57:	data_out=16'h9d0;
17'hca58:	data_out=16'h9df;
17'hca59:	data_out=16'h9a9;
17'hca5a:	data_out=16'h89d4;
17'hca5b:	data_out=16'h570;
17'hca5c:	data_out=16'h87a2;
17'hca5d:	data_out=16'h89c0;
17'hca5e:	data_out=16'h887f;
17'hca5f:	data_out=16'h8a00;
17'hca60:	data_out=16'h89ff;
17'hca61:	data_out=16'ha00;
17'hca62:	data_out=16'h89fd;
17'hca63:	data_out=16'h89fe;
17'hca64:	data_out=16'h8a00;
17'hca65:	data_out=16'h89f0;
17'hca66:	data_out=16'h3e6;
17'hca67:	data_out=16'h8a00;
17'hca68:	data_out=16'ha00;
17'hca69:	data_out=16'h8a00;
17'hca6a:	data_out=16'ha00;
17'hca6b:	data_out=16'hb8;
17'hca6c:	data_out=16'h8a00;
17'hca6d:	data_out=16'h89ff;
17'hca6e:	data_out=16'ha00;
17'hca6f:	data_out=16'h279;
17'hca70:	data_out=16'ha00;
17'hca71:	data_out=16'h89fe;
17'hca72:	data_out=16'h9c0;
17'hca73:	data_out=16'h9e8;
17'hca74:	data_out=16'ha00;
17'hca75:	data_out=16'ha00;
17'hca76:	data_out=16'h8a00;
17'hca77:	data_out=16'h89da;
17'hca78:	data_out=16'h473;
17'hca79:	data_out=16'h89fd;
17'hca7a:	data_out=16'h89f4;
17'hca7b:	data_out=16'ha00;
17'hca7c:	data_out=16'h89fd;
17'hca7d:	data_out=16'h9ff;
17'hca7e:	data_out=16'h92a;
17'hca7f:	data_out=16'h9f1;
17'hca80:	data_out=16'h89ff;
17'hca81:	data_out=16'h89fc;
17'hca82:	data_out=16'h972;
17'hca83:	data_out=16'h89e7;
17'hca84:	data_out=16'h23e;
17'hca85:	data_out=16'ha00;
17'hca86:	data_out=16'h9e9;
17'hca87:	data_out=16'h8a00;
17'hca88:	data_out=16'h8a00;
17'hca89:	data_out=16'h8a00;
17'hca8a:	data_out=16'h89e4;
17'hca8b:	data_out=16'h8a00;
17'hca8c:	data_out=16'h8a00;
17'hca8d:	data_out=16'h8a00;
17'hca8e:	data_out=16'ha00;
17'hca8f:	data_out=16'h89ff;
17'hca90:	data_out=16'h89f8;
17'hca91:	data_out=16'h7b6;
17'hca92:	data_out=16'h8a00;
17'hca93:	data_out=16'h840c;
17'hca94:	data_out=16'h8527;
17'hca95:	data_out=16'h88f3;
17'hca96:	data_out=16'h89f9;
17'hca97:	data_out=16'h864f;
17'hca98:	data_out=16'h8a00;
17'hca99:	data_out=16'h8a00;
17'hca9a:	data_out=16'ha00;
17'hca9b:	data_out=16'h89f0;
17'hca9c:	data_out=16'h9f8;
17'hca9d:	data_out=16'h89ff;
17'hca9e:	data_out=16'h8984;
17'hca9f:	data_out=16'h9ce;
17'hcaa0:	data_out=16'h88b9;
17'hcaa1:	data_out=16'ha00;
17'hcaa2:	data_out=16'h7e0;
17'hcaa3:	data_out=16'h8a00;
17'hcaa4:	data_out=16'h8a00;
17'hcaa5:	data_out=16'h9ce;
17'hcaa6:	data_out=16'h8a00;
17'hcaa7:	data_out=16'h89ff;
17'hcaa8:	data_out=16'ha00;
17'hcaa9:	data_out=16'h8a00;
17'hcaaa:	data_out=16'h89fe;
17'hcaab:	data_out=16'h8a00;
17'hcaac:	data_out=16'h89e5;
17'hcaad:	data_out=16'h8a00;
17'hcaae:	data_out=16'h89d2;
17'hcaaf:	data_out=16'h89f8;
17'hcab0:	data_out=16'h9fc;
17'hcab1:	data_out=16'h83f5;
17'hcab2:	data_out=16'h9f9;
17'hcab3:	data_out=16'h8866;
17'hcab4:	data_out=16'h8a00;
17'hcab5:	data_out=16'h89fc;
17'hcab6:	data_out=16'h89fd;
17'hcab7:	data_out=16'h980;
17'hcab8:	data_out=16'ha00;
17'hcab9:	data_out=16'h89a5;
17'hcaba:	data_out=16'h8a00;
17'hcabb:	data_out=16'h89f5;
17'hcabc:	data_out=16'h9e3;
17'hcabd:	data_out=16'h87d2;
17'hcabe:	data_out=16'ha00;
17'hcabf:	data_out=16'ha00;
17'hcac0:	data_out=16'h9ee;
17'hcac1:	data_out=16'h89e4;
17'hcac2:	data_out=16'h8a00;
17'hcac3:	data_out=16'ha00;
17'hcac4:	data_out=16'h8495;
17'hcac5:	data_out=16'h8901;
17'hcac6:	data_out=16'h8a00;
17'hcac7:	data_out=16'h8a00;
17'hcac8:	data_out=16'h89ff;
17'hcac9:	data_out=16'h89a;
17'hcaca:	data_out=16'h8a00;
17'hcacb:	data_out=16'h8a00;
17'hcacc:	data_out=16'h8759;
17'hcacd:	data_out=16'h8547;
17'hcace:	data_out=16'h8a00;
17'hcacf:	data_out=16'h8a00;
17'hcad0:	data_out=16'h6a9;
17'hcad1:	data_out=16'h9f2;
17'hcad2:	data_out=16'h8a00;
17'hcad3:	data_out=16'h89db;
17'hcad4:	data_out=16'h89ef;
17'hcad5:	data_out=16'h8ff;
17'hcad6:	data_out=16'h824e;
17'hcad7:	data_out=16'h9d8;
17'hcad8:	data_out=16'ha00;
17'hcad9:	data_out=16'h9c9;
17'hcada:	data_out=16'h8ce;
17'hcadb:	data_out=16'h9f5;
17'hcadc:	data_out=16'ha00;
17'hcadd:	data_out=16'h8932;
17'hcade:	data_out=16'h8758;
17'hcadf:	data_out=16'h8a00;
17'hcae0:	data_out=16'h8a00;
17'hcae1:	data_out=16'ha00;
17'hcae2:	data_out=16'h8974;
17'hcae3:	data_out=16'h888e;
17'hcae4:	data_out=16'h8a00;
17'hcae5:	data_out=16'h89fe;
17'hcae6:	data_out=16'h89ef;
17'hcae7:	data_out=16'h89f9;
17'hcae8:	data_out=16'ha00;
17'hcae9:	data_out=16'h8a00;
17'hcaea:	data_out=16'ha00;
17'hcaeb:	data_out=16'ha00;
17'hcaec:	data_out=16'h89fb;
17'hcaed:	data_out=16'h88b1;
17'hcaee:	data_out=16'ha00;
17'hcaef:	data_out=16'h9fc;
17'hcaf0:	data_out=16'ha00;
17'hcaf1:	data_out=16'h8a00;
17'hcaf2:	data_out=16'ha00;
17'hcaf3:	data_out=16'ha00;
17'hcaf4:	data_out=16'h9fb;
17'hcaf5:	data_out=16'ha00;
17'hcaf6:	data_out=16'h8a00;
17'hcaf7:	data_out=16'h89ff;
17'hcaf8:	data_out=16'ha00;
17'hcaf9:	data_out=16'h8a00;
17'hcafa:	data_out=16'h8870;
17'hcafb:	data_out=16'ha00;
17'hcafc:	data_out=16'h8a00;
17'hcafd:	data_out=16'ha00;
17'hcafe:	data_out=16'ha00;
17'hcaff:	data_out=16'ha00;
17'hcb00:	data_out=16'h89fc;
17'hcb01:	data_out=16'h8a00;
17'hcb02:	data_out=16'h89fe;
17'hcb03:	data_out=16'h98c;
17'hcb04:	data_out=16'h89f2;
17'hcb05:	data_out=16'ha00;
17'hcb06:	data_out=16'ha00;
17'hcb07:	data_out=16'h8a00;
17'hcb08:	data_out=16'h8a00;
17'hcb09:	data_out=16'h8a00;
17'hcb0a:	data_out=16'h8a00;
17'hcb0b:	data_out=16'h8a00;
17'hcb0c:	data_out=16'h8a00;
17'hcb0d:	data_out=16'h89f8;
17'hcb0e:	data_out=16'ha00;
17'hcb0f:	data_out=16'h8a00;
17'hcb10:	data_out=16'h89ec;
17'hcb11:	data_out=16'h89fc;
17'hcb12:	data_out=16'h89ff;
17'hcb13:	data_out=16'ha00;
17'hcb14:	data_out=16'h9f2;
17'hcb15:	data_out=16'h897f;
17'hcb16:	data_out=16'h89f7;
17'hcb17:	data_out=16'h9cd;
17'hcb18:	data_out=16'h8a00;
17'hcb19:	data_out=16'h8a00;
17'hcb1a:	data_out=16'ha00;
17'hcb1b:	data_out=16'h475;
17'hcb1c:	data_out=16'ha00;
17'hcb1d:	data_out=16'h8a00;
17'hcb1e:	data_out=16'h5da;
17'hcb1f:	data_out=16'h9ff;
17'hcb20:	data_out=16'h8671;
17'hcb21:	data_out=16'ha00;
17'hcb22:	data_out=16'h9e9;
17'hcb23:	data_out=16'h8a00;
17'hcb24:	data_out=16'h8a00;
17'hcb25:	data_out=16'h89c6;
17'hcb26:	data_out=16'h8a00;
17'hcb27:	data_out=16'h8a00;
17'hcb28:	data_out=16'ha00;
17'hcb29:	data_out=16'h89ff;
17'hcb2a:	data_out=16'h89ff;
17'hcb2b:	data_out=16'h8a00;
17'hcb2c:	data_out=16'h8897;
17'hcb2d:	data_out=16'h8a00;
17'hcb2e:	data_out=16'h826e;
17'hcb2f:	data_out=16'h877b;
17'hcb30:	data_out=16'h41f;
17'hcb31:	data_out=16'h8a00;
17'hcb32:	data_out=16'h817;
17'hcb33:	data_out=16'ha00;
17'hcb34:	data_out=16'h8a00;
17'hcb35:	data_out=16'h8a00;
17'hcb36:	data_out=16'h89ff;
17'hcb37:	data_out=16'h89fc;
17'hcb38:	data_out=16'ha00;
17'hcb39:	data_out=16'ha00;
17'hcb3a:	data_out=16'h8a00;
17'hcb3b:	data_out=16'h8a00;
17'hcb3c:	data_out=16'h9b8;
17'hcb3d:	data_out=16'h869d;
17'hcb3e:	data_out=16'ha00;
17'hcb3f:	data_out=16'ha00;
17'hcb40:	data_out=16'h9b7;
17'hcb41:	data_out=16'h8a00;
17'hcb42:	data_out=16'h8a00;
17'hcb43:	data_out=16'ha00;
17'hcb44:	data_out=16'h89ff;
17'hcb45:	data_out=16'h896e;
17'hcb46:	data_out=16'h8a00;
17'hcb47:	data_out=16'h8a00;
17'hcb48:	data_out=16'h8426;
17'hcb49:	data_out=16'h89fd;
17'hcb4a:	data_out=16'h8a00;
17'hcb4b:	data_out=16'h8a00;
17'hcb4c:	data_out=16'h89fc;
17'hcb4d:	data_out=16'h9f3;
17'hcb4e:	data_out=16'h8a00;
17'hcb4f:	data_out=16'h8a00;
17'hcb50:	data_out=16'h9c8;
17'hcb51:	data_out=16'ha00;
17'hcb52:	data_out=16'h8a00;
17'hcb53:	data_out=16'h8995;
17'hcb54:	data_out=16'h8993;
17'hcb55:	data_out=16'h8e0;
17'hcb56:	data_out=16'h8a00;
17'hcb57:	data_out=16'h941;
17'hcb58:	data_out=16'ha00;
17'hcb59:	data_out=16'h9ab;
17'hcb5a:	data_out=16'h9d9;
17'hcb5b:	data_out=16'h89f9;
17'hcb5c:	data_out=16'ha00;
17'hcb5d:	data_out=16'h87f7;
17'hcb5e:	data_out=16'h849a;
17'hcb5f:	data_out=16'h89fe;
17'hcb60:	data_out=16'h8a00;
17'hcb61:	data_out=16'h9e3;
17'hcb62:	data_out=16'h86e1;
17'hcb63:	data_out=16'ha00;
17'hcb64:	data_out=16'h8a00;
17'hcb65:	data_out=16'h8a00;
17'hcb66:	data_out=16'h8a00;
17'hcb67:	data_out=16'h8900;
17'hcb68:	data_out=16'ha00;
17'hcb69:	data_out=16'h8a00;
17'hcb6a:	data_out=16'ha00;
17'hcb6b:	data_out=16'ha00;
17'hcb6c:	data_out=16'h89f7;
17'hcb6d:	data_out=16'ha00;
17'hcb6e:	data_out=16'ha00;
17'hcb6f:	data_out=16'h9cf;
17'hcb70:	data_out=16'ha00;
17'hcb71:	data_out=16'h8a00;
17'hcb72:	data_out=16'h9df;
17'hcb73:	data_out=16'h9e4;
17'hcb74:	data_out=16'h3c0;
17'hcb75:	data_out=16'ha00;
17'hcb76:	data_out=16'h8a00;
17'hcb77:	data_out=16'h8a00;
17'hcb78:	data_out=16'ha00;
17'hcb79:	data_out=16'h8a00;
17'hcb7a:	data_out=16'h9f5;
17'hcb7b:	data_out=16'ha00;
17'hcb7c:	data_out=16'h8a00;
17'hcb7d:	data_out=16'ha00;
17'hcb7e:	data_out=16'ha00;
17'hcb7f:	data_out=16'ha00;
17'hcb80:	data_out=16'h8a00;
17'hcb81:	data_out=16'h8a00;
17'hcb82:	data_out=16'h8a00;
17'hcb83:	data_out=16'h9af;
17'hcb84:	data_out=16'h8a00;
17'hcb85:	data_out=16'h9de;
17'hcb86:	data_out=16'ha00;
17'hcb87:	data_out=16'h8a00;
17'hcb88:	data_out=16'h8a00;
17'hcb89:	data_out=16'h89ff;
17'hcb8a:	data_out=16'h8a00;
17'hcb8b:	data_out=16'h8a00;
17'hcb8c:	data_out=16'h8a00;
17'hcb8d:	data_out=16'h991;
17'hcb8e:	data_out=16'ha00;
17'hcb8f:	data_out=16'h8a00;
17'hcb90:	data_out=16'h89c2;
17'hcb91:	data_out=16'h8a00;
17'hcb92:	data_out=16'h912;
17'hcb93:	data_out=16'ha00;
17'hcb94:	data_out=16'ha00;
17'hcb95:	data_out=16'h89fe;
17'hcb96:	data_out=16'h89fd;
17'hcb97:	data_out=16'h9dd;
17'hcb98:	data_out=16'h8a00;
17'hcb99:	data_out=16'h8a00;
17'hcb9a:	data_out=16'h9e4;
17'hcb9b:	data_out=16'h8c0;
17'hcb9c:	data_out=16'h9e2;
17'hcb9d:	data_out=16'h8a00;
17'hcb9e:	data_out=16'h9e5;
17'hcb9f:	data_out=16'h9f9;
17'hcba0:	data_out=16'h897a;
17'hcba1:	data_out=16'ha00;
17'hcba2:	data_out=16'h9f4;
17'hcba3:	data_out=16'h8a00;
17'hcba4:	data_out=16'h8a00;
17'hcba5:	data_out=16'h89a2;
17'hcba6:	data_out=16'h8a00;
17'hcba7:	data_out=16'h8a00;
17'hcba8:	data_out=16'ha00;
17'hcba9:	data_out=16'h7ed;
17'hcbaa:	data_out=16'h8a00;
17'hcbab:	data_out=16'h8a00;
17'hcbac:	data_out=16'h89fb;
17'hcbad:	data_out=16'h8a00;
17'hcbae:	data_out=16'h9ea;
17'hcbaf:	data_out=16'h85f5;
17'hcbb0:	data_out=16'h8a00;
17'hcbb1:	data_out=16'h8a00;
17'hcbb2:	data_out=16'h8a00;
17'hcbb3:	data_out=16'ha00;
17'hcbb4:	data_out=16'h8a00;
17'hcbb5:	data_out=16'h8a00;
17'hcbb6:	data_out=16'h8a00;
17'hcbb7:	data_out=16'h8907;
17'hcbb8:	data_out=16'ha00;
17'hcbb9:	data_out=16'ha00;
17'hcbba:	data_out=16'h8a00;
17'hcbbb:	data_out=16'h8a00;
17'hcbbc:	data_out=16'h959;
17'hcbbd:	data_out=16'h89aa;
17'hcbbe:	data_out=16'ha00;
17'hcbbf:	data_out=16'h9de;
17'hcbc0:	data_out=16'h88e4;
17'hcbc1:	data_out=16'h8a00;
17'hcbc2:	data_out=16'h8a00;
17'hcbc3:	data_out=16'ha00;
17'hcbc4:	data_out=16'h8a00;
17'hcbc5:	data_out=16'h89fe;
17'hcbc6:	data_out=16'h8a00;
17'hcbc7:	data_out=16'h8a00;
17'hcbc8:	data_out=16'h9c1;
17'hcbc9:	data_out=16'h89fb;
17'hcbca:	data_out=16'h8a00;
17'hcbcb:	data_out=16'h8a00;
17'hcbcc:	data_out=16'h89d7;
17'hcbcd:	data_out=16'h9ef;
17'hcbce:	data_out=16'h8215;
17'hcbcf:	data_out=16'h8a00;
17'hcbd0:	data_out=16'ha00;
17'hcbd1:	data_out=16'h9fb;
17'hcbd2:	data_out=16'h8a00;
17'hcbd3:	data_out=16'h8a00;
17'hcbd4:	data_out=16'h89c9;
17'hcbd5:	data_out=16'h981;
17'hcbd6:	data_out=16'h8a00;
17'hcbd7:	data_out=16'h89d2;
17'hcbd8:	data_out=16'h9fe;
17'hcbd9:	data_out=16'h8907;
17'hcbda:	data_out=16'h9da;
17'hcbdb:	data_out=16'h8a00;
17'hcbdc:	data_out=16'h9f4;
17'hcbdd:	data_out=16'h87d4;
17'hcbde:	data_out=16'h8319;
17'hcbdf:	data_out=16'h8a00;
17'hcbe0:	data_out=16'h8a00;
17'hcbe1:	data_out=16'h8a00;
17'hcbe2:	data_out=16'h9c0;
17'hcbe3:	data_out=16'ha00;
17'hcbe4:	data_out=16'h8a00;
17'hcbe5:	data_out=16'h8a00;
17'hcbe6:	data_out=16'h8a00;
17'hcbe7:	data_out=16'h9da;
17'hcbe8:	data_out=16'ha00;
17'hcbe9:	data_out=16'h8a00;
17'hcbea:	data_out=16'ha00;
17'hcbeb:	data_out=16'h9eb;
17'hcbec:	data_out=16'h89ff;
17'hcbed:	data_out=16'ha00;
17'hcbee:	data_out=16'ha00;
17'hcbef:	data_out=16'h9ae;
17'hcbf0:	data_out=16'ha00;
17'hcbf1:	data_out=16'h8a00;
17'hcbf2:	data_out=16'h9c8;
17'hcbf3:	data_out=16'h99f;
17'hcbf4:	data_out=16'h8a00;
17'hcbf5:	data_out=16'h9e3;
17'hcbf6:	data_out=16'h8a00;
17'hcbf7:	data_out=16'h89f0;
17'hcbf8:	data_out=16'ha00;
17'hcbf9:	data_out=16'h89c7;
17'hcbfa:	data_out=16'ha00;
17'hcbfb:	data_out=16'ha00;
17'hcbfc:	data_out=16'h8a00;
17'hcbfd:	data_out=16'ha00;
17'hcbfe:	data_out=16'h9ff;
17'hcbff:	data_out=16'ha00;
17'hcc00:	data_out=16'h8a00;
17'hcc01:	data_out=16'h8a00;
17'hcc02:	data_out=16'h9b8;
17'hcc03:	data_out=16'ha00;
17'hcc04:	data_out=16'h8a00;
17'hcc05:	data_out=16'h89dc;
17'hcc06:	data_out=16'ha00;
17'hcc07:	data_out=16'h8a00;
17'hcc08:	data_out=16'h8a00;
17'hcc09:	data_out=16'h874f;
17'hcc0a:	data_out=16'h8a00;
17'hcc0b:	data_out=16'h896d;
17'hcc0c:	data_out=16'h8a00;
17'hcc0d:	data_out=16'h9de;
17'hcc0e:	data_out=16'ha00;
17'hcc0f:	data_out=16'h464;
17'hcc10:	data_out=16'h81c6;
17'hcc11:	data_out=16'h8a00;
17'hcc12:	data_out=16'h9de;
17'hcc13:	data_out=16'ha00;
17'hcc14:	data_out=16'ha00;
17'hcc15:	data_out=16'h8a00;
17'hcc16:	data_out=16'h8a00;
17'hcc17:	data_out=16'ha00;
17'hcc18:	data_out=16'h8a00;
17'hcc19:	data_out=16'h8a00;
17'hcc1a:	data_out=16'h89fd;
17'hcc1b:	data_out=16'h9cd;
17'hcc1c:	data_out=16'ha00;
17'hcc1d:	data_out=16'h8a00;
17'hcc1e:	data_out=16'h9fe;
17'hcc1f:	data_out=16'h9e1;
17'hcc20:	data_out=16'h89fc;
17'hcc21:	data_out=16'ha00;
17'hcc22:	data_out=16'ha00;
17'hcc23:	data_out=16'h8a00;
17'hcc24:	data_out=16'h8a00;
17'hcc25:	data_out=16'h8967;
17'hcc26:	data_out=16'h8a00;
17'hcc27:	data_out=16'h8a00;
17'hcc28:	data_out=16'ha00;
17'hcc29:	data_out=16'h8d3;
17'hcc2a:	data_out=16'h89ff;
17'hcc2b:	data_out=16'h8a00;
17'hcc2c:	data_out=16'h8a00;
17'hcc2d:	data_out=16'h8a00;
17'hcc2e:	data_out=16'h9dc;
17'hcc2f:	data_out=16'h86bc;
17'hcc30:	data_out=16'h8a00;
17'hcc31:	data_out=16'h8a00;
17'hcc32:	data_out=16'h8a00;
17'hcc33:	data_out=16'ha00;
17'hcc34:	data_out=16'h8a00;
17'hcc35:	data_out=16'h8a00;
17'hcc36:	data_out=16'h8a00;
17'hcc37:	data_out=16'h9b7;
17'hcc38:	data_out=16'ha00;
17'hcc39:	data_out=16'ha00;
17'hcc3a:	data_out=16'h8a00;
17'hcc3b:	data_out=16'h8a00;
17'hcc3c:	data_out=16'h976;
17'hcc3d:	data_out=16'h89f4;
17'hcc3e:	data_out=16'ha00;
17'hcc3f:	data_out=16'h89e1;
17'hcc40:	data_out=16'h89fc;
17'hcc41:	data_out=16'h8a00;
17'hcc42:	data_out=16'h8a00;
17'hcc43:	data_out=16'ha00;
17'hcc44:	data_out=16'h8a00;
17'hcc45:	data_out=16'h8a00;
17'hcc46:	data_out=16'h8a00;
17'hcc47:	data_out=16'h89e9;
17'hcc48:	data_out=16'h9f4;
17'hcc49:	data_out=16'h89e9;
17'hcc4a:	data_out=16'h8a00;
17'hcc4b:	data_out=16'h8a00;
17'hcc4c:	data_out=16'h890d;
17'hcc4d:	data_out=16'ha00;
17'hcc4e:	data_out=16'h9da;
17'hcc4f:	data_out=16'h8a00;
17'hcc50:	data_out=16'ha00;
17'hcc51:	data_out=16'h9f8;
17'hcc52:	data_out=16'h8a00;
17'hcc53:	data_out=16'h8a00;
17'hcc54:	data_out=16'h89e8;
17'hcc55:	data_out=16'h9ce;
17'hcc56:	data_out=16'h8a00;
17'hcc57:	data_out=16'h6ec;
17'hcc58:	data_out=16'h9f3;
17'hcc59:	data_out=16'h8995;
17'hcc5a:	data_out=16'h9ff;
17'hcc5b:	data_out=16'h8a00;
17'hcc5c:	data_out=16'h9e6;
17'hcc5d:	data_out=16'h87f9;
17'hcc5e:	data_out=16'h82cc;
17'hcc5f:	data_out=16'h89ef;
17'hcc60:	data_out=16'h8a00;
17'hcc61:	data_out=16'h8a00;
17'hcc62:	data_out=16'h9f2;
17'hcc63:	data_out=16'ha00;
17'hcc64:	data_out=16'h8a00;
17'hcc65:	data_out=16'h8a00;
17'hcc66:	data_out=16'h8a00;
17'hcc67:	data_out=16'h96c;
17'hcc68:	data_out=16'ha00;
17'hcc69:	data_out=16'h8a00;
17'hcc6a:	data_out=16'ha00;
17'hcc6b:	data_out=16'h8928;
17'hcc6c:	data_out=16'h89ff;
17'hcc6d:	data_out=16'ha00;
17'hcc6e:	data_out=16'ha00;
17'hcc6f:	data_out=16'h8108;
17'hcc70:	data_out=16'ha00;
17'hcc71:	data_out=16'h88c5;
17'hcc72:	data_out=16'h886e;
17'hcc73:	data_out=16'h87d3;
17'hcc74:	data_out=16'h8a00;
17'hcc75:	data_out=16'h98f;
17'hcc76:	data_out=16'h8a00;
17'hcc77:	data_out=16'h8186;
17'hcc78:	data_out=16'ha00;
17'hcc79:	data_out=16'h879c;
17'hcc7a:	data_out=16'ha00;
17'hcc7b:	data_out=16'ha00;
17'hcc7c:	data_out=16'h8a00;
17'hcc7d:	data_out=16'h9fd;
17'hcc7e:	data_out=16'ha00;
17'hcc7f:	data_out=16'ha00;
17'hcc80:	data_out=16'h8a00;
17'hcc81:	data_out=16'h89fd;
17'hcc82:	data_out=16'ha00;
17'hcc83:	data_out=16'ha00;
17'hcc84:	data_out=16'h8a00;
17'hcc85:	data_out=16'h8a00;
17'hcc86:	data_out=16'h9ff;
17'hcc87:	data_out=16'h8a00;
17'hcc88:	data_out=16'h100;
17'hcc89:	data_out=16'h9c4;
17'hcc8a:	data_out=16'h89f7;
17'hcc8b:	data_out=16'ha00;
17'hcc8c:	data_out=16'h898f;
17'hcc8d:	data_out=16'h2a5;
17'hcc8e:	data_out=16'ha00;
17'hcc8f:	data_out=16'ha00;
17'hcc90:	data_out=16'ha00;
17'hcc91:	data_out=16'h89a1;
17'hcc92:	data_out=16'h9fa;
17'hcc93:	data_out=16'h9ff;
17'hcc94:	data_out=16'ha00;
17'hcc95:	data_out=16'h8a00;
17'hcc96:	data_out=16'h89f8;
17'hcc97:	data_out=16'ha00;
17'hcc98:	data_out=16'h7b5;
17'hcc99:	data_out=16'h5b8;
17'hcc9a:	data_out=16'h8a00;
17'hcc9b:	data_out=16'ha00;
17'hcc9c:	data_out=16'h123;
17'hcc9d:	data_out=16'h89ff;
17'hcc9e:	data_out=16'ha00;
17'hcc9f:	data_out=16'h9d8;
17'hcca0:	data_out=16'h89b4;
17'hcca1:	data_out=16'ha00;
17'hcca2:	data_out=16'ha00;
17'hcca3:	data_out=16'h8a00;
17'hcca4:	data_out=16'h8a00;
17'hcca5:	data_out=16'h9df;
17'hcca6:	data_out=16'h9f4;
17'hcca7:	data_out=16'h89f2;
17'hcca8:	data_out=16'ha00;
17'hcca9:	data_out=16'h9e9;
17'hccaa:	data_out=16'h9f3;
17'hccab:	data_out=16'h9fd;
17'hccac:	data_out=16'h8a00;
17'hccad:	data_out=16'h8711;
17'hccae:	data_out=16'ha00;
17'hccaf:	data_out=16'h87ef;
17'hccb0:	data_out=16'h8836;
17'hccb1:	data_out=16'h8a00;
17'hccb2:	data_out=16'h8a00;
17'hccb3:	data_out=16'ha00;
17'hccb4:	data_out=16'h8a00;
17'hccb5:	data_out=16'h8a00;
17'hccb6:	data_out=16'h26c;
17'hccb7:	data_out=16'ha00;
17'hccb8:	data_out=16'h897b;
17'hccb9:	data_out=16'ha00;
17'hccba:	data_out=16'h99a;
17'hccbb:	data_out=16'h8a00;
17'hccbc:	data_out=16'h9cc;
17'hccbd:	data_out=16'h8977;
17'hccbe:	data_out=16'ha00;
17'hccbf:	data_out=16'h8a00;
17'hccc0:	data_out=16'h89da;
17'hccc1:	data_out=16'h8708;
17'hccc2:	data_out=16'h89b1;
17'hccc3:	data_out=16'ha00;
17'hccc4:	data_out=16'h8a00;
17'hccc5:	data_out=16'h8a00;
17'hccc6:	data_out=16'ha00;
17'hccc7:	data_out=16'h9d0;
17'hccc8:	data_out=16'h9fe;
17'hccc9:	data_out=16'h9ca;
17'hccca:	data_out=16'h89db;
17'hcccb:	data_out=16'h89a2;
17'hcccc:	data_out=16'h9ea;
17'hcccd:	data_out=16'ha00;
17'hccce:	data_out=16'ha00;
17'hcccf:	data_out=16'h607;
17'hccd0:	data_out=16'h8915;
17'hccd1:	data_out=16'h9e8;
17'hccd2:	data_out=16'h89ff;
17'hccd3:	data_out=16'h88d8;
17'hccd4:	data_out=16'h893f;
17'hccd5:	data_out=16'h9fc;
17'hccd6:	data_out=16'h354;
17'hccd7:	data_out=16'h9b5;
17'hccd8:	data_out=16'ha00;
17'hccd9:	data_out=16'h8976;
17'hccda:	data_out=16'ha00;
17'hccdb:	data_out=16'h8a00;
17'hccdc:	data_out=16'h862a;
17'hccdd:	data_out=16'h88d2;
17'hccde:	data_out=16'h84aa;
17'hccdf:	data_out=16'h891a;
17'hcce0:	data_out=16'h810f;
17'hcce1:	data_out=16'h8a00;
17'hcce2:	data_out=16'ha00;
17'hcce3:	data_out=16'ha00;
17'hcce4:	data_out=16'h8a00;
17'hcce5:	data_out=16'h89df;
17'hcce6:	data_out=16'h9fc;
17'hcce7:	data_out=16'h9e8;
17'hcce8:	data_out=16'ha00;
17'hcce9:	data_out=16'h9f7;
17'hccea:	data_out=16'ha00;
17'hcceb:	data_out=16'h89b1;
17'hccec:	data_out=16'h89dc;
17'hcced:	data_out=16'ha00;
17'hccee:	data_out=16'ha00;
17'hccef:	data_out=16'h89f2;
17'hccf0:	data_out=16'ha00;
17'hccf1:	data_out=16'h9ee;
17'hccf2:	data_out=16'h8995;
17'hccf3:	data_out=16'h8989;
17'hccf4:	data_out=16'h89f9;
17'hccf5:	data_out=16'h8960;
17'hccf6:	data_out=16'ha00;
17'hccf7:	data_out=16'ha00;
17'hccf8:	data_out=16'h9aa;
17'hccf9:	data_out=16'ha00;
17'hccfa:	data_out=16'ha00;
17'hccfb:	data_out=16'ha00;
17'hccfc:	data_out=16'h89f5;
17'hccfd:	data_out=16'h9df;
17'hccfe:	data_out=16'ha00;
17'hccff:	data_out=16'h8a00;
17'hcd00:	data_out=16'h8a00;
17'hcd01:	data_out=16'h89df;
17'hcd02:	data_out=16'ha00;
17'hcd03:	data_out=16'h86cd;
17'hcd04:	data_out=16'h8a00;
17'hcd05:	data_out=16'h8a00;
17'hcd06:	data_out=16'h9f;
17'hcd07:	data_out=16'h997;
17'hcd08:	data_out=16'ha00;
17'hcd09:	data_out=16'h9e1;
17'hcd0a:	data_out=16'h899f;
17'hcd0b:	data_out=16'ha00;
17'hcd0c:	data_out=16'h9c2;
17'hcd0d:	data_out=16'h89e8;
17'hcd0e:	data_out=16'h9ff;
17'hcd0f:	data_out=16'ha00;
17'hcd10:	data_out=16'h392;
17'hcd11:	data_out=16'h8968;
17'hcd12:	data_out=16'h9f0;
17'hcd13:	data_out=16'h83fe;
17'hcd14:	data_out=16'ha00;
17'hcd15:	data_out=16'h8a00;
17'hcd16:	data_out=16'h8a00;
17'hcd17:	data_out=16'ha00;
17'hcd18:	data_out=16'h9ec;
17'hcd19:	data_out=16'ha00;
17'hcd1a:	data_out=16'h8a00;
17'hcd1b:	data_out=16'ha00;
17'hcd1c:	data_out=16'h8992;
17'hcd1d:	data_out=16'h89cc;
17'hcd1e:	data_out=16'ha00;
17'hcd1f:	data_out=16'h99b;
17'hcd20:	data_out=16'h89dd;
17'hcd21:	data_out=16'h9ff;
17'hcd22:	data_out=16'h9ea;
17'hcd23:	data_out=16'h9fe;
17'hcd24:	data_out=16'h9ff;
17'hcd25:	data_out=16'h9f3;
17'hcd26:	data_out=16'ha00;
17'hcd27:	data_out=16'h8964;
17'hcd28:	data_out=16'ha00;
17'hcd29:	data_out=16'h9f9;
17'hcd2a:	data_out=16'ha00;
17'hcd2b:	data_out=16'ha00;
17'hcd2c:	data_out=16'h8a00;
17'hcd2d:	data_out=16'h882f;
17'hcd2e:	data_out=16'ha00;
17'hcd2f:	data_out=16'h895f;
17'hcd30:	data_out=16'h82a4;
17'hcd31:	data_out=16'h89ff;
17'hcd32:	data_out=16'h89c0;
17'hcd33:	data_out=16'ha00;
17'hcd34:	data_out=16'h89ef;
17'hcd35:	data_out=16'h896b;
17'hcd36:	data_out=16'ha00;
17'hcd37:	data_out=16'ha00;
17'hcd38:	data_out=16'h8a00;
17'hcd39:	data_out=16'h9ff;
17'hcd3a:	data_out=16'h9d7;
17'hcd3b:	data_out=16'h89d4;
17'hcd3c:	data_out=16'h9fe;
17'hcd3d:	data_out=16'h89c9;
17'hcd3e:	data_out=16'ha00;
17'hcd3f:	data_out=16'h8a00;
17'hcd40:	data_out=16'h89ff;
17'hcd41:	data_out=16'h9a2;
17'hcd42:	data_out=16'h8794;
17'hcd43:	data_out=16'h9da;
17'hcd44:	data_out=16'h89f9;
17'hcd45:	data_out=16'h8a00;
17'hcd46:	data_out=16'ha00;
17'hcd47:	data_out=16'h9c6;
17'hcd48:	data_out=16'h99b;
17'hcd49:	data_out=16'h9e4;
17'hcd4a:	data_out=16'h9a4;
17'hcd4b:	data_out=16'h874c;
17'hcd4c:	data_out=16'h9e8;
17'hcd4d:	data_out=16'h9f4;
17'hcd4e:	data_out=16'ha00;
17'hcd4f:	data_out=16'h9fa;
17'hcd50:	data_out=16'h89d7;
17'hcd51:	data_out=16'h85cd;
17'hcd52:	data_out=16'h83b1;
17'hcd53:	data_out=16'ha00;
17'hcd54:	data_out=16'h88fc;
17'hcd55:	data_out=16'h9f0;
17'hcd56:	data_out=16'h9ee;
17'hcd57:	data_out=16'h9c4;
17'hcd58:	data_out=16'h9f4;
17'hcd59:	data_out=16'h89c8;
17'hcd5a:	data_out=16'ha00;
17'hcd5b:	data_out=16'h89e1;
17'hcd5c:	data_out=16'h8995;
17'hcd5d:	data_out=16'h8987;
17'hcd5e:	data_out=16'h882a;
17'hcd5f:	data_out=16'h643;
17'hcd60:	data_out=16'h9fd;
17'hcd61:	data_out=16'h89e2;
17'hcd62:	data_out=16'h9fc;
17'hcd63:	data_out=16'ha00;
17'hcd64:	data_out=16'h8a00;
17'hcd65:	data_out=16'h88c1;
17'hcd66:	data_out=16'ha00;
17'hcd67:	data_out=16'h9ff;
17'hcd68:	data_out=16'ha00;
17'hcd69:	data_out=16'h9fd;
17'hcd6a:	data_out=16'h9ff;
17'hcd6b:	data_out=16'h89ff;
17'hcd6c:	data_out=16'h89d1;
17'hcd6d:	data_out=16'ha00;
17'hcd6e:	data_out=16'h9ff;
17'hcd6f:	data_out=16'h89ff;
17'hcd70:	data_out=16'h9ff;
17'hcd71:	data_out=16'h9fd;
17'hcd72:	data_out=16'h8a00;
17'hcd73:	data_out=16'h89e8;
17'hcd74:	data_out=16'h8369;
17'hcd75:	data_out=16'h89ff;
17'hcd76:	data_out=16'ha00;
17'hcd77:	data_out=16'h9df;
17'hcd78:	data_out=16'h8385;
17'hcd79:	data_out=16'ha00;
17'hcd7a:	data_out=16'ha00;
17'hcd7b:	data_out=16'ha00;
17'hcd7c:	data_out=16'h9db;
17'hcd7d:	data_out=16'h8815;
17'hcd7e:	data_out=16'h81f7;
17'hcd7f:	data_out=16'h8a00;
17'hcd80:	data_out=16'h8a00;
17'hcd81:	data_out=16'h8a00;
17'hcd82:	data_out=16'h9e3;
17'hcd83:	data_out=16'h8948;
17'hcd84:	data_out=16'h8a00;
17'hcd85:	data_out=16'h8a00;
17'hcd86:	data_out=16'h8959;
17'hcd87:	data_out=16'ha00;
17'hcd88:	data_out=16'ha00;
17'hcd89:	data_out=16'h9da;
17'hcd8a:	data_out=16'h8a00;
17'hcd8b:	data_out=16'ha00;
17'hcd8c:	data_out=16'ha00;
17'hcd8d:	data_out=16'h89fa;
17'hcd8e:	data_out=16'h888a;
17'hcd8f:	data_out=16'ha00;
17'hcd90:	data_out=16'h953;
17'hcd91:	data_out=16'h89ff;
17'hcd92:	data_out=16'h9c4;
17'hcd93:	data_out=16'h8917;
17'hcd94:	data_out=16'h85e8;
17'hcd95:	data_out=16'h8a00;
17'hcd96:	data_out=16'h8a00;
17'hcd97:	data_out=16'h86ef;
17'hcd98:	data_out=16'h9dc;
17'hcd99:	data_out=16'ha00;
17'hcd9a:	data_out=16'h8a00;
17'hcd9b:	data_out=16'ha00;
17'hcd9c:	data_out=16'h89fb;
17'hcd9d:	data_out=16'h89f1;
17'hcd9e:	data_out=16'h865f;
17'hcd9f:	data_out=16'h89f4;
17'hcda0:	data_out=16'h89fa;
17'hcda1:	data_out=16'h8715;
17'hcda2:	data_out=16'h395;
17'hcda3:	data_out=16'ha00;
17'hcda4:	data_out=16'ha00;
17'hcda5:	data_out=16'h8309;
17'hcda6:	data_out=16'h9fd;
17'hcda7:	data_out=16'h8693;
17'hcda8:	data_out=16'h84b6;
17'hcda9:	data_out=16'h9ff;
17'hcdaa:	data_out=16'ha00;
17'hcdab:	data_out=16'ha00;
17'hcdac:	data_out=16'h8a00;
17'hcdad:	data_out=16'h89ad;
17'hcdae:	data_out=16'h9ab;
17'hcdaf:	data_out=16'h89ed;
17'hcdb0:	data_out=16'h87de;
17'hcdb1:	data_out=16'h8a00;
17'hcdb2:	data_out=16'h8a00;
17'hcdb3:	data_out=16'h81e1;
17'hcdb4:	data_out=16'h89f5;
17'hcdb5:	data_out=16'h89fc;
17'hcdb6:	data_out=16'ha00;
17'hcdb7:	data_out=16'h9f3;
17'hcdb8:	data_out=16'h8a00;
17'hcdb9:	data_out=16'h8621;
17'hcdba:	data_out=16'h9f0;
17'hcdbb:	data_out=16'h89f4;
17'hcdbc:	data_out=16'h8603;
17'hcdbd:	data_out=16'h89fa;
17'hcdbe:	data_out=16'h84af;
17'hcdbf:	data_out=16'h8a00;
17'hcdc0:	data_out=16'h8a00;
17'hcdc1:	data_out=16'h976;
17'hcdc2:	data_out=16'h8264;
17'hcdc3:	data_out=16'h8920;
17'hcdc4:	data_out=16'h89ff;
17'hcdc5:	data_out=16'h8a00;
17'hcdc6:	data_out=16'h9fa;
17'hcdc7:	data_out=16'h9f6;
17'hcdc8:	data_out=16'h988;
17'hcdc9:	data_out=16'h8737;
17'hcdca:	data_out=16'h9fa;
17'hcdcb:	data_out=16'h9a0;
17'hcdcc:	data_out=16'h82a;
17'hcdcd:	data_out=16'h9ed;
17'hcdce:	data_out=16'ha00;
17'hcdcf:	data_out=16'h9f9;
17'hcdd0:	data_out=16'h8a00;
17'hcdd1:	data_out=16'h89f6;
17'hcdd2:	data_out=16'h8118;
17'hcdd3:	data_out=16'h429;
17'hcdd4:	data_out=16'h84e8;
17'hcdd5:	data_out=16'h8111;
17'hcdd6:	data_out=16'h8689;
17'hcdd7:	data_out=16'h89b8;
17'hcdd8:	data_out=16'h882b;
17'hcdd9:	data_out=16'h8a00;
17'hcdda:	data_out=16'h9fe;
17'hcddb:	data_out=16'h8a00;
17'hcddc:	data_out=16'h8a00;
17'hcddd:	data_out=16'h89f9;
17'hcdde:	data_out=16'h89f4;
17'hcddf:	data_out=16'h6ad;
17'hcde0:	data_out=16'h856a;
17'hcde1:	data_out=16'h8a00;
17'hcde2:	data_out=16'h896;
17'hcde3:	data_out=16'h8184;
17'hcde4:	data_out=16'h89ff;
17'hcde5:	data_out=16'h89c8;
17'hcde6:	data_out=16'ha00;
17'hcde7:	data_out=16'ha00;
17'hcde8:	data_out=16'h861e;
17'hcde9:	data_out=16'ha00;
17'hcdea:	data_out=16'h8942;
17'hcdeb:	data_out=16'h8a00;
17'hcdec:	data_out=16'h8a00;
17'hcded:	data_out=16'h8218;
17'hcdee:	data_out=16'h8942;
17'hcdef:	data_out=16'h8a00;
17'hcdf0:	data_out=16'h8901;
17'hcdf1:	data_out=16'h9b9;
17'hcdf2:	data_out=16'h8a00;
17'hcdf3:	data_out=16'h8a00;
17'hcdf4:	data_out=16'h87cd;
17'hcdf5:	data_out=16'h8a00;
17'hcdf6:	data_out=16'ha00;
17'hcdf7:	data_out=16'h9c1;
17'hcdf8:	data_out=16'h89fd;
17'hcdf9:	data_out=16'h9fd;
17'hcdfa:	data_out=16'h841d;
17'hcdfb:	data_out=16'h84ab;
17'hcdfc:	data_out=16'h9c7;
17'hcdfd:	data_out=16'h89f3;
17'hcdfe:	data_out=16'h8a00;
17'hcdff:	data_out=16'h8a00;
17'hce00:	data_out=16'h89fd;
17'hce01:	data_out=16'h8a00;
17'hce02:	data_out=16'h8813;
17'hce03:	data_out=16'h8937;
17'hce04:	data_out=16'h8a00;
17'hce05:	data_out=16'h8a00;
17'hce06:	data_out=16'h89fb;
17'hce07:	data_out=16'ha00;
17'hce08:	data_out=16'h9c4;
17'hce09:	data_out=16'h9ef;
17'hce0a:	data_out=16'h8a00;
17'hce0b:	data_out=16'ha00;
17'hce0c:	data_out=16'ha00;
17'hce0d:	data_out=16'h89c5;
17'hce0e:	data_out=16'h89ff;
17'hce0f:	data_out=16'h2d3;
17'hce10:	data_out=16'h95b;
17'hce11:	data_out=16'h8a00;
17'hce12:	data_out=16'h814e;
17'hce13:	data_out=16'h8718;
17'hce14:	data_out=16'h8975;
17'hce15:	data_out=16'h89ff;
17'hce16:	data_out=16'h89fd;
17'hce17:	data_out=16'h8900;
17'hce18:	data_out=16'h89fb;
17'hce19:	data_out=16'ha00;
17'hce1a:	data_out=16'h8a00;
17'hce1b:	data_out=16'h8192;
17'hce1c:	data_out=16'h89ff;
17'hce1d:	data_out=16'h89f1;
17'hce1e:	data_out=16'h89dc;
17'hce1f:	data_out=16'h89f8;
17'hce20:	data_out=16'h89f8;
17'hce21:	data_out=16'h89ff;
17'hce22:	data_out=16'h86ca;
17'hce23:	data_out=16'ha00;
17'hce24:	data_out=16'ha00;
17'hce25:	data_out=16'h89e9;
17'hce26:	data_out=16'h9ed;
17'hce27:	data_out=16'h89fc;
17'hce28:	data_out=16'h89ff;
17'hce29:	data_out=16'h83a1;
17'hce2a:	data_out=16'h9e3;
17'hce2b:	data_out=16'ha00;
17'hce2c:	data_out=16'h89fe;
17'hce2d:	data_out=16'h851c;
17'hce2e:	data_out=16'h8806;
17'hce2f:	data_out=16'h89f4;
17'hce30:	data_out=16'h89d8;
17'hce31:	data_out=16'h8a00;
17'hce32:	data_out=16'h8a00;
17'hce33:	data_out=16'h89f1;
17'hce34:	data_out=16'h89e5;
17'hce35:	data_out=16'h89ff;
17'hce36:	data_out=16'h9b8;
17'hce37:	data_out=16'h870a;
17'hce38:	data_out=16'h8a00;
17'hce39:	data_out=16'h89f1;
17'hce3a:	data_out=16'h9f3;
17'hce3b:	data_out=16'h89dc;
17'hce3c:	data_out=16'h8940;
17'hce3d:	data_out=16'h89f5;
17'hce3e:	data_out=16'h89ff;
17'hce3f:	data_out=16'h8a00;
17'hce40:	data_out=16'h8a00;
17'hce41:	data_out=16'h810b;
17'hce42:	data_out=16'h9fa;
17'hce43:	data_out=16'h89ca;
17'hce44:	data_out=16'h89ff;
17'hce45:	data_out=16'h89ff;
17'hce46:	data_out=16'h6d5;
17'hce47:	data_out=16'ha00;
17'hce48:	data_out=16'h8710;
17'hce49:	data_out=16'h89c0;
17'hce4a:	data_out=16'ha00;
17'hce4b:	data_out=16'h9f4;
17'hce4c:	data_out=16'h8b2;
17'hce4d:	data_out=16'h17;
17'hce4e:	data_out=16'h70c;
17'hce4f:	data_out=16'h9f0;
17'hce50:	data_out=16'h89fc;
17'hce51:	data_out=16'h89f8;
17'hce52:	data_out=16'h11a;
17'hce53:	data_out=16'h84ca;
17'hce54:	data_out=16'h87e4;
17'hce55:	data_out=16'h88b6;
17'hce56:	data_out=16'h8945;
17'hce57:	data_out=16'h89f2;
17'hce58:	data_out=16'h89f6;
17'hce59:	data_out=16'h89fd;
17'hce5a:	data_out=16'h884c;
17'hce5b:	data_out=16'h8a00;
17'hce5c:	data_out=16'h8a00;
17'hce5d:	data_out=16'h89f8;
17'hce5e:	data_out=16'h89fa;
17'hce5f:	data_out=16'h882d;
17'hce60:	data_out=16'h85f3;
17'hce61:	data_out=16'h8a00;
17'hce62:	data_out=16'h80eb;
17'hce63:	data_out=16'h89de;
17'hce64:	data_out=16'h86c1;
17'hce65:	data_out=16'h89c4;
17'hce66:	data_out=16'ha00;
17'hce67:	data_out=16'ha00;
17'hce68:	data_out=16'h89ff;
17'hce69:	data_out=16'h9e5;
17'hce6a:	data_out=16'h89ff;
17'hce6b:	data_out=16'h8a00;
17'hce6c:	data_out=16'h89ff;
17'hce6d:	data_out=16'h89e3;
17'hce6e:	data_out=16'h89ff;
17'hce6f:	data_out=16'h8a00;
17'hce70:	data_out=16'h89ff;
17'hce71:	data_out=16'h8453;
17'hce72:	data_out=16'h8a00;
17'hce73:	data_out=16'h8a00;
17'hce74:	data_out=16'h89da;
17'hce75:	data_out=16'h8a00;
17'hce76:	data_out=16'ha00;
17'hce77:	data_out=16'h544;
17'hce78:	data_out=16'h89fa;
17'hce79:	data_out=16'h392;
17'hce7a:	data_out=16'h899e;
17'hce7b:	data_out=16'h89ff;
17'hce7c:	data_out=16'h89fd;
17'hce7d:	data_out=16'h89f8;
17'hce7e:	data_out=16'h8a00;
17'hce7f:	data_out=16'h8a00;
17'hce80:	data_out=16'h89fb;
17'hce81:	data_out=16'h8a00;
17'hce82:	data_out=16'h89f5;
17'hce83:	data_out=16'h883e;
17'hce84:	data_out=16'h89fc;
17'hce85:	data_out=16'h8a00;
17'hce86:	data_out=16'h89da;
17'hce87:	data_out=16'ha00;
17'hce88:	data_out=16'h98f;
17'hce89:	data_out=16'ha00;
17'hce8a:	data_out=16'h8a00;
17'hce8b:	data_out=16'ha00;
17'hce8c:	data_out=16'ha00;
17'hce8d:	data_out=16'h89f4;
17'hce8e:	data_out=16'h8a00;
17'hce8f:	data_out=16'h81d2;
17'hce90:	data_out=16'h757;
17'hce91:	data_out=16'h8a00;
17'hce92:	data_out=16'h89f4;
17'hce93:	data_out=16'h84a8;
17'hce94:	data_out=16'h89e4;
17'hce95:	data_out=16'h8a00;
17'hce96:	data_out=16'h89fc;
17'hce97:	data_out=16'h87d4;
17'hce98:	data_out=16'h89ff;
17'hce99:	data_out=16'ha00;
17'hce9a:	data_out=16'h8a00;
17'hce9b:	data_out=16'h86f9;
17'hce9c:	data_out=16'h8a00;
17'hce9d:	data_out=16'h89e8;
17'hce9e:	data_out=16'h89f9;
17'hce9f:	data_out=16'h89fe;
17'hcea0:	data_out=16'h89fe;
17'hcea1:	data_out=16'h8a00;
17'hcea2:	data_out=16'h5e6;
17'hcea3:	data_out=16'h9fd;
17'hcea4:	data_out=16'h9fd;
17'hcea5:	data_out=16'h853d;
17'hcea6:	data_out=16'h9ff;
17'hcea7:	data_out=16'h89fc;
17'hcea8:	data_out=16'h8a00;
17'hcea9:	data_out=16'h874e;
17'hceaa:	data_out=16'ha00;
17'hceab:	data_out=16'ha00;
17'hceac:	data_out=16'h89fe;
17'hcead:	data_out=16'ha00;
17'hceae:	data_out=16'h165;
17'hceaf:	data_out=16'h89fb;
17'hceb0:	data_out=16'h89e7;
17'hceb1:	data_out=16'h8a00;
17'hceb2:	data_out=16'h8985;
17'hceb3:	data_out=16'h89ff;
17'hceb4:	data_out=16'h89dc;
17'hceb5:	data_out=16'h8a00;
17'hceb6:	data_out=16'h821c;
17'hceb7:	data_out=16'h89d5;
17'hceb8:	data_out=16'h8a00;
17'hceb9:	data_out=16'h89ff;
17'hceba:	data_out=16'ha00;
17'hcebb:	data_out=16'h82e8;
17'hcebc:	data_out=16'h89ff;
17'hcebd:	data_out=16'h89fd;
17'hcebe:	data_out=16'h8a00;
17'hcebf:	data_out=16'h8a00;
17'hcec0:	data_out=16'h89f9;
17'hcec1:	data_out=16'h884c;
17'hcec2:	data_out=16'ha00;
17'hcec3:	data_out=16'h8318;
17'hcec4:	data_out=16'h8a00;
17'hcec5:	data_out=16'h8a00;
17'hcec6:	data_out=16'h896d;
17'hcec7:	data_out=16'ha00;
17'hcec8:	data_out=16'h9df;
17'hcec9:	data_out=16'h89c7;
17'hceca:	data_out=16'ha00;
17'hcecb:	data_out=16'ha00;
17'hcecc:	data_out=16'h9dc;
17'hcecd:	data_out=16'h230;
17'hcece:	data_out=16'ha00;
17'hcecf:	data_out=16'h9fe;
17'hced0:	data_out=16'h89e2;
17'hced1:	data_out=16'h8a00;
17'hced2:	data_out=16'h4e0;
17'hced3:	data_out=16'h886c;
17'hced4:	data_out=16'h89fa;
17'hced5:	data_out=16'h893d;
17'hced6:	data_out=16'h89fc;
17'hced7:	data_out=16'h8a00;
17'hced8:	data_out=16'h8a00;
17'hced9:	data_out=16'h89fb;
17'hceda:	data_out=16'h89d6;
17'hcedb:	data_out=16'h8a00;
17'hcedc:	data_out=16'h8a00;
17'hcedd:	data_out=16'h89fa;
17'hcede:	data_out=16'h8836;
17'hcedf:	data_out=16'h89fe;
17'hcee0:	data_out=16'h9fd;
17'hcee1:	data_out=16'h8a00;
17'hcee2:	data_out=16'ha00;
17'hcee3:	data_out=16'h89fa;
17'hcee4:	data_out=16'h86b8;
17'hcee5:	data_out=16'h820d;
17'hcee6:	data_out=16'ha00;
17'hcee7:	data_out=16'ha00;
17'hcee8:	data_out=16'h8a00;
17'hcee9:	data_out=16'h9b9;
17'hceea:	data_out=16'h8a00;
17'hceeb:	data_out=16'h8a00;
17'hceec:	data_out=16'h89fc;
17'hceed:	data_out=16'h89fc;
17'hceee:	data_out=16'h8a00;
17'hceef:	data_out=16'h8988;
17'hcef0:	data_out=16'h8a00;
17'hcef1:	data_out=16'h848b;
17'hcef2:	data_out=16'h8a00;
17'hcef3:	data_out=16'h8a00;
17'hcef4:	data_out=16'h89ee;
17'hcef5:	data_out=16'h8a00;
17'hcef6:	data_out=16'ha00;
17'hcef7:	data_out=16'h462;
17'hcef8:	data_out=16'h33b;
17'hcef9:	data_out=16'h876b;
17'hcefa:	data_out=16'h89ee;
17'hcefb:	data_out=16'h8a00;
17'hcefc:	data_out=16'h8a00;
17'hcefd:	data_out=16'h8a00;
17'hcefe:	data_out=16'h7e;
17'hceff:	data_out=16'h8a00;
17'hcf00:	data_out=16'h89fd;
17'hcf01:	data_out=16'h8a00;
17'hcf02:	data_out=16'h89f4;
17'hcf03:	data_out=16'h87fc;
17'hcf04:	data_out=16'h89fc;
17'hcf05:	data_out=16'h8a00;
17'hcf06:	data_out=16'h80c;
17'hcf07:	data_out=16'ha00;
17'hcf08:	data_out=16'h8568;
17'hcf09:	data_out=16'ha00;
17'hcf0a:	data_out=16'h8a00;
17'hcf0b:	data_out=16'ha00;
17'hcf0c:	data_out=16'ha00;
17'hcf0d:	data_out=16'h89e7;
17'hcf0e:	data_out=16'h8a00;
17'hcf0f:	data_out=16'h8069;
17'hcf10:	data_out=16'h882;
17'hcf11:	data_out=16'h8a00;
17'hcf12:	data_out=16'h276;
17'hcf13:	data_out=16'h9f2;
17'hcf14:	data_out=16'h89f2;
17'hcf15:	data_out=16'h8a00;
17'hcf16:	data_out=16'h89f9;
17'hcf17:	data_out=16'hcc;
17'hcf18:	data_out=16'h8a00;
17'hcf19:	data_out=16'ha00;
17'hcf1a:	data_out=16'h8a00;
17'hcf1b:	data_out=16'h89e7;
17'hcf1c:	data_out=16'h8a00;
17'hcf1d:	data_out=16'h89df;
17'hcf1e:	data_out=16'h89f9;
17'hcf1f:	data_out=16'h89f6;
17'hcf20:	data_out=16'h8a00;
17'hcf21:	data_out=16'h8a00;
17'hcf22:	data_out=16'h9d6;
17'hcf23:	data_out=16'h98f;
17'hcf24:	data_out=16'h993;
17'hcf25:	data_out=16'h463;
17'hcf26:	data_out=16'ha00;
17'hcf27:	data_out=16'h89fd;
17'hcf28:	data_out=16'h8a00;
17'hcf29:	data_out=16'h8387;
17'hcf2a:	data_out=16'ha00;
17'hcf2b:	data_out=16'ha00;
17'hcf2c:	data_out=16'h89fe;
17'hcf2d:	data_out=16'ha00;
17'hcf2e:	data_out=16'ha00;
17'hcf2f:	data_out=16'h89f7;
17'hcf30:	data_out=16'h66b;
17'hcf31:	data_out=16'h8a00;
17'hcf32:	data_out=16'h7d6;
17'hcf33:	data_out=16'h8a00;
17'hcf34:	data_out=16'h85a0;
17'hcf35:	data_out=16'h89ff;
17'hcf36:	data_out=16'h8955;
17'hcf37:	data_out=16'h89ed;
17'hcf38:	data_out=16'h8a00;
17'hcf39:	data_out=16'h8a00;
17'hcf3a:	data_out=16'ha00;
17'hcf3b:	data_out=16'h809;
17'hcf3c:	data_out=16'h8a00;
17'hcf3d:	data_out=16'h8a00;
17'hcf3e:	data_out=16'h8a00;
17'hcf3f:	data_out=16'h8a00;
17'hcf40:	data_out=16'h89ea;
17'hcf41:	data_out=16'h89fb;
17'hcf42:	data_out=16'ha00;
17'hcf43:	data_out=16'h166;
17'hcf44:	data_out=16'h8a00;
17'hcf45:	data_out=16'h8a00;
17'hcf46:	data_out=16'h89ff;
17'hcf47:	data_out=16'ha00;
17'hcf48:	data_out=16'ha00;
17'hcf49:	data_out=16'h8204;
17'hcf4a:	data_out=16'ha00;
17'hcf4b:	data_out=16'ha00;
17'hcf4c:	data_out=16'h9f9;
17'hcf4d:	data_out=16'h793;
17'hcf4e:	data_out=16'h9f3;
17'hcf4f:	data_out=16'ha00;
17'hcf50:	data_out=16'h89e2;
17'hcf51:	data_out=16'h89ff;
17'hcf52:	data_out=16'h904;
17'hcf53:	data_out=16'h89f6;
17'hcf54:	data_out=16'h89ff;
17'hcf55:	data_out=16'h89d8;
17'hcf56:	data_out=16'h89fe;
17'hcf57:	data_out=16'h8a00;
17'hcf58:	data_out=16'h8a00;
17'hcf59:	data_out=16'h89ff;
17'hcf5a:	data_out=16'h89e6;
17'hcf5b:	data_out=16'h89ff;
17'hcf5c:	data_out=16'h8a00;
17'hcf5d:	data_out=16'h89fb;
17'hcf5e:	data_out=16'h8872;
17'hcf5f:	data_out=16'h89fd;
17'hcf60:	data_out=16'ha00;
17'hcf61:	data_out=16'h8a00;
17'hcf62:	data_out=16'ha00;
17'hcf63:	data_out=16'h89fa;
17'hcf64:	data_out=16'h838f;
17'hcf65:	data_out=16'h99c;
17'hcf66:	data_out=16'ha00;
17'hcf67:	data_out=16'ha00;
17'hcf68:	data_out=16'h8a00;
17'hcf69:	data_out=16'h9b7;
17'hcf6a:	data_out=16'h8a00;
17'hcf6b:	data_out=16'h8a00;
17'hcf6c:	data_out=16'h89fd;
17'hcf6d:	data_out=16'h89fc;
17'hcf6e:	data_out=16'h8a00;
17'hcf6f:	data_out=16'h9fa;
17'hcf70:	data_out=16'h8a00;
17'hcf71:	data_out=16'h806f;
17'hcf72:	data_out=16'h8a00;
17'hcf73:	data_out=16'h8a00;
17'hcf74:	data_out=16'h5ed;
17'hcf75:	data_out=16'h8a00;
17'hcf76:	data_out=16'ha00;
17'hcf77:	data_out=16'ha00;
17'hcf78:	data_out=16'h9ea;
17'hcf79:	data_out=16'h82bf;
17'hcf7a:	data_out=16'h89f3;
17'hcf7b:	data_out=16'h8a00;
17'hcf7c:	data_out=16'h8a00;
17'hcf7d:	data_out=16'h8a00;
17'hcf7e:	data_out=16'h7bf;
17'hcf7f:	data_out=16'h8a00;
17'hcf80:	data_out=16'h89ff;
17'hcf81:	data_out=16'h8a00;
17'hcf82:	data_out=16'h8a00;
17'hcf83:	data_out=16'h89ab;
17'hcf84:	data_out=16'h840f;
17'hcf85:	data_out=16'h8a00;
17'hcf86:	data_out=16'h9a5;
17'hcf87:	data_out=16'ha00;
17'hcf88:	data_out=16'h8a00;
17'hcf89:	data_out=16'ha00;
17'hcf8a:	data_out=16'h8a00;
17'hcf8b:	data_out=16'ha00;
17'hcf8c:	data_out=16'ha00;
17'hcf8d:	data_out=16'h8a00;
17'hcf8e:	data_out=16'h8a00;
17'hcf8f:	data_out=16'h8423;
17'hcf90:	data_out=16'h395;
17'hcf91:	data_out=16'h89ff;
17'hcf92:	data_out=16'h3e6;
17'hcf93:	data_out=16'h97f;
17'hcf94:	data_out=16'h89f8;
17'hcf95:	data_out=16'h8a00;
17'hcf96:	data_out=16'h89fe;
17'hcf97:	data_out=16'h810f;
17'hcf98:	data_out=16'h8a00;
17'hcf99:	data_out=16'ha00;
17'hcf9a:	data_out=16'h89b5;
17'hcf9b:	data_out=16'h8a00;
17'hcf9c:	data_out=16'h8a00;
17'hcf9d:	data_out=16'h894e;
17'hcf9e:	data_out=16'h8a00;
17'hcf9f:	data_out=16'h89f0;
17'hcfa0:	data_out=16'h8a00;
17'hcfa1:	data_out=16'h8a00;
17'hcfa2:	data_out=16'h9e2;
17'hcfa3:	data_out=16'h755;
17'hcfa4:	data_out=16'h747;
17'hcfa5:	data_out=16'h67c;
17'hcfa6:	data_out=16'h9e3;
17'hcfa7:	data_out=16'h89fd;
17'hcfa8:	data_out=16'h8a00;
17'hcfa9:	data_out=16'h8a00;
17'hcfaa:	data_out=16'ha00;
17'hcfab:	data_out=16'ha00;
17'hcfac:	data_out=16'h89ff;
17'hcfad:	data_out=16'ha00;
17'hcfae:	data_out=16'ha00;
17'hcfaf:	data_out=16'h89fc;
17'hcfb0:	data_out=16'h951;
17'hcfb1:	data_out=16'h8a00;
17'hcfb2:	data_out=16'h9fc;
17'hcfb3:	data_out=16'h8a00;
17'hcfb4:	data_out=16'h9aa;
17'hcfb5:	data_out=16'h89ff;
17'hcfb6:	data_out=16'h8a00;
17'hcfb7:	data_out=16'h8a00;
17'hcfb8:	data_out=16'h8a00;
17'hcfb9:	data_out=16'h8a00;
17'hcfba:	data_out=16'ha00;
17'hcfbb:	data_out=16'h8a4;
17'hcfbc:	data_out=16'h8a00;
17'hcfbd:	data_out=16'h8a00;
17'hcfbe:	data_out=16'h8a00;
17'hcfbf:	data_out=16'h8a00;
17'hcfc0:	data_out=16'h9b3;
17'hcfc1:	data_out=16'h8a00;
17'hcfc2:	data_out=16'ha00;
17'hcfc3:	data_out=16'h4bf;
17'hcfc4:	data_out=16'h8a00;
17'hcfc5:	data_out=16'h8a00;
17'hcfc6:	data_out=16'h8a00;
17'hcfc7:	data_out=16'ha00;
17'hcfc8:	data_out=16'ha00;
17'hcfc9:	data_out=16'h189;
17'hcfca:	data_out=16'ha00;
17'hcfcb:	data_out=16'ha00;
17'hcfcc:	data_out=16'h9fe;
17'hcfcd:	data_out=16'h7f2;
17'hcfce:	data_out=16'h9e5;
17'hcfcf:	data_out=16'ha00;
17'hcfd0:	data_out=16'h899f;
17'hcfd1:	data_out=16'h8a00;
17'hcfd2:	data_out=16'h939;
17'hcfd3:	data_out=16'h89ff;
17'hcfd4:	data_out=16'h8a00;
17'hcfd5:	data_out=16'h89f7;
17'hcfd6:	data_out=16'h8a00;
17'hcfd7:	data_out=16'h8a00;
17'hcfd8:	data_out=16'h8a00;
17'hcfd9:	data_out=16'h89d5;
17'hcfda:	data_out=16'h8a00;
17'hcfdb:	data_out=16'h8a00;
17'hcfdc:	data_out=16'h8a00;
17'hcfdd:	data_out=16'h89f0;
17'hcfde:	data_out=16'h8740;
17'hcfdf:	data_out=16'h8a00;
17'hcfe0:	data_out=16'h9ff;
17'hcfe1:	data_out=16'h8a00;
17'hcfe2:	data_out=16'ha00;
17'hcfe3:	data_out=16'h8a00;
17'hcfe4:	data_out=16'h9c5;
17'hcfe5:	data_out=16'ha00;
17'hcfe6:	data_out=16'ha00;
17'hcfe7:	data_out=16'ha00;
17'hcfe8:	data_out=16'h8a00;
17'hcfe9:	data_out=16'h8626;
17'hcfea:	data_out=16'h8a00;
17'hcfeb:	data_out=16'h8a00;
17'hcfec:	data_out=16'h89ff;
17'hcfed:	data_out=16'h8a00;
17'hcfee:	data_out=16'h8a00;
17'hcfef:	data_out=16'h9fd;
17'hcff0:	data_out=16'h8a00;
17'hcff1:	data_out=16'h823b;
17'hcff2:	data_out=16'h8a00;
17'hcff3:	data_out=16'h89ff;
17'hcff4:	data_out=16'h8e5;
17'hcff5:	data_out=16'h8a00;
17'hcff6:	data_out=16'ha00;
17'hcff7:	data_out=16'h477;
17'hcff8:	data_out=16'h9fc;
17'hcff9:	data_out=16'h82c7;
17'hcffa:	data_out=16'h89fc;
17'hcffb:	data_out=16'h8a00;
17'hcffc:	data_out=16'h8a00;
17'hcffd:	data_out=16'h8a00;
17'hcffe:	data_out=16'h928;
17'hcfff:	data_out=16'h8a00;
17'hd000:	data_out=16'h89fe;
17'hd001:	data_out=16'h8644;
17'hd002:	data_out=16'h8a00;
17'hd003:	data_out=16'h89ee;
17'hd004:	data_out=16'h9fb;
17'hd005:	data_out=16'h89fd;
17'hd006:	data_out=16'h9e1;
17'hd007:	data_out=16'ha00;
17'hd008:	data_out=16'h8a00;
17'hd009:	data_out=16'ha00;
17'hd00a:	data_out=16'h38e;
17'hd00b:	data_out=16'ha00;
17'hd00c:	data_out=16'ha00;
17'hd00d:	data_out=16'h8a00;
17'hd00e:	data_out=16'h8a00;
17'hd00f:	data_out=16'h89dc;
17'hd010:	data_out=16'h6c0;
17'hd011:	data_out=16'h9ed;
17'hd012:	data_out=16'h182;
17'hd013:	data_out=16'h503;
17'hd014:	data_out=16'h89f8;
17'hd015:	data_out=16'h8a00;
17'hd016:	data_out=16'h89fe;
17'hd017:	data_out=16'h89e5;
17'hd018:	data_out=16'h8a00;
17'hd019:	data_out=16'ha00;
17'hd01a:	data_out=16'h8d3;
17'hd01b:	data_out=16'h8a00;
17'hd01c:	data_out=16'h8a00;
17'hd01d:	data_out=16'h1fe;
17'hd01e:	data_out=16'h89fd;
17'hd01f:	data_out=16'h89ee;
17'hd020:	data_out=16'h8a00;
17'hd021:	data_out=16'h8a00;
17'hd022:	data_out=16'h9fe;
17'hd023:	data_out=16'h10a;
17'hd024:	data_out=16'hf6;
17'hd025:	data_out=16'h8aa;
17'hd026:	data_out=16'h9d9;
17'hd027:	data_out=16'h85a7;
17'hd028:	data_out=16'h8a00;
17'hd029:	data_out=16'h8a00;
17'hd02a:	data_out=16'h829b;
17'hd02b:	data_out=16'ha00;
17'hd02c:	data_out=16'h8a00;
17'hd02d:	data_out=16'ha00;
17'hd02e:	data_out=16'h83bf;
17'hd02f:	data_out=16'h894a;
17'hd030:	data_out=16'h951;
17'hd031:	data_out=16'h744;
17'hd032:	data_out=16'h9db;
17'hd033:	data_out=16'h8a00;
17'hd034:	data_out=16'h9e3;
17'hd035:	data_out=16'h59b;
17'hd036:	data_out=16'h8a00;
17'hd037:	data_out=16'h8a00;
17'hd038:	data_out=16'h632;
17'hd039:	data_out=16'h8a00;
17'hd03a:	data_out=16'ha00;
17'hd03b:	data_out=16'h878;
17'hd03c:	data_out=16'h8a00;
17'hd03d:	data_out=16'h8a00;
17'hd03e:	data_out=16'h8a00;
17'hd03f:	data_out=16'h89fe;
17'hd040:	data_out=16'h9ff;
17'hd041:	data_out=16'h8a00;
17'hd042:	data_out=16'ha00;
17'hd043:	data_out=16'h8193;
17'hd044:	data_out=16'h89ff;
17'hd045:	data_out=16'h8a00;
17'hd046:	data_out=16'h8a00;
17'hd047:	data_out=16'ha00;
17'hd048:	data_out=16'ha00;
17'hd049:	data_out=16'h74b;
17'hd04a:	data_out=16'ha00;
17'hd04b:	data_out=16'ha00;
17'hd04c:	data_out=16'h9ff;
17'hd04d:	data_out=16'h9c4;
17'hd04e:	data_out=16'h8066;
17'hd04f:	data_out=16'ha00;
17'hd050:	data_out=16'h89ba;
17'hd051:	data_out=16'h8a00;
17'hd052:	data_out=16'h318;
17'hd053:	data_out=16'h89f4;
17'hd054:	data_out=16'h89f8;
17'hd055:	data_out=16'h89fe;
17'hd056:	data_out=16'h8a00;
17'hd057:	data_out=16'h8a00;
17'hd058:	data_out=16'h8a00;
17'hd059:	data_out=16'ha00;
17'hd05a:	data_out=16'h8a00;
17'hd05b:	data_out=16'h89fd;
17'hd05c:	data_out=16'h8a00;
17'hd05d:	data_out=16'h8985;
17'hd05e:	data_out=16'h107;
17'hd05f:	data_out=16'h89d7;
17'hd060:	data_out=16'h9f7;
17'hd061:	data_out=16'h8a00;
17'hd062:	data_out=16'h810d;
17'hd063:	data_out=16'h89fb;
17'hd064:	data_out=16'h9ec;
17'hd065:	data_out=16'ha00;
17'hd066:	data_out=16'h9ff;
17'hd067:	data_out=16'ha00;
17'hd068:	data_out=16'h8a00;
17'hd069:	data_out=16'h8a00;
17'hd06a:	data_out=16'h8a00;
17'hd06b:	data_out=16'h81ba;
17'hd06c:	data_out=16'h85c8;
17'hd06d:	data_out=16'h89fc;
17'hd06e:	data_out=16'h8a00;
17'hd06f:	data_out=16'h9fd;
17'hd070:	data_out=16'h8a00;
17'hd071:	data_out=16'h89dc;
17'hd072:	data_out=16'h8840;
17'hd073:	data_out=16'h8229;
17'hd074:	data_out=16'h8cf;
17'hd075:	data_out=16'h8a00;
17'hd076:	data_out=16'ha00;
17'hd077:	data_out=16'h85e2;
17'hd078:	data_out=16'h490;
17'hd079:	data_out=16'h8a00;
17'hd07a:	data_out=16'h89f7;
17'hd07b:	data_out=16'h8a00;
17'hd07c:	data_out=16'h8a00;
17'hd07d:	data_out=16'h8930;
17'hd07e:	data_out=16'h9dc;
17'hd07f:	data_out=16'h8a00;
17'hd080:	data_out=16'h9fa;
17'hd081:	data_out=16'h9fa;
17'hd082:	data_out=16'h8a00;
17'hd083:	data_out=16'h89fe;
17'hd084:	data_out=16'ha00;
17'hd085:	data_out=16'h44d;
17'hd086:	data_out=16'h882a;
17'hd087:	data_out=16'h8217;
17'hd088:	data_out=16'h8a00;
17'hd089:	data_out=16'h9fd;
17'hd08a:	data_out=16'h991;
17'hd08b:	data_out=16'h8514;
17'hd08c:	data_out=16'h8a00;
17'hd08d:	data_out=16'h8a00;
17'hd08e:	data_out=16'h8602;
17'hd08f:	data_out=16'h89fc;
17'hd090:	data_out=16'hbd;
17'hd091:	data_out=16'ha00;
17'hd092:	data_out=16'h89ff;
17'hd093:	data_out=16'h89fc;
17'hd094:	data_out=16'h89fc;
17'hd095:	data_out=16'h8009;
17'hd096:	data_out=16'h89ff;
17'hd097:	data_out=16'h89fd;
17'hd098:	data_out=16'h88cb;
17'hd099:	data_out=16'ha00;
17'hd09a:	data_out=16'h9ff;
17'hd09b:	data_out=16'h8a00;
17'hd09c:	data_out=16'h6f5;
17'hd09d:	data_out=16'ha00;
17'hd09e:	data_out=16'h89fa;
17'hd09f:	data_out=16'h86cb;
17'hd0a0:	data_out=16'ha00;
17'hd0a1:	data_out=16'h861a;
17'hd0a2:	data_out=16'ha00;
17'hd0a3:	data_out=16'h8a00;
17'hd0a4:	data_out=16'h8a00;
17'hd0a5:	data_out=16'h841;
17'hd0a6:	data_out=16'h89fe;
17'hd0a7:	data_out=16'h9ff;
17'hd0a8:	data_out=16'h865d;
17'hd0a9:	data_out=16'h8a00;
17'hd0aa:	data_out=16'h89f9;
17'hd0ab:	data_out=16'ha00;
17'hd0ac:	data_out=16'h89fe;
17'hd0ad:	data_out=16'h5ec;
17'hd0ae:	data_out=16'h89f9;
17'hd0af:	data_out=16'h9f6;
17'hd0b0:	data_out=16'h8a00;
17'hd0b1:	data_out=16'h9fa;
17'hd0b2:	data_out=16'h89fe;
17'hd0b3:	data_out=16'h893d;
17'hd0b4:	data_out=16'ha00;
17'hd0b5:	data_out=16'h859b;
17'hd0b6:	data_out=16'h89fc;
17'hd0b7:	data_out=16'h8a00;
17'hd0b8:	data_out=16'ha00;
17'hd0b9:	data_out=16'h8869;
17'hd0ba:	data_out=16'h9f9;
17'hd0bb:	data_out=16'h8475;
17'hd0bc:	data_out=16'h89f9;
17'hd0bd:	data_out=16'ha00;
17'hd0be:	data_out=16'h8662;
17'hd0bf:	data_out=16'h447;
17'hd0c0:	data_out=16'ha00;
17'hd0c1:	data_out=16'h8a00;
17'hd0c2:	data_out=16'h9f7;
17'hd0c3:	data_out=16'h89fe;
17'hd0c4:	data_out=16'ha00;
17'hd0c5:	data_out=16'h808a;
17'hd0c6:	data_out=16'h89fe;
17'hd0c7:	data_out=16'h9fd;
17'hd0c8:	data_out=16'h80f7;
17'hd0c9:	data_out=16'h7bf;
17'hd0ca:	data_out=16'h84ea;
17'hd0cb:	data_out=16'h86b6;
17'hd0cc:	data_out=16'ha00;
17'hd0cd:	data_out=16'ha00;
17'hd0ce:	data_out=16'h89fe;
17'hd0cf:	data_out=16'ha00;
17'hd0d0:	data_out=16'h240;
17'hd0d1:	data_out=16'h8a00;
17'hd0d2:	data_out=16'h8a00;
17'hd0d3:	data_out=16'h31b;
17'hd0d4:	data_out=16'ha00;
17'hd0d5:	data_out=16'h8a00;
17'hd0d6:	data_out=16'h81fe;
17'hd0d7:	data_out=16'h470;
17'hd0d8:	data_out=16'h8a00;
17'hd0d9:	data_out=16'ha00;
17'hd0da:	data_out=16'h8a00;
17'hd0db:	data_out=16'h74;
17'hd0dc:	data_out=16'h67b;
17'hd0dd:	data_out=16'h8729;
17'hd0de:	data_out=16'h9f1;
17'hd0df:	data_out=16'h1a9;
17'hd0e0:	data_out=16'h8a00;
17'hd0e1:	data_out=16'h947;
17'hd0e2:	data_out=16'h89f9;
17'hd0e3:	data_out=16'h89e3;
17'hd0e4:	data_out=16'ha00;
17'hd0e5:	data_out=16'ha00;
17'hd0e6:	data_out=16'h9fd;
17'hd0e7:	data_out=16'h117;
17'hd0e8:	data_out=16'h8628;
17'hd0e9:	data_out=16'h8a00;
17'hd0ea:	data_out=16'h85f1;
17'hd0eb:	data_out=16'ha00;
17'hd0ec:	data_out=16'h378;
17'hd0ed:	data_out=16'h8983;
17'hd0ee:	data_out=16'h85f2;
17'hd0ef:	data_out=16'h83ca;
17'hd0f0:	data_out=16'h8601;
17'hd0f1:	data_out=16'h89fd;
17'hd0f2:	data_out=16'ha00;
17'hd0f3:	data_out=16'ha00;
17'hd0f4:	data_out=16'h8a00;
17'hd0f5:	data_out=16'h8a00;
17'hd0f6:	data_out=16'ha00;
17'hd0f7:	data_out=16'h837e;
17'hd0f8:	data_out=16'h89f9;
17'hd0f9:	data_out=16'h8a00;
17'hd0fa:	data_out=16'h89fb;
17'hd0fb:	data_out=16'h8664;
17'hd0fc:	data_out=16'h839b;
17'hd0fd:	data_out=16'h8733;
17'hd0fe:	data_out=16'h76c;
17'hd0ff:	data_out=16'h9ff;
17'hd100:	data_out=16'ha00;
17'hd101:	data_out=16'ha00;
17'hd102:	data_out=16'h898c;
17'hd103:	data_out=16'h57a;
17'hd104:	data_out=16'h9eb;
17'hd105:	data_out=16'h90d;
17'hd106:	data_out=16'h813b;
17'hd107:	data_out=16'h83f8;
17'hd108:	data_out=16'h89e4;
17'hd109:	data_out=16'h6eb;
17'hd10a:	data_out=16'ha00;
17'hd10b:	data_out=16'h88a3;
17'hd10c:	data_out=16'h8a00;
17'hd10d:	data_out=16'h86db;
17'hd10e:	data_out=16'h8170;
17'hd10f:	data_out=16'h89cd;
17'hd110:	data_out=16'h397;
17'hd111:	data_out=16'ha00;
17'hd112:	data_out=16'h8644;
17'hd113:	data_out=16'h80a2;
17'hd114:	data_out=16'h39a;
17'hd115:	data_out=16'h56c;
17'hd116:	data_out=16'h8071;
17'hd117:	data_out=16'h81c6;
17'hd118:	data_out=16'h815a;
17'hd119:	data_out=16'h72b;
17'hd11a:	data_out=16'h65d;
17'hd11b:	data_out=16'h81f6;
17'hd11c:	data_out=16'h9f9;
17'hd11d:	data_out=16'ha00;
17'hd11e:	data_out=16'h2ee;
17'hd11f:	data_out=16'h44b;
17'hd120:	data_out=16'ha00;
17'hd121:	data_out=16'h8180;
17'hd122:	data_out=16'h876;
17'hd123:	data_out=16'h858f;
17'hd124:	data_out=16'h858c;
17'hd125:	data_out=16'h8100;
17'hd126:	data_out=16'h8474;
17'hd127:	data_out=16'ha00;
17'hd128:	data_out=16'h818c;
17'hd129:	data_out=16'h1b5;
17'hd12a:	data_out=16'h89ff;
17'hd12b:	data_out=16'ha00;
17'hd12c:	data_out=16'h1f2;
17'hd12d:	data_out=16'h813b;
17'hd12e:	data_out=16'h8981;
17'hd12f:	data_out=16'ha00;
17'hd130:	data_out=16'h8813;
17'hd131:	data_out=16'ha00;
17'hd132:	data_out=16'h8664;
17'hd133:	data_out=16'h772;
17'hd134:	data_out=16'ha00;
17'hd135:	data_out=16'h8231;
17'hd136:	data_out=16'h8465;
17'hd137:	data_out=16'h898c;
17'hd138:	data_out=16'ha00;
17'hd139:	data_out=16'h7a9;
17'hd13a:	data_out=16'h2ab;
17'hd13b:	data_out=16'h38b;
17'hd13c:	data_out=16'h89b0;
17'hd13d:	data_out=16'ha00;
17'hd13e:	data_out=16'h818c;
17'hd13f:	data_out=16'h8eb;
17'hd140:	data_out=16'h35f;
17'hd141:	data_out=16'h89ff;
17'hd142:	data_out=16'h8726;
17'hd143:	data_out=16'h80b9;
17'hd144:	data_out=16'ha00;
17'hd145:	data_out=16'h552;
17'hd146:	data_out=16'h83be;
17'hd147:	data_out=16'hf;
17'hd148:	data_out=16'h83b6;
17'hd149:	data_out=16'h8024;
17'hd14a:	data_out=16'h864c;
17'hd14b:	data_out=16'h8a00;
17'hd14c:	data_out=16'h84be;
17'hd14d:	data_out=16'h91d;
17'hd14e:	data_out=16'h89ff;
17'hd14f:	data_out=16'h8323;
17'hd150:	data_out=16'h2ce;
17'hd151:	data_out=16'h8764;
17'hd152:	data_out=16'h845b;
17'hd153:	data_out=16'ha00;
17'hd154:	data_out=16'ha00;
17'hd155:	data_out=16'h8a00;
17'hd156:	data_out=16'h3b1;
17'hd157:	data_out=16'h52a;
17'hd158:	data_out=16'h8a00;
17'hd159:	data_out=16'h490;
17'hd15a:	data_out=16'h85e4;
17'hd15b:	data_out=16'ha00;
17'hd15c:	data_out=16'h9e1;
17'hd15d:	data_out=16'h80ed;
17'hd15e:	data_out=16'h8cf;
17'hd15f:	data_out=16'h11a;
17'hd160:	data_out=16'h85cf;
17'hd161:	data_out=16'ha00;
17'hd162:	data_out=16'h89ff;
17'hd163:	data_out=16'h6c6;
17'hd164:	data_out=16'ha00;
17'hd165:	data_out=16'h6a8;
17'hd166:	data_out=16'h655;
17'hd167:	data_out=16'h8070;
17'hd168:	data_out=16'h8184;
17'hd169:	data_out=16'h89ff;
17'hd16a:	data_out=16'h8168;
17'hd16b:	data_out=16'ha00;
17'hd16c:	data_out=16'h3a2;
17'hd16d:	data_out=16'h71b;
17'hd16e:	data_out=16'h8168;
17'hd16f:	data_out=16'h80ac;
17'hd170:	data_out=16'h816e;
17'hd171:	data_out=16'h89ff;
17'hd172:	data_out=16'ha00;
17'hd173:	data_out=16'ha00;
17'hd174:	data_out=16'h88b8;
17'hd175:	data_out=16'h883c;
17'hd176:	data_out=16'ha00;
17'hd177:	data_out=16'hfb;
17'hd178:	data_out=16'h810f;
17'hd179:	data_out=16'h89ff;
17'hd17a:	data_out=16'h477;
17'hd17b:	data_out=16'h818d;
17'hd17c:	data_out=16'h8030;
17'hd17d:	data_out=16'haf;
17'hd17e:	data_out=16'h816;
17'hd17f:	data_out=16'h5bc;
17'hd180:	data_out=16'h129;
17'hd181:	data_out=16'h4d;
17'hd182:	data_out=16'h806a;
17'hd183:	data_out=16'h40;
17'hd184:	data_out=16'h3a;
17'hd185:	data_out=16'h2a;
17'hd186:	data_out=16'h801d;
17'hd187:	data_out=16'h1d;
17'hd188:	data_out=16'ha;
17'hd189:	data_out=16'ha0;
17'hd18a:	data_out=16'h20;
17'hd18b:	data_out=16'h8052;
17'hd18c:	data_out=16'h8070;
17'hd18d:	data_out=16'h1c;
17'hd18e:	data_out=16'h8014;
17'hd18f:	data_out=16'h800f;
17'hd190:	data_out=16'h3;
17'hd191:	data_out=16'h73;
17'hd192:	data_out=16'h803f;
17'hd193:	data_out=16'h54;
17'hd194:	data_out=16'h8027;
17'hd195:	data_out=16'h8e;
17'hd196:	data_out=16'h6d;
17'hd197:	data_out=16'h804b;
17'hd198:	data_out=16'h8009;
17'hd199:	data_out=16'h5a;
17'hd19a:	data_out=16'h19;
17'hd19b:	data_out=16'h18;
17'hd19c:	data_out=16'h87;
17'hd19d:	data_out=16'h2b;
17'hd19e:	data_out=16'he;
17'hd19f:	data_out=16'h8001;
17'hd1a0:	data_out=16'ha3;
17'hd1a1:	data_out=16'h8009;
17'hd1a2:	data_out=16'h61;
17'hd1a3:	data_out=16'h803e;
17'hd1a4:	data_out=16'h8041;
17'hd1a5:	data_out=16'h10;
17'hd1a6:	data_out=16'h4a;
17'hd1a7:	data_out=16'h35;
17'hd1a8:	data_out=16'h8016;
17'hd1a9:	data_out=16'h31;
17'hd1aa:	data_out=16'h8043;
17'hd1ab:	data_out=16'hf4;
17'hd1ac:	data_out=16'h24;
17'hd1ad:	data_out=16'h800e;
17'hd1ae:	data_out=16'h805e;
17'hd1af:	data_out=16'h5d;
17'hd1b0:	data_out=16'h8034;
17'hd1b1:	data_out=16'ha8;
17'hd1b2:	data_out=16'h8021;
17'hd1b3:	data_out=16'h2;
17'hd1b4:	data_out=16'hb7;
17'hd1b5:	data_out=16'h8046;
17'hd1b6:	data_out=16'h8051;
17'hd1b7:	data_out=16'h8067;
17'hd1b8:	data_out=16'hcf;
17'hd1b9:	data_out=16'h2e;
17'hd1ba:	data_out=16'h8002;
17'hd1bb:	data_out=16'h4f;
17'hd1bc:	data_out=16'h8080;
17'hd1bd:	data_out=16'h12f;
17'hd1be:	data_out=16'h800b;
17'hd1bf:	data_out=16'h37;
17'hd1c0:	data_out=16'h1a;
17'hd1c1:	data_out=16'h8067;
17'hd1c2:	data_out=16'h800f;
17'hd1c3:	data_out=16'h8032;
17'hd1c4:	data_out=16'h5c;
17'hd1c5:	data_out=16'ha6;
17'hd1c6:	data_out=16'h8036;
17'hd1c7:	data_out=16'h3;
17'hd1c8:	data_out=16'h8039;
17'hd1c9:	data_out=16'h1b;
17'hd1ca:	data_out=16'h801d;
17'hd1cb:	data_out=16'h8098;
17'hd1cc:	data_out=16'h8011;
17'hd1cd:	data_out=16'h84;
17'hd1ce:	data_out=16'h8034;
17'hd1cf:	data_out=16'h8008;
17'hd1d0:	data_out=16'hc;
17'hd1d1:	data_out=16'h27;
17'hd1d2:	data_out=16'h8028;
17'hd1d3:	data_out=16'h16;
17'hd1d4:	data_out=16'h5e;
17'hd1d5:	data_out=16'h80a0;
17'hd1d6:	data_out=16'h4;
17'hd1d7:	data_out=16'h15;
17'hd1d8:	data_out=16'h809a;
17'hd1d9:	data_out=16'h18;
17'hd1da:	data_out=16'h8080;
17'hd1db:	data_out=16'h18;
17'hd1dc:	data_out=16'h10;
17'hd1dd:	data_out=16'h8;
17'hd1de:	data_out=16'h36;
17'hd1df:	data_out=16'h10;
17'hd1e0:	data_out=16'h2e;
17'hd1e1:	data_out=16'h7a;
17'hd1e2:	data_out=16'h807c;
17'hd1e3:	data_out=16'h800b;
17'hd1e4:	data_out=16'hd9;
17'hd1e5:	data_out=16'h41;
17'hd1e6:	data_out=16'h3f;
17'hd1e7:	data_out=16'h8027;
17'hd1e8:	data_out=16'h8010;
17'hd1e9:	data_out=16'h806f;
17'hd1ea:	data_out=16'h800d;
17'hd1eb:	data_out=16'h9b;
17'hd1ec:	data_out=16'h4;
17'hd1ed:	data_out=16'h4;
17'hd1ee:	data_out=16'h800a;
17'hd1ef:	data_out=16'h1a;
17'hd1f0:	data_out=16'h800e;
17'hd1f1:	data_out=16'h806f;
17'hd1f2:	data_out=16'h5e;
17'hd1f3:	data_out=16'h96;
17'hd1f4:	data_out=16'h802e;
17'hd1f5:	data_out=16'h8063;
17'hd1f6:	data_out=16'h83;
17'hd1f7:	data_out=16'h25;
17'hd1f8:	data_out=16'h37;
17'hd1f9:	data_out=16'h8085;
17'hd1fa:	data_out=16'h8023;
17'hd1fb:	data_out=16'h800f;
17'hd1fc:	data_out=16'h8021;
17'hd1fd:	data_out=16'h8026;
17'hd1fe:	data_out=16'ha1;
17'hd1ff:	data_out=16'h2c;
17'hd200:	data_out=16'h8010;
17'hd201:	data_out=16'h10;
17'hd202:	data_out=16'h3;
17'hd203:	data_out=16'h2;
17'hd204:	data_out=16'h4;
17'hd205:	data_out=16'h8004;
17'hd206:	data_out=16'h1;
17'hd207:	data_out=16'h8007;
17'hd208:	data_out=16'h800b;
17'hd209:	data_out=16'h8004;
17'hd20a:	data_out=16'h800c;
17'hd20b:	data_out=16'h800e;
17'hd20c:	data_out=16'h800a;
17'hd20d:	data_out=16'h8005;
17'hd20e:	data_out=16'h8008;
17'hd20f:	data_out=16'h800c;
17'hd210:	data_out=16'h800e;
17'hd211:	data_out=16'h0;
17'hd212:	data_out=16'h8009;
17'hd213:	data_out=16'h800a;
17'hd214:	data_out=16'h800f;
17'hd215:	data_out=16'h8005;
17'hd216:	data_out=16'h8007;
17'hd217:	data_out=16'h800a;
17'hd218:	data_out=16'h8008;
17'hd219:	data_out=16'h8024;
17'hd21a:	data_out=16'h4;
17'hd21b:	data_out=16'h8007;
17'hd21c:	data_out=16'h8010;
17'hd21d:	data_out=16'h6;
17'hd21e:	data_out=16'h800b;
17'hd21f:	data_out=16'ha;
17'hd220:	data_out=16'h800a;
17'hd221:	data_out=16'h8007;
17'hd222:	data_out=16'h8006;
17'hd223:	data_out=16'h1a;
17'hd224:	data_out=16'h25;
17'hd225:	data_out=16'h800b;
17'hd226:	data_out=16'h800d;
17'hd227:	data_out=16'h8002;
17'hd228:	data_out=16'h6;
17'hd229:	data_out=16'h800c;
17'hd22a:	data_out=16'h8008;
17'hd22b:	data_out=16'h8008;
17'hd22c:	data_out=16'h8007;
17'hd22d:	data_out=16'h8006;
17'hd22e:	data_out=16'h800c;
17'hd22f:	data_out=16'h14;
17'hd230:	data_out=16'h8011;
17'hd231:	data_out=16'h8011;
17'hd232:	data_out=16'h8018;
17'hd233:	data_out=16'h8012;
17'hd234:	data_out=16'h800e;
17'hd235:	data_out=16'h1;
17'hd236:	data_out=16'he;
17'hd237:	data_out=16'h800c;
17'hd238:	data_out=16'h26;
17'hd239:	data_out=16'h800f;
17'hd23a:	data_out=16'h16;
17'hd23b:	data_out=16'h2;
17'hd23c:	data_out=16'h800c;
17'hd23d:	data_out=16'h8004;
17'hd23e:	data_out=16'h2;
17'hd23f:	data_out=16'h8000;
17'hd240:	data_out=16'h27;
17'hd241:	data_out=16'h8004;
17'hd242:	data_out=16'h5;
17'hd243:	data_out=16'ha;
17'hd244:	data_out=16'h8002;
17'hd245:	data_out=16'hb;
17'hd246:	data_out=16'h8016;
17'hd247:	data_out=16'h20;
17'hd248:	data_out=16'h801a;
17'hd249:	data_out=16'h6;
17'hd24a:	data_out=16'h8003;
17'hd24b:	data_out=16'h10;
17'hd24c:	data_out=16'h7;
17'hd24d:	data_out=16'h800b;
17'hd24e:	data_out=16'h8005;
17'hd24f:	data_out=16'h6;
17'hd250:	data_out=16'h21;
17'hd251:	data_out=16'h800c;
17'hd252:	data_out=16'h16;
17'hd253:	data_out=16'h8008;
17'hd254:	data_out=16'h3;
17'hd255:	data_out=16'h4;
17'hd256:	data_out=16'h800c;
17'hd257:	data_out=16'h8003;
17'hd258:	data_out=16'h800a;
17'hd259:	data_out=16'h7;
17'hd25a:	data_out=16'h800f;
17'hd25b:	data_out=16'h13;
17'hd25c:	data_out=16'h8003;
17'hd25d:	data_out=16'h8006;
17'hd25e:	data_out=16'h8004;
17'hd25f:	data_out=16'h800a;
17'hd260:	data_out=16'h800c;
17'hd261:	data_out=16'h8004;
17'hd262:	data_out=16'h8003;
17'hd263:	data_out=16'h8012;
17'hd264:	data_out=16'h8011;
17'hd265:	data_out=16'h4;
17'hd266:	data_out=16'h8021;
17'hd267:	data_out=16'h800b;
17'hd268:	data_out=16'h2;
17'hd269:	data_out=16'h2;
17'hd26a:	data_out=16'h3;
17'hd26b:	data_out=16'h8005;
17'hd26c:	data_out=16'h9;
17'hd26d:	data_out=16'h800f;
17'hd26e:	data_out=16'h8001;
17'hd26f:	data_out=16'h800b;
17'hd270:	data_out=16'h6;
17'hd271:	data_out=16'h8005;
17'hd272:	data_out=16'h8013;
17'hd273:	data_out=16'h8008;
17'hd274:	data_out=16'h8016;
17'hd275:	data_out=16'h800a;
17'hd276:	data_out=16'h8016;
17'hd277:	data_out=16'h12;
17'hd278:	data_out=16'h8005;
17'hd279:	data_out=16'h800b;
17'hd27a:	data_out=16'h800f;
17'hd27b:	data_out=16'h5;
17'hd27c:	data_out=16'h8004;
17'hd27d:	data_out=16'hd;
17'hd27e:	data_out=16'h8003;
17'hd27f:	data_out=16'h8002;
17'hd280:	data_out=16'h82e5;
17'hd281:	data_out=16'h8027;
17'hd282:	data_out=16'h80b1;
17'hd283:	data_out=16'h816c;
17'hd284:	data_out=16'h80fe;
17'hd285:	data_out=16'h87;
17'hd286:	data_out=16'h8080;
17'hd287:	data_out=16'h81c9;
17'hd288:	data_out=16'h8070;
17'hd289:	data_out=16'h832d;
17'hd28a:	data_out=16'h80d6;
17'hd28b:	data_out=16'heb;
17'hd28c:	data_out=16'hd1;
17'hd28d:	data_out=16'h80db;
17'hd28e:	data_out=16'h8039;
17'hd28f:	data_out=16'h80e8;
17'hd290:	data_out=16'h8292;
17'hd291:	data_out=16'h8053;
17'hd292:	data_out=16'h812e;
17'hd293:	data_out=16'h8227;
17'hd294:	data_out=16'h8028;
17'hd295:	data_out=16'h8131;
17'hd296:	data_out=16'h81bc;
17'hd297:	data_out=16'h1e;
17'hd298:	data_out=16'h80b0;
17'hd299:	data_out=16'h41;
17'hd29a:	data_out=16'h80b6;
17'hd29b:	data_out=16'h170;
17'hd29c:	data_out=16'h48;
17'hd29d:	data_out=16'h8011;
17'hd29e:	data_out=16'h805a;
17'hd29f:	data_out=16'h80e3;
17'hd2a0:	data_out=16'h800c;
17'hd2a1:	data_out=16'h8038;
17'hd2a2:	data_out=16'h82cb;
17'hd2a3:	data_out=16'h807b;
17'hd2a4:	data_out=16'h8080;
17'hd2a5:	data_out=16'h8274;
17'hd2a6:	data_out=16'h827b;
17'hd2a7:	data_out=16'h77;
17'hd2a8:	data_out=16'h8025;
17'hd2a9:	data_out=16'h8133;
17'hd2aa:	data_out=16'h8291;
17'hd2ab:	data_out=16'h69;
17'hd2ac:	data_out=16'h813b;
17'hd2ad:	data_out=16'h8324;
17'hd2ae:	data_out=16'h81a9;
17'hd2af:	data_out=16'h808f;
17'hd2b0:	data_out=16'h808b;
17'hd2b1:	data_out=16'h1e;
17'hd2b2:	data_out=16'h80a9;
17'hd2b3:	data_out=16'h8049;
17'hd2b4:	data_out=16'h80a7;
17'hd2b5:	data_out=16'hfa;
17'hd2b6:	data_out=16'h8079;
17'hd2b7:	data_out=16'h809a;
17'hd2b8:	data_out=16'h6;
17'hd2b9:	data_out=16'h8029;
17'hd2ba:	data_out=16'h837e;
17'hd2bb:	data_out=16'hf;
17'hd2bc:	data_out=16'h4e;
17'hd2bd:	data_out=16'h82e4;
17'hd2be:	data_out=16'h802d;
17'hd2bf:	data_out=16'h26;
17'hd2c0:	data_out=16'h8322;
17'hd2c1:	data_out=16'hff;
17'hd2c2:	data_out=16'h8287;
17'hd2c3:	data_out=16'h22;
17'hd2c4:	data_out=16'h8086;
17'hd2c5:	data_out=16'h8156;
17'hd2c6:	data_out=16'h48;
17'hd2c7:	data_out=16'h8377;
17'hd2c8:	data_out=16'h810d;
17'hd2c9:	data_out=16'h8289;
17'hd2ca:	data_out=16'h814e;
17'hd2cb:	data_out=16'h80c0;
17'hd2cc:	data_out=16'h82e1;
17'hd2cd:	data_out=16'h82bf;
17'hd2ce:	data_out=16'h81a9;
17'hd2cf:	data_out=16'h8315;
17'hd2d0:	data_out=16'h82d6;
17'hd2d1:	data_out=16'h3f;
17'hd2d2:	data_out=16'h80f3;
17'hd2d3:	data_out=16'h1f6;
17'hd2d4:	data_out=16'h80d8;
17'hd2d5:	data_out=16'h8e;
17'hd2d6:	data_out=16'h832b;
17'hd2d7:	data_out=16'h8379;
17'hd2d8:	data_out=16'h31;
17'hd2d9:	data_out=16'h83b3;
17'hd2da:	data_out=16'h239;
17'hd2db:	data_out=16'hc7;
17'hd2dc:	data_out=16'h16b;
17'hd2dd:	data_out=16'h81f4;
17'hd2de:	data_out=16'h80ce;
17'hd2df:	data_out=16'h80b7;
17'hd2e0:	data_out=16'h82d2;
17'hd2e1:	data_out=16'h8052;
17'hd2e2:	data_out=16'h13f;
17'hd2e3:	data_out=16'h8026;
17'hd2e4:	data_out=16'h812e;
17'hd2e5:	data_out=16'h80e0;
17'hd2e6:	data_out=16'h38;
17'hd2e7:	data_out=16'h816f;
17'hd2e8:	data_out=16'h802a;
17'hd2e9:	data_out=16'h80ad;
17'hd2ea:	data_out=16'h8042;
17'hd2eb:	data_out=16'h80da;
17'hd2ec:	data_out=16'h83a2;
17'hd2ed:	data_out=16'h802d;
17'hd2ee:	data_out=16'h8045;
17'hd2ef:	data_out=16'h8097;
17'hd2f0:	data_out=16'h8040;
17'hd2f1:	data_out=16'h80d9;
17'hd2f2:	data_out=16'h81a8;
17'hd2f3:	data_out=16'h80d0;
17'hd2f4:	data_out=16'h8085;
17'hd2f5:	data_out=16'h1d4;
17'hd2f6:	data_out=16'h18;
17'hd2f7:	data_out=16'h83a5;
17'hd2f8:	data_out=16'h28;
17'hd2f9:	data_out=16'h81c1;
17'hd2fa:	data_out=16'h801d;
17'hd2fb:	data_out=16'h802a;
17'hd2fc:	data_out=16'hf;
17'hd2fd:	data_out=16'hbb;
17'hd2fe:	data_out=16'h82fc;
17'hd2ff:	data_out=16'h8316;
17'hd300:	data_out=16'h80db;
17'hd301:	data_out=16'h272;
17'hd302:	data_out=16'h8129;
17'hd303:	data_out=16'h801a;
17'hd304:	data_out=16'h8352;
17'hd305:	data_out=16'hb4;
17'hd306:	data_out=16'h81b9;
17'hd307:	data_out=16'h812d;
17'hd308:	data_out=16'h8182;
17'hd309:	data_out=16'h833b;
17'hd30a:	data_out=16'h80b4;
17'hd30b:	data_out=16'h6a;
17'hd30c:	data_out=16'h830a;
17'hd30d:	data_out=16'h7e;
17'hd30e:	data_out=16'h80d7;
17'hd30f:	data_out=16'h8057;
17'hd310:	data_out=16'h82ab;
17'hd311:	data_out=16'h829e;
17'hd312:	data_out=16'h2bd;
17'hd313:	data_out=16'h8119;
17'hd314:	data_out=16'h267;
17'hd315:	data_out=16'h8152;
17'hd316:	data_out=16'h80ea;
17'hd317:	data_out=16'h335;
17'hd318:	data_out=16'h80fb;
17'hd319:	data_out=16'h816d;
17'hd31a:	data_out=16'h82a6;
17'hd31b:	data_out=16'h3d8;
17'hd31c:	data_out=16'h48;
17'hd31d:	data_out=16'h1d4;
17'hd31e:	data_out=16'h2fc;
17'hd31f:	data_out=16'h81fb;
17'hd320:	data_out=16'h504;
17'hd321:	data_out=16'h80d2;
17'hd322:	data_out=16'h17;
17'hd323:	data_out=16'h82eb;
17'hd324:	data_out=16'h82eb;
17'hd325:	data_out=16'h820f;
17'hd326:	data_out=16'h83f1;
17'hd327:	data_out=16'h27c;
17'hd328:	data_out=16'h80d0;
17'hd329:	data_out=16'h29;
17'hd32a:	data_out=16'h810a;
17'hd32b:	data_out=16'h8082;
17'hd32c:	data_out=16'h80f3;
17'hd32d:	data_out=16'h81c9;
17'hd32e:	data_out=16'h65;
17'hd32f:	data_out=16'h452;
17'hd330:	data_out=16'h82db;
17'hd331:	data_out=16'h179;
17'hd332:	data_out=16'h82d0;
17'hd333:	data_out=16'h263;
17'hd334:	data_out=16'h80db;
17'hd335:	data_out=16'h8291;
17'hd336:	data_out=16'hd2;
17'hd337:	data_out=16'h8055;
17'hd338:	data_out=16'h8099;
17'hd339:	data_out=16'h1b6;
17'hd33a:	data_out=16'h805f;
17'hd33b:	data_out=16'h81e8;
17'hd33c:	data_out=16'h77;
17'hd33d:	data_out=16'h81d8;
17'hd33e:	data_out=16'h80c3;
17'hd33f:	data_out=16'h807e;
17'hd340:	data_out=16'h8301;
17'hd341:	data_out=16'hf8;
17'hd342:	data_out=16'h81b1;
17'hd343:	data_out=16'h8269;
17'hd344:	data_out=16'h817e;
17'hd345:	data_out=16'h81db;
17'hd346:	data_out=16'h4c;
17'hd347:	data_out=16'h81cf;
17'hd348:	data_out=16'h17c;
17'hd349:	data_out=16'h8249;
17'hd34a:	data_out=16'h8123;
17'hd34b:	data_out=16'h8047;
17'hd34c:	data_out=16'h8120;
17'hd34d:	data_out=16'h47;
17'hd34e:	data_out=16'h92;
17'hd34f:	data_out=16'h81fe;
17'hd350:	data_out=16'h8327;
17'hd351:	data_out=16'h8236;
17'hd352:	data_out=16'h83bc;
17'hd353:	data_out=16'h534;
17'hd354:	data_out=16'h3b3;
17'hd355:	data_out=16'h81be;
17'hd356:	data_out=16'h82a7;
17'hd357:	data_out=16'h8459;
17'hd358:	data_out=16'h81d0;
17'hd359:	data_out=16'h8450;
17'hd35a:	data_out=16'h343;
17'hd35b:	data_out=16'h8093;
17'hd35c:	data_out=16'h330;
17'hd35d:	data_out=16'he5;
17'hd35e:	data_out=16'h3ae;
17'hd35f:	data_out=16'h147;
17'hd360:	data_out=16'h842f;
17'hd361:	data_out=16'h81c9;
17'hd362:	data_out=16'h24f;
17'hd363:	data_out=16'h28f;
17'hd364:	data_out=16'h81ef;
17'hd365:	data_out=16'h8068;
17'hd366:	data_out=16'h815e;
17'hd367:	data_out=16'h8081;
17'hd368:	data_out=16'h80d9;
17'hd369:	data_out=16'h814b;
17'hd36a:	data_out=16'h80dc;
17'hd36b:	data_out=16'h8166;
17'hd36c:	data_out=16'h20d;
17'hd36d:	data_out=16'h28a;
17'hd36e:	data_out=16'h80e3;
17'hd36f:	data_out=16'h90;
17'hd370:	data_out=16'h80e4;
17'hd371:	data_out=16'h16;
17'hd372:	data_out=16'h825a;
17'hd373:	data_out=16'h80b0;
17'hd374:	data_out=16'h82e3;
17'hd375:	data_out=16'h808c;
17'hd376:	data_out=16'h80c2;
17'hd377:	data_out=16'h86cb;
17'hd378:	data_out=16'h81cb;
17'hd379:	data_out=16'h49;
17'hd37a:	data_out=16'h293;
17'hd37b:	data_out=16'h80c5;
17'hd37c:	data_out=16'h7f;
17'hd37d:	data_out=16'h806c;
17'hd37e:	data_out=16'h83a4;
17'hd37f:	data_out=16'h83ee;
17'hd380:	data_out=16'h829a;
17'hd381:	data_out=16'h10b;
17'hd382:	data_out=16'h2ae;
17'hd383:	data_out=16'h80ae;
17'hd384:	data_out=16'h8999;
17'hd385:	data_out=16'h84b0;
17'hd386:	data_out=16'h80e3;
17'hd387:	data_out=16'h89ff;
17'hd388:	data_out=16'h8669;
17'hd389:	data_out=16'h8107;
17'hd38a:	data_out=16'h8a00;
17'hd38b:	data_out=16'h3cf;
17'hd38c:	data_out=16'h89fd;
17'hd38d:	data_out=16'h3c5;
17'hd38e:	data_out=16'h8094;
17'hd38f:	data_out=16'h38c;
17'hd390:	data_out=16'h45b;
17'hd391:	data_out=16'h8940;
17'hd392:	data_out=16'h839;
17'hd393:	data_out=16'h81aa;
17'hd394:	data_out=16'h9fe;
17'hd395:	data_out=16'h84f5;
17'hd396:	data_out=16'h8a00;
17'hd397:	data_out=16'h9fb;
17'hd398:	data_out=16'h307;
17'hd399:	data_out=16'h85ab;
17'hd39a:	data_out=16'h898c;
17'hd39b:	data_out=16'ha00;
17'hd39c:	data_out=16'h826b;
17'hd39d:	data_out=16'h159;
17'hd39e:	data_out=16'h9fb;
17'hd39f:	data_out=16'h83d6;
17'hd3a0:	data_out=16'h9ff;
17'hd3a1:	data_out=16'h8097;
17'hd3a2:	data_out=16'h7ff;
17'hd3a3:	data_out=16'h8a00;
17'hd3a4:	data_out=16'h8a00;
17'hd3a5:	data_out=16'h833f;
17'hd3a6:	data_out=16'h8a00;
17'hd3a7:	data_out=16'h8f9;
17'hd3a8:	data_out=16'h80a1;
17'hd3a9:	data_out=16'h77e;
17'hd3aa:	data_out=16'h8230;
17'hd3ab:	data_out=16'h50d;
17'hd3ac:	data_out=16'h8a00;
17'hd3ad:	data_out=16'h8766;
17'hd3ae:	data_out=16'h9ca;
17'hd3af:	data_out=16'h9ff;
17'hd3b0:	data_out=16'h8a00;
17'hd3b1:	data_out=16'h89fd;
17'hd3b2:	data_out=16'h8a00;
17'hd3b3:	data_out=16'ha00;
17'hd3b4:	data_out=16'h86e2;
17'hd3b5:	data_out=16'h89fe;
17'hd3b6:	data_out=16'h54a;
17'hd3b7:	data_out=16'h319;
17'hd3b8:	data_out=16'h138;
17'hd3b9:	data_out=16'ha00;
17'hd3ba:	data_out=16'h544;
17'hd3bb:	data_out=16'h89ff;
17'hd3bc:	data_out=16'h48d;
17'hd3bd:	data_out=16'h258;
17'hd3be:	data_out=16'h80a3;
17'hd3bf:	data_out=16'h84b0;
17'hd3c0:	data_out=16'h89ec;
17'hd3c1:	data_out=16'h445;
17'hd3c2:	data_out=16'h8a00;
17'hd3c3:	data_out=16'h82c7;
17'hd3c4:	data_out=16'h88ac;
17'hd3c5:	data_out=16'h8551;
17'hd3c6:	data_out=16'h2e;
17'hd3c7:	data_out=16'h87ab;
17'hd3c8:	data_out=16'h9ff;
17'hd3c9:	data_out=16'h83db;
17'hd3ca:	data_out=16'h8847;
17'hd3cb:	data_out=16'h8a00;
17'hd3cc:	data_out=16'h880e;
17'hd3cd:	data_out=16'h9fd;
17'hd3ce:	data_out=16'h905;
17'hd3cf:	data_out=16'h885c;
17'hd3d0:	data_out=16'h873e;
17'hd3d1:	data_out=16'h8804;
17'hd3d2:	data_out=16'h8a00;
17'hd3d3:	data_out=16'ha00;
17'hd3d4:	data_out=16'h9ff;
17'hd3d5:	data_out=16'h8145;
17'hd3d6:	data_out=16'h844b;
17'hd3d7:	data_out=16'h8405;
17'hd3d8:	data_out=16'h1ac;
17'hd3d9:	data_out=16'h89e9;
17'hd3da:	data_out=16'ha00;
17'hd3db:	data_out=16'h86cd;
17'hd3dc:	data_out=16'h9fd;
17'hd3dd:	data_out=16'h49f;
17'hd3de:	data_out=16'h9fe;
17'hd3df:	data_out=16'h7cd;
17'hd3e0:	data_out=16'h8a00;
17'hd3e1:	data_out=16'h89fb;
17'hd3e2:	data_out=16'h72a;
17'hd3e3:	data_out=16'ha00;
17'hd3e4:	data_out=16'h8341;
17'hd3e5:	data_out=16'h8681;
17'hd3e6:	data_out=16'h84e0;
17'hd3e7:	data_out=16'h14b;
17'hd3e8:	data_out=16'h809a;
17'hd3e9:	data_out=16'h88e6;
17'hd3ea:	data_out=16'h808f;
17'hd3eb:	data_out=16'h878a;
17'hd3ec:	data_out=16'h87f2;
17'hd3ed:	data_out=16'ha00;
17'hd3ee:	data_out=16'h8090;
17'hd3ef:	data_out=16'h89ff;
17'hd3f0:	data_out=16'h8093;
17'hd3f1:	data_out=16'h24f;
17'hd3f2:	data_out=16'h89fd;
17'hd3f3:	data_out=16'h89fe;
17'hd3f4:	data_out=16'h8a00;
17'hd3f5:	data_out=16'h89c7;
17'hd3f6:	data_out=16'h82e3;
17'hd3f7:	data_out=16'h890b;
17'hd3f8:	data_out=16'h86f0;
17'hd3f9:	data_out=16'h9fa;
17'hd3fa:	data_out=16'ha00;
17'hd3fb:	data_out=16'h80a4;
17'hd3fc:	data_out=16'h49a;
17'hd3fd:	data_out=16'h53;
17'hd3fe:	data_out=16'h8057;
17'hd3ff:	data_out=16'h8819;
17'hd400:	data_out=16'h89c7;
17'hd401:	data_out=16'h89f9;
17'hd402:	data_out=16'h505;
17'hd403:	data_out=16'h8074;
17'hd404:	data_out=16'h89ff;
17'hd405:	data_out=16'h8a00;
17'hd406:	data_out=16'h595;
17'hd407:	data_out=16'h2d;
17'hd408:	data_out=16'h509;
17'hd409:	data_out=16'h9fe;
17'hd40a:	data_out=16'h8a00;
17'hd40b:	data_out=16'ha00;
17'hd40c:	data_out=16'h80f8;
17'hd40d:	data_out=16'h7a8;
17'hd40e:	data_out=16'h81cb;
17'hd40f:	data_out=16'h755;
17'hd410:	data_out=16'h9ec;
17'hd411:	data_out=16'h89c5;
17'hd412:	data_out=16'h9f8;
17'hd413:	data_out=16'h69b;
17'hd414:	data_out=16'h9f9;
17'hd415:	data_out=16'h8a00;
17'hd416:	data_out=16'h8a00;
17'hd417:	data_out=16'h9f9;
17'hd418:	data_out=16'h70c;
17'hd419:	data_out=16'h83b0;
17'hd41a:	data_out=16'h8a00;
17'hd41b:	data_out=16'h9ff;
17'hd41c:	data_out=16'h856d;
17'hd41d:	data_out=16'h89ea;
17'hd41e:	data_out=16'h9f4;
17'hd41f:	data_out=16'h9dc;
17'hd420:	data_out=16'h27f;
17'hd421:	data_out=16'h81b2;
17'hd422:	data_out=16'h445;
17'hd423:	data_out=16'h83b0;
17'hd424:	data_out=16'h83ac;
17'hd425:	data_out=16'h5ad;
17'hd426:	data_out=16'h9f9;
17'hd427:	data_out=16'h25f;
17'hd428:	data_out=16'h8161;
17'hd429:	data_out=16'h821d;
17'hd42a:	data_out=16'h784;
17'hd42b:	data_out=16'ha00;
17'hd42c:	data_out=16'h8a00;
17'hd42d:	data_out=16'h8260;
17'hd42e:	data_out=16'h953;
17'hd42f:	data_out=16'h8337;
17'hd430:	data_out=16'h8a00;
17'hd431:	data_out=16'h89f2;
17'hd432:	data_out=16'h8a00;
17'hd433:	data_out=16'h9ff;
17'hd434:	data_out=16'h89ed;
17'hd435:	data_out=16'h89f2;
17'hd436:	data_out=16'h9ff;
17'hd437:	data_out=16'h912;
17'hd438:	data_out=16'h89d3;
17'hd439:	data_out=16'ha00;
17'hd43a:	data_out=16'h9ee;
17'hd43b:	data_out=16'h89f0;
17'hd43c:	data_out=16'h636;
17'hd43d:	data_out=16'h89f7;
17'hd43e:	data_out=16'h8160;
17'hd43f:	data_out=16'h8a00;
17'hd440:	data_out=16'h8a00;
17'hd441:	data_out=16'h9f6;
17'hd442:	data_out=16'h89f3;
17'hd443:	data_out=16'h45f;
17'hd444:	data_out=16'h897f;
17'hd445:	data_out=16'h8a00;
17'hd446:	data_out=16'h8675;
17'hd447:	data_out=16'h9f0;
17'hd448:	data_out=16'ha00;
17'hd449:	data_out=16'h4ad;
17'hd44a:	data_out=16'h89e2;
17'hd44b:	data_out=16'h88e8;
17'hd44c:	data_out=16'h8a00;
17'hd44d:	data_out=16'h610;
17'hd44e:	data_out=16'ha00;
17'hd44f:	data_out=16'h81eb;
17'hd450:	data_out=16'h8a00;
17'hd451:	data_out=16'h9dc;
17'hd452:	data_out=16'h856a;
17'hd453:	data_out=16'h9ff;
17'hd454:	data_out=16'h82c5;
17'hd455:	data_out=16'h9e1;
17'hd456:	data_out=16'h483;
17'hd457:	data_out=16'h302;
17'hd458:	data_out=16'h9eb;
17'hd459:	data_out=16'h8a00;
17'hd45a:	data_out=16'h9ff;
17'hd45b:	data_out=16'h8911;
17'hd45c:	data_out=16'h6f8;
17'hd45d:	data_out=16'h89fc;
17'hd45e:	data_out=16'h84ec;
17'hd45f:	data_out=16'h806a;
17'hd460:	data_out=16'h9fd;
17'hd461:	data_out=16'h8a00;
17'hd462:	data_out=16'h9ff;
17'hd463:	data_out=16'h9ff;
17'hd464:	data_out=16'ha00;
17'hd465:	data_out=16'h8a00;
17'hd466:	data_out=16'h3e3;
17'hd467:	data_out=16'h83e8;
17'hd468:	data_out=16'h8186;
17'hd469:	data_out=16'h656;
17'hd46a:	data_out=16'h81d5;
17'hd46b:	data_out=16'h8a00;
17'hd46c:	data_out=16'h89f1;
17'hd46d:	data_out=16'h9ff;
17'hd46e:	data_out=16'h81d6;
17'hd46f:	data_out=16'h8a00;
17'hd470:	data_out=16'h81d2;
17'hd471:	data_out=16'h895;
17'hd472:	data_out=16'h8a00;
17'hd473:	data_out=16'h8a00;
17'hd474:	data_out=16'h8a00;
17'hd475:	data_out=16'h8a00;
17'hd476:	data_out=16'ha00;
17'hd477:	data_out=16'h80bd;
17'hd478:	data_out=16'h8a00;
17'hd479:	data_out=16'h9f3;
17'hd47a:	data_out=16'h9fb;
17'hd47b:	data_out=16'h8160;
17'hd47c:	data_out=16'h38b;
17'hd47d:	data_out=16'h80a8;
17'hd47e:	data_out=16'h9f0;
17'hd47f:	data_out=16'h8a00;
17'hd480:	data_out=16'h89fe;
17'hd481:	data_out=16'h8a00;
17'hd482:	data_out=16'h8a00;
17'hd483:	data_out=16'h863c;
17'hd484:	data_out=16'h89bd;
17'hd485:	data_out=16'h8a00;
17'hd486:	data_out=16'h9f1;
17'hd487:	data_out=16'ha00;
17'hd488:	data_out=16'h84c7;
17'hd489:	data_out=16'ha00;
17'hd48a:	data_out=16'h8a00;
17'hd48b:	data_out=16'ha00;
17'hd48c:	data_out=16'ha00;
17'hd48d:	data_out=16'h8795;
17'hd48e:	data_out=16'h8a00;
17'hd48f:	data_out=16'h8a00;
17'hd490:	data_out=16'h9b7;
17'hd491:	data_out=16'h8a00;
17'hd492:	data_out=16'h7b3;
17'hd493:	data_out=16'h9ff;
17'hd494:	data_out=16'h80f5;
17'hd495:	data_out=16'h8a00;
17'hd496:	data_out=16'h8a00;
17'hd497:	data_out=16'h9d8;
17'hd498:	data_out=16'h8a00;
17'hd499:	data_out=16'ha00;
17'hd49a:	data_out=16'h8a00;
17'hd49b:	data_out=16'h826d;
17'hd49c:	data_out=16'h8a00;
17'hd49d:	data_out=16'h89f7;
17'hd49e:	data_out=16'h8a00;
17'hd49f:	data_out=16'h75f;
17'hd4a0:	data_out=16'h8a00;
17'hd4a1:	data_out=16'h8a00;
17'hd4a2:	data_out=16'h1f3;
17'hd4a3:	data_out=16'ha00;
17'hd4a4:	data_out=16'ha00;
17'hd4a5:	data_out=16'h8c4;
17'hd4a6:	data_out=16'h9fb;
17'hd4a7:	data_out=16'h89be;
17'hd4a8:	data_out=16'h8a00;
17'hd4a9:	data_out=16'h8a00;
17'hd4aa:	data_out=16'h83aa;
17'hd4ab:	data_out=16'ha00;
17'hd4ac:	data_out=16'h8a00;
17'hd4ad:	data_out=16'ha00;
17'hd4ae:	data_out=16'h813c;
17'hd4af:	data_out=16'h8a00;
17'hd4b0:	data_out=16'h89cb;
17'hd4b1:	data_out=16'h8a00;
17'hd4b2:	data_out=16'h89ed;
17'hd4b3:	data_out=16'h87a0;
17'hd4b4:	data_out=16'h89fb;
17'hd4b5:	data_out=16'h89ff;
17'hd4b6:	data_out=16'h8a00;
17'hd4b7:	data_out=16'h8a00;
17'hd4b8:	data_out=16'h8a00;
17'hd4b9:	data_out=16'h8a00;
17'hd4ba:	data_out=16'ha00;
17'hd4bb:	data_out=16'h84bf;
17'hd4bc:	data_out=16'h8a00;
17'hd4bd:	data_out=16'h8a00;
17'hd4be:	data_out=16'h8a00;
17'hd4bf:	data_out=16'h8a00;
17'hd4c0:	data_out=16'h89fe;
17'hd4c1:	data_out=16'h88f7;
17'hd4c2:	data_out=16'ha00;
17'hd4c3:	data_out=16'h7af;
17'hd4c4:	data_out=16'h89fe;
17'hd4c5:	data_out=16'h8a00;
17'hd4c6:	data_out=16'h8a00;
17'hd4c7:	data_out=16'ha00;
17'hd4c8:	data_out=16'h9ec;
17'hd4c9:	data_out=16'h98e;
17'hd4ca:	data_out=16'ha00;
17'hd4cb:	data_out=16'ha00;
17'hd4cc:	data_out=16'h619;
17'hd4cd:	data_out=16'h1c6;
17'hd4ce:	data_out=16'h8720;
17'hd4cf:	data_out=16'h9fe;
17'hd4d0:	data_out=16'h89fd;
17'hd4d1:	data_out=16'h81f6;
17'hd4d2:	data_out=16'ha00;
17'hd4d3:	data_out=16'h89fd;
17'hd4d4:	data_out=16'h8a00;
17'hd4d5:	data_out=16'h9a6;
17'hd4d6:	data_out=16'h89ff;
17'hd4d7:	data_out=16'h8a00;
17'hd4d8:	data_out=16'h8a00;
17'hd4d9:	data_out=16'h8a00;
17'hd4da:	data_out=16'h1c;
17'hd4db:	data_out=16'h89fd;
17'hd4dc:	data_out=16'h8a00;
17'hd4dd:	data_out=16'h8a00;
17'hd4de:	data_out=16'h8a00;
17'hd4df:	data_out=16'h8a00;
17'hd4e0:	data_out=16'ha00;
17'hd4e1:	data_out=16'h8a00;
17'hd4e2:	data_out=16'h9ff;
17'hd4e3:	data_out=16'h871c;
17'hd4e4:	data_out=16'h9e5;
17'hd4e5:	data_out=16'h89d3;
17'hd4e6:	data_out=16'ha00;
17'hd4e7:	data_out=16'h89fb;
17'hd4e8:	data_out=16'h8a00;
17'hd4e9:	data_out=16'h9d8;
17'hd4ea:	data_out=16'h8a00;
17'hd4eb:	data_out=16'h8a00;
17'hd4ec:	data_out=16'h8a00;
17'hd4ed:	data_out=16'h8804;
17'hd4ee:	data_out=16'h8a00;
17'hd4ef:	data_out=16'h89ef;
17'hd4f0:	data_out=16'h8a00;
17'hd4f1:	data_out=16'h89f9;
17'hd4f2:	data_out=16'h8a00;
17'hd4f3:	data_out=16'h8a00;
17'hd4f4:	data_out=16'h89b1;
17'hd4f5:	data_out=16'h8a00;
17'hd4f6:	data_out=16'ha00;
17'hd4f7:	data_out=16'h9ec;
17'hd4f8:	data_out=16'h8a00;
17'hd4f9:	data_out=16'h8a00;
17'hd4fa:	data_out=16'h86cb;
17'hd4fb:	data_out=16'h8a00;
17'hd4fc:	data_out=16'h8a00;
17'hd4fd:	data_out=16'h8871;
17'hd4fe:	data_out=16'h9cd;
17'hd4ff:	data_out=16'h8a00;
17'hd500:	data_out=16'h8a00;
17'hd501:	data_out=16'h8a00;
17'hd502:	data_out=16'h8a00;
17'hd503:	data_out=16'h83c7;
17'hd504:	data_out=16'h8980;
17'hd505:	data_out=16'h8a00;
17'hd506:	data_out=16'h9fa;
17'hd507:	data_out=16'ha00;
17'hd508:	data_out=16'h89ff;
17'hd509:	data_out=16'ha00;
17'hd50a:	data_out=16'h89f4;
17'hd50b:	data_out=16'ha00;
17'hd50c:	data_out=16'ha00;
17'hd50d:	data_out=16'h84a8;
17'hd50e:	data_out=16'h8a00;
17'hd50f:	data_out=16'h81da;
17'hd510:	data_out=16'h976;
17'hd511:	data_out=16'h8a00;
17'hd512:	data_out=16'h696;
17'hd513:	data_out=16'h9f6;
17'hd514:	data_out=16'h365;
17'hd515:	data_out=16'h8a00;
17'hd516:	data_out=16'h8a00;
17'hd517:	data_out=16'h7a0;
17'hd518:	data_out=16'h8a00;
17'hd519:	data_out=16'h9ce;
17'hd51a:	data_out=16'h8a00;
17'hd51b:	data_out=16'h81ea;
17'hd51c:	data_out=16'h8a00;
17'hd51d:	data_out=16'h8a00;
17'hd51e:	data_out=16'h8941;
17'hd51f:	data_out=16'h975;
17'hd520:	data_out=16'h8a00;
17'hd521:	data_out=16'h8a00;
17'hd522:	data_out=16'h427;
17'hd523:	data_out=16'ha00;
17'hd524:	data_out=16'ha00;
17'hd525:	data_out=16'h9e0;
17'hd526:	data_out=16'ha00;
17'hd527:	data_out=16'h89f6;
17'hd528:	data_out=16'h8a00;
17'hd529:	data_out=16'h8a00;
17'hd52a:	data_out=16'h19c;
17'hd52b:	data_out=16'ha00;
17'hd52c:	data_out=16'h8a00;
17'hd52d:	data_out=16'ha00;
17'hd52e:	data_out=16'h4a1;
17'hd52f:	data_out=16'h8a00;
17'hd530:	data_out=16'h877b;
17'hd531:	data_out=16'h8a00;
17'hd532:	data_out=16'h8a00;
17'hd533:	data_out=16'h89c8;
17'hd534:	data_out=16'h8a00;
17'hd535:	data_out=16'h8728;
17'hd536:	data_out=16'h89ff;
17'hd537:	data_out=16'h8a00;
17'hd538:	data_out=16'h8a00;
17'hd539:	data_out=16'h89fe;
17'hd53a:	data_out=16'ha00;
17'hd53b:	data_out=16'h905;
17'hd53c:	data_out=16'h8a00;
17'hd53d:	data_out=16'h8a00;
17'hd53e:	data_out=16'h8a00;
17'hd53f:	data_out=16'h8a00;
17'hd540:	data_out=16'h8a00;
17'hd541:	data_out=16'h8a00;
17'hd542:	data_out=16'ha00;
17'hd543:	data_out=16'h541;
17'hd544:	data_out=16'h8a00;
17'hd545:	data_out=16'h8a00;
17'hd546:	data_out=16'h8a00;
17'hd547:	data_out=16'ha00;
17'hd548:	data_out=16'h9de;
17'hd549:	data_out=16'h9e8;
17'hd54a:	data_out=16'h94b;
17'hd54b:	data_out=16'ha00;
17'hd54c:	data_out=16'h975;
17'hd54d:	data_out=16'h243;
17'hd54e:	data_out=16'h85f8;
17'hd54f:	data_out=16'ha00;
17'hd550:	data_out=16'h8a00;
17'hd551:	data_out=16'h297;
17'hd552:	data_out=16'ha00;
17'hd553:	data_out=16'h8a00;
17'hd554:	data_out=16'h8a00;
17'hd555:	data_out=16'h9cf;
17'hd556:	data_out=16'h985;
17'hd557:	data_out=16'h8a00;
17'hd558:	data_out=16'h8a00;
17'hd559:	data_out=16'h8a00;
17'hd55a:	data_out=16'h82db;
17'hd55b:	data_out=16'h89e7;
17'hd55c:	data_out=16'h8a00;
17'hd55d:	data_out=16'h8a00;
17'hd55e:	data_out=16'h8a00;
17'hd55f:	data_out=16'h89ff;
17'hd560:	data_out=16'ha00;
17'hd561:	data_out=16'h8a00;
17'hd562:	data_out=16'h9f1;
17'hd563:	data_out=16'h89fe;
17'hd564:	data_out=16'h89ec;
17'hd565:	data_out=16'h89cf;
17'hd566:	data_out=16'ha00;
17'hd567:	data_out=16'h9f1;
17'hd568:	data_out=16'h8a00;
17'hd569:	data_out=16'h9a9;
17'hd56a:	data_out=16'h8a00;
17'hd56b:	data_out=16'h8a00;
17'hd56c:	data_out=16'h8a00;
17'hd56d:	data_out=16'h89fe;
17'hd56e:	data_out=16'h8a00;
17'hd56f:	data_out=16'h8a00;
17'hd570:	data_out=16'h8a00;
17'hd571:	data_out=16'h8c0;
17'hd572:	data_out=16'h8a00;
17'hd573:	data_out=16'h8a00;
17'hd574:	data_out=16'h874b;
17'hd575:	data_out=16'h8a00;
17'hd576:	data_out=16'ha00;
17'hd577:	data_out=16'h9e5;
17'hd578:	data_out=16'h8a00;
17'hd579:	data_out=16'h8a00;
17'hd57a:	data_out=16'h8646;
17'hd57b:	data_out=16'h8a00;
17'hd57c:	data_out=16'h8a00;
17'hd57d:	data_out=16'h85fc;
17'hd57e:	data_out=16'h9ec;
17'hd57f:	data_out=16'h8a00;
17'hd580:	data_out=16'h8a00;
17'hd581:	data_out=16'h8a00;
17'hd582:	data_out=16'h89fe;
17'hd583:	data_out=16'h853b;
17'hd584:	data_out=16'h89e4;
17'hd585:	data_out=16'h8a00;
17'hd586:	data_out=16'h9dd;
17'hd587:	data_out=16'ha00;
17'hd588:	data_out=16'h8a00;
17'hd589:	data_out=16'ha00;
17'hd58a:	data_out=16'h89d7;
17'hd58b:	data_out=16'ha00;
17'hd58c:	data_out=16'ha00;
17'hd58d:	data_out=16'h847f;
17'hd58e:	data_out=16'h8a00;
17'hd58f:	data_out=16'h81d3;
17'hd590:	data_out=16'h883;
17'hd591:	data_out=16'h89fe;
17'hd592:	data_out=16'h2aa;
17'hd593:	data_out=16'h9b5;
17'hd594:	data_out=16'h74a;
17'hd595:	data_out=16'h8a00;
17'hd596:	data_out=16'h89fe;
17'hd597:	data_out=16'h597;
17'hd598:	data_out=16'h875d;
17'hd599:	data_out=16'h9ff;
17'hd59a:	data_out=16'h8a00;
17'hd59b:	data_out=16'h8343;
17'hd59c:	data_out=16'h8a00;
17'hd59d:	data_out=16'h8a00;
17'hd59e:	data_out=16'h8904;
17'hd59f:	data_out=16'h9ad;
17'hd5a0:	data_out=16'h8a00;
17'hd5a1:	data_out=16'h89ff;
17'hd5a2:	data_out=16'h8;
17'hd5a3:	data_out=16'ha00;
17'hd5a4:	data_out=16'ha00;
17'hd5a5:	data_out=16'h9bf;
17'hd5a6:	data_out=16'ha00;
17'hd5a7:	data_out=16'h89e4;
17'hd5a8:	data_out=16'h8a00;
17'hd5a9:	data_out=16'h8a00;
17'hd5aa:	data_out=16'h8846;
17'hd5ab:	data_out=16'ha00;
17'hd5ac:	data_out=16'h89fe;
17'hd5ad:	data_out=16'h9ff;
17'hd5ae:	data_out=16'h4e4;
17'hd5af:	data_out=16'h8a00;
17'hd5b0:	data_out=16'h83d7;
17'hd5b1:	data_out=16'h8a00;
17'hd5b2:	data_out=16'h8a00;
17'hd5b3:	data_out=16'h89f9;
17'hd5b4:	data_out=16'h8a00;
17'hd5b5:	data_out=16'h450;
17'hd5b6:	data_out=16'h8a00;
17'hd5b7:	data_out=16'h88c6;
17'hd5b8:	data_out=16'h8a00;
17'hd5b9:	data_out=16'h89fb;
17'hd5ba:	data_out=16'ha00;
17'hd5bb:	data_out=16'h9ff;
17'hd5bc:	data_out=16'h8a00;
17'hd5bd:	data_out=16'h8a00;
17'hd5be:	data_out=16'h8a00;
17'hd5bf:	data_out=16'h8a00;
17'hd5c0:	data_out=16'h89ff;
17'hd5c1:	data_out=16'h8a00;
17'hd5c2:	data_out=16'ha00;
17'hd5c3:	data_out=16'h81ed;
17'hd5c4:	data_out=16'h86f4;
17'hd5c5:	data_out=16'h8a00;
17'hd5c6:	data_out=16'h8a00;
17'hd5c7:	data_out=16'ha00;
17'hd5c8:	data_out=16'h8ec;
17'hd5c9:	data_out=16'h9d7;
17'hd5ca:	data_out=16'h4e6;
17'hd5cb:	data_out=16'ha00;
17'hd5cc:	data_out=16'h954;
17'hd5cd:	data_out=16'h827b;
17'hd5ce:	data_out=16'h89f2;
17'hd5cf:	data_out=16'ha00;
17'hd5d0:	data_out=16'h89fc;
17'hd5d1:	data_out=16'h970;
17'hd5d2:	data_out=16'ha00;
17'hd5d3:	data_out=16'h8a00;
17'hd5d4:	data_out=16'h8a00;
17'hd5d5:	data_out=16'h9e1;
17'hd5d6:	data_out=16'h9d7;
17'hd5d7:	data_out=16'h454;
17'hd5d8:	data_out=16'h89ff;
17'hd5d9:	data_out=16'h8a00;
17'hd5da:	data_out=16'h894c;
17'hd5db:	data_out=16'h89d5;
17'hd5dc:	data_out=16'h8a00;
17'hd5dd:	data_out=16'h8a00;
17'hd5de:	data_out=16'h8a00;
17'hd5df:	data_out=16'h8a00;
17'hd5e0:	data_out=16'ha00;
17'hd5e1:	data_out=16'h8a00;
17'hd5e2:	data_out=16'h9e7;
17'hd5e3:	data_out=16'h89fb;
17'hd5e4:	data_out=16'h89f5;
17'hd5e5:	data_out=16'h88a1;
17'hd5e6:	data_out=16'ha00;
17'hd5e7:	data_out=16'ha00;
17'hd5e8:	data_out=16'h89ff;
17'hd5e9:	data_out=16'h999;
17'hd5ea:	data_out=16'h8a00;
17'hd5eb:	data_out=16'h8a00;
17'hd5ec:	data_out=16'h8a00;
17'hd5ed:	data_out=16'h89fb;
17'hd5ee:	data_out=16'h8a00;
17'hd5ef:	data_out=16'h89ff;
17'hd5f0:	data_out=16'h8a00;
17'hd5f1:	data_out=16'h6d8;
17'hd5f2:	data_out=16'h8a00;
17'hd5f3:	data_out=16'h8a00;
17'hd5f4:	data_out=16'h83eb;
17'hd5f5:	data_out=16'h8a00;
17'hd5f6:	data_out=16'ha00;
17'hd5f7:	data_out=16'h9bf;
17'hd5f8:	data_out=16'h8a00;
17'hd5f9:	data_out=16'h8a00;
17'hd5fa:	data_out=16'h87a7;
17'hd5fb:	data_out=16'h8a00;
17'hd5fc:	data_out=16'h8a00;
17'hd5fd:	data_out=16'h3b9;
17'hd5fe:	data_out=16'h9ee;
17'hd5ff:	data_out=16'h8a00;
17'hd600:	data_out=16'h8a00;
17'hd601:	data_out=16'h8a00;
17'hd602:	data_out=16'h85d8;
17'hd603:	data_out=16'h82f8;
17'hd604:	data_out=16'h89c5;
17'hd605:	data_out=16'h8a00;
17'hd606:	data_out=16'h9ae;
17'hd607:	data_out=16'ha00;
17'hd608:	data_out=16'h89e9;
17'hd609:	data_out=16'h9e9;
17'hd60a:	data_out=16'h899a;
17'hd60b:	data_out=16'ha00;
17'hd60c:	data_out=16'h9f7;
17'hd60d:	data_out=16'h4ba;
17'hd60e:	data_out=16'h829e;
17'hd60f:	data_out=16'h9f2;
17'hd610:	data_out=16'h7a7;
17'hd611:	data_out=16'h89f1;
17'hd612:	data_out=16'h462;
17'hd613:	data_out=16'h9b6;
17'hd614:	data_out=16'h9a8;
17'hd615:	data_out=16'h89f8;
17'hd616:	data_out=16'h872c;
17'hd617:	data_out=16'h117;
17'hd618:	data_out=16'h85;
17'hd619:	data_out=16'h809a;
17'hd61a:	data_out=16'h89ff;
17'hd61b:	data_out=16'h137;
17'hd61c:	data_out=16'h8a00;
17'hd61d:	data_out=16'h8a00;
17'hd61e:	data_out=16'h82b9;
17'hd61f:	data_out=16'h9d6;
17'hd620:	data_out=16'h8a00;
17'hd621:	data_out=16'h8209;
17'hd622:	data_out=16'h128;
17'hd623:	data_out=16'ha00;
17'hd624:	data_out=16'ha00;
17'hd625:	data_out=16'h9df;
17'hd626:	data_out=16'h9fd;
17'hd627:	data_out=16'h89b4;
17'hd628:	data_out=16'h80b1;
17'hd629:	data_out=16'h2af;
17'hd62a:	data_out=16'h811d;
17'hd62b:	data_out=16'h6d8;
17'hd62c:	data_out=16'h887d;
17'hd62d:	data_out=16'h9fa;
17'hd62e:	data_out=16'h7b4;
17'hd62f:	data_out=16'h8a00;
17'hd630:	data_out=16'h22c;
17'hd631:	data_out=16'h89b0;
17'hd632:	data_out=16'h89f8;
17'hd633:	data_out=16'h88a8;
17'hd634:	data_out=16'h8a00;
17'hd635:	data_out=16'h9fd;
17'hd636:	data_out=16'h89de;
17'hd637:	data_out=16'h312;
17'hd638:	data_out=16'h8a00;
17'hd639:	data_out=16'h89d9;
17'hd63a:	data_out=16'ha00;
17'hd63b:	data_out=16'ha00;
17'hd63c:	data_out=16'h8a00;
17'hd63d:	data_out=16'h89ea;
17'hd63e:	data_out=16'h80a6;
17'hd63f:	data_out=16'h8a00;
17'hd640:	data_out=16'h89fe;
17'hd641:	data_out=16'h89c2;
17'hd642:	data_out=16'h9e9;
17'hd643:	data_out=16'h112;
17'hd644:	data_out=16'h80d5;
17'hd645:	data_out=16'h89f8;
17'hd646:	data_out=16'h8a00;
17'hd647:	data_out=16'ha00;
17'hd648:	data_out=16'h8d0;
17'hd649:	data_out=16'h9f8;
17'hd64a:	data_out=16'h6c;
17'hd64b:	data_out=16'h9e9;
17'hd64c:	data_out=16'h9ce;
17'hd64d:	data_out=16'h8562;
17'hd64e:	data_out=16'h89e7;
17'hd64f:	data_out=16'h9fe;
17'hd650:	data_out=16'h89f7;
17'hd651:	data_out=16'ha00;
17'hd652:	data_out=16'ha00;
17'hd653:	data_out=16'h89d5;
17'hd654:	data_out=16'h8a00;
17'hd655:	data_out=16'ha00;
17'hd656:	data_out=16'h9ff;
17'hd657:	data_out=16'h9ec;
17'hd658:	data_out=16'h89be;
17'hd659:	data_out=16'h89fe;
17'hd65a:	data_out=16'h877c;
17'hd65b:	data_out=16'h896d;
17'hd65c:	data_out=16'h8a00;
17'hd65d:	data_out=16'h8a00;
17'hd65e:	data_out=16'h8a00;
17'hd65f:	data_out=16'h89fc;
17'hd660:	data_out=16'h9f6;
17'hd661:	data_out=16'h89e2;
17'hd662:	data_out=16'h9f3;
17'hd663:	data_out=16'h89cb;
17'hd664:	data_out=16'h8a00;
17'hd665:	data_out=16'h8a00;
17'hd666:	data_out=16'ha00;
17'hd667:	data_out=16'ha00;
17'hd668:	data_out=16'h8123;
17'hd669:	data_out=16'h157;
17'hd66a:	data_out=16'h82d7;
17'hd66b:	data_out=16'h89fe;
17'hd66c:	data_out=16'h8a00;
17'hd66d:	data_out=16'h89da;
17'hd66e:	data_out=16'h82da;
17'hd66f:	data_out=16'h89f8;
17'hd670:	data_out=16'h82cb;
17'hd671:	data_out=16'h9e9;
17'hd672:	data_out=16'h8a00;
17'hd673:	data_out=16'h8a00;
17'hd674:	data_out=16'h248;
17'hd675:	data_out=16'h8a00;
17'hd676:	data_out=16'ha00;
17'hd677:	data_out=16'h9b0;
17'hd678:	data_out=16'h8a00;
17'hd679:	data_out=16'h8a00;
17'hd67a:	data_out=16'h857c;
17'hd67b:	data_out=16'h80a6;
17'hd67c:	data_out=16'h89f5;
17'hd67d:	data_out=16'h9a9;
17'hd67e:	data_out=16'h9d9;
17'hd67f:	data_out=16'h8a00;
17'hd680:	data_out=16'h8a00;
17'hd681:	data_out=16'h89fe;
17'hd682:	data_out=16'h151;
17'hd683:	data_out=16'h81f0;
17'hd684:	data_out=16'h895f;
17'hd685:	data_out=16'h8951;
17'hd686:	data_out=16'h9c7;
17'hd687:	data_out=16'ha00;
17'hd688:	data_out=16'h89b0;
17'hd689:	data_out=16'ha00;
17'hd68a:	data_out=16'h89dd;
17'hd68b:	data_out=16'ha00;
17'hd68c:	data_out=16'h9fe;
17'hd68d:	data_out=16'h8198;
17'hd68e:	data_out=16'ha00;
17'hd68f:	data_out=16'h9e9;
17'hd690:	data_out=16'h87d;
17'hd691:	data_out=16'h884c;
17'hd692:	data_out=16'h89bb;
17'hd693:	data_out=16'h814a;
17'hd694:	data_out=16'h235;
17'hd695:	data_out=16'h89de;
17'hd696:	data_out=16'h8420;
17'hd697:	data_out=16'h8281;
17'hd698:	data_out=16'h87;
17'hd699:	data_out=16'h89fc;
17'hd69a:	data_out=16'h8976;
17'hd69b:	data_out=16'h3b3;
17'hd69c:	data_out=16'h89dc;
17'hd69d:	data_out=16'h8a00;
17'hd69e:	data_out=16'h8140;
17'hd69f:	data_out=16'h9f4;
17'hd6a0:	data_out=16'h89e3;
17'hd6a1:	data_out=16'ha00;
17'hd6a2:	data_out=16'h88c;
17'hd6a3:	data_out=16'ha00;
17'hd6a4:	data_out=16'ha00;
17'hd6a5:	data_out=16'h9ff;
17'hd6a6:	data_out=16'h9fb;
17'hd6a7:	data_out=16'h8980;
17'hd6a8:	data_out=16'ha00;
17'hd6a9:	data_out=16'h8c5;
17'hd6aa:	data_out=16'h3cc;
17'hd6ab:	data_out=16'h330;
17'hd6ac:	data_out=16'h857d;
17'hd6ad:	data_out=16'h9bd;
17'hd6ae:	data_out=16'h52c;
17'hd6af:	data_out=16'h89c9;
17'hd6b0:	data_out=16'ha00;
17'hd6b1:	data_out=16'h8215;
17'hd6b2:	data_out=16'h8959;
17'hd6b3:	data_out=16'h8708;
17'hd6b4:	data_out=16'h8a00;
17'hd6b5:	data_out=16'h9ff;
17'hd6b6:	data_out=16'h8989;
17'hd6b7:	data_out=16'h6c1;
17'hd6b8:	data_out=16'h8a00;
17'hd6b9:	data_out=16'h892a;
17'hd6ba:	data_out=16'ha00;
17'hd6bb:	data_out=16'ha00;
17'hd6bc:	data_out=16'h8a00;
17'hd6bd:	data_out=16'h89cc;
17'hd6be:	data_out=16'ha00;
17'hd6bf:	data_out=16'h8953;
17'hd6c0:	data_out=16'h8977;
17'hd6c1:	data_out=16'h8956;
17'hd6c2:	data_out=16'h9d7;
17'hd6c3:	data_out=16'h85f4;
17'hd6c4:	data_out=16'ha00;
17'hd6c5:	data_out=16'h89dd;
17'hd6c6:	data_out=16'h8a00;
17'hd6c7:	data_out=16'h9d0;
17'hd6c8:	data_out=16'h933;
17'hd6c9:	data_out=16'ha00;
17'hd6ca:	data_out=16'h4e6;
17'hd6cb:	data_out=16'h9e7;
17'hd6cc:	data_out=16'h9df;
17'hd6cd:	data_out=16'h84ad;
17'hd6ce:	data_out=16'h89ee;
17'hd6cf:	data_out=16'h9fb;
17'hd6d0:	data_out=16'h8738;
17'hd6d1:	data_out=16'ha00;
17'hd6d2:	data_out=16'h9ff;
17'hd6d3:	data_out=16'h897e;
17'hd6d4:	data_out=16'h89e7;
17'hd6d5:	data_out=16'ha00;
17'hd6d6:	data_out=16'h9f1;
17'hd6d7:	data_out=16'h9d2;
17'hd6d8:	data_out=16'h87a4;
17'hd6d9:	data_out=16'h89d1;
17'hd6da:	data_out=16'h8761;
17'hd6db:	data_out=16'h84e4;
17'hd6dc:	data_out=16'h89bb;
17'hd6dd:	data_out=16'h89cb;
17'hd6de:	data_out=16'h89a5;
17'hd6df:	data_out=16'h89fb;
17'hd6e0:	data_out=16'h9ea;
17'hd6e1:	data_out=16'h8517;
17'hd6e2:	data_out=16'h72d;
17'hd6e3:	data_out=16'h880f;
17'hd6e4:	data_out=16'h8a00;
17'hd6e5:	data_out=16'h86bb;
17'hd6e6:	data_out=16'ha00;
17'hd6e7:	data_out=16'ha00;
17'hd6e8:	data_out=16'ha00;
17'hd6e9:	data_out=16'h89cb;
17'hd6ea:	data_out=16'ha00;
17'hd6eb:	data_out=16'h89c0;
17'hd6ec:	data_out=16'h8a00;
17'hd6ed:	data_out=16'h8827;
17'hd6ee:	data_out=16'ha00;
17'hd6ef:	data_out=16'h87bf;
17'hd6f0:	data_out=16'ha00;
17'hd6f1:	data_out=16'hf7;
17'hd6f2:	data_out=16'h8a00;
17'hd6f3:	data_out=16'h89d7;
17'hd6f4:	data_out=16'h9fe;
17'hd6f5:	data_out=16'h89a7;
17'hd6f6:	data_out=16'ha00;
17'hd6f7:	data_out=16'h9fa;
17'hd6f8:	data_out=16'h8a00;
17'hd6f9:	data_out=16'h89fc;
17'hd6fa:	data_out=16'h8480;
17'hd6fb:	data_out=16'ha00;
17'hd6fc:	data_out=16'h89ed;
17'hd6fd:	data_out=16'h9ff;
17'hd6fe:	data_out=16'h9e9;
17'hd6ff:	data_out=16'h8a00;
17'hd700:	data_out=16'h8a00;
17'hd701:	data_out=16'h8a00;
17'hd702:	data_out=16'h86a8;
17'hd703:	data_out=16'h88cf;
17'hd704:	data_out=16'h80c8;
17'hd705:	data_out=16'h894d;
17'hd706:	data_out=16'h9a9;
17'hd707:	data_out=16'ha00;
17'hd708:	data_out=16'h89c0;
17'hd709:	data_out=16'ha00;
17'hd70a:	data_out=16'h8a00;
17'hd70b:	data_out=16'ha00;
17'hd70c:	data_out=16'ha00;
17'hd70d:	data_out=16'h892a;
17'hd70e:	data_out=16'ha00;
17'hd70f:	data_out=16'h8544;
17'hd710:	data_out=16'h8636;
17'hd711:	data_out=16'h3ca;
17'hd712:	data_out=16'h89f7;
17'hd713:	data_out=16'h8a00;
17'hd714:	data_out=16'h8997;
17'hd715:	data_out=16'h89ea;
17'hd716:	data_out=16'h896c;
17'hd717:	data_out=16'h89a8;
17'hd718:	data_out=16'h89f9;
17'hd719:	data_out=16'h8a00;
17'hd71a:	data_out=16'h8986;
17'hd71b:	data_out=16'h8695;
17'hd71c:	data_out=16'h89d2;
17'hd71d:	data_out=16'h8a00;
17'hd71e:	data_out=16'h896e;
17'hd71f:	data_out=16'h94c;
17'hd720:	data_out=16'h89f9;
17'hd721:	data_out=16'ha00;
17'hd722:	data_out=16'h9ea;
17'hd723:	data_out=16'ha00;
17'hd724:	data_out=16'ha00;
17'hd725:	data_out=16'ha00;
17'hd726:	data_out=16'h9f6;
17'hd727:	data_out=16'h89e4;
17'hd728:	data_out=16'ha00;
17'hd729:	data_out=16'h810a;
17'hd72a:	data_out=16'h8707;
17'hd72b:	data_out=16'h89db;
17'hd72c:	data_out=16'h8986;
17'hd72d:	data_out=16'h995;
17'hd72e:	data_out=16'h89d3;
17'hd72f:	data_out=16'h89ea;
17'hd730:	data_out=16'h9fe;
17'hd731:	data_out=16'h89cb;
17'hd732:	data_out=16'h8572;
17'hd733:	data_out=16'h89db;
17'hd734:	data_out=16'h8a00;
17'hd735:	data_out=16'h9fd;
17'hd736:	data_out=16'h89c1;
17'hd737:	data_out=16'h8647;
17'hd738:	data_out=16'h8a00;
17'hd739:	data_out=16'h89eb;
17'hd73a:	data_out=16'h9fd;
17'hd73b:	data_out=16'ha00;
17'hd73c:	data_out=16'h8a00;
17'hd73d:	data_out=16'h89ee;
17'hd73e:	data_out=16'ha00;
17'hd73f:	data_out=16'h894e;
17'hd740:	data_out=16'h897d;
17'hd741:	data_out=16'h8957;
17'hd742:	data_out=16'ha00;
17'hd743:	data_out=16'h889d;
17'hd744:	data_out=16'h9ff;
17'hd745:	data_out=16'h89e9;
17'hd746:	data_out=16'h8a00;
17'hd747:	data_out=16'h981;
17'hd748:	data_out=16'h89e9;
17'hd749:	data_out=16'ha00;
17'hd74a:	data_out=16'h8933;
17'hd74b:	data_out=16'ha00;
17'hd74c:	data_out=16'h9ed;
17'hd74d:	data_out=16'h80;
17'hd74e:	data_out=16'h8a00;
17'hd74f:	data_out=16'ha00;
17'hd750:	data_out=16'h88c2;
17'hd751:	data_out=16'h8329;
17'hd752:	data_out=16'ha00;
17'hd753:	data_out=16'h89d3;
17'hd754:	data_out=16'h89ff;
17'hd755:	data_out=16'h90c;
17'hd756:	data_out=16'h8263;
17'hd757:	data_out=16'h9d4;
17'hd758:	data_out=16'h8976;
17'hd759:	data_out=16'h89f8;
17'hd75a:	data_out=16'h89b2;
17'hd75b:	data_out=16'h89a9;
17'hd75c:	data_out=16'h89d3;
17'hd75d:	data_out=16'h89df;
17'hd75e:	data_out=16'h89a4;
17'hd75f:	data_out=16'h8a00;
17'hd760:	data_out=16'h9eb;
17'hd761:	data_out=16'h835c;
17'hd762:	data_out=16'h8914;
17'hd763:	data_out=16'h89d5;
17'hd764:	data_out=16'h8a00;
17'hd765:	data_out=16'h89f7;
17'hd766:	data_out=16'ha00;
17'hd767:	data_out=16'h5b9;
17'hd768:	data_out=16'ha00;
17'hd769:	data_out=16'h89bc;
17'hd76a:	data_out=16'ha00;
17'hd76b:	data_out=16'h89e2;
17'hd76c:	data_out=16'h8a00;
17'hd76d:	data_out=16'h89d8;
17'hd76e:	data_out=16'ha00;
17'hd76f:	data_out=16'h8980;
17'hd770:	data_out=16'ha00;
17'hd771:	data_out=16'h89c6;
17'hd772:	data_out=16'h8a00;
17'hd773:	data_out=16'h8a00;
17'hd774:	data_out=16'h9fd;
17'hd775:	data_out=16'h8922;
17'hd776:	data_out=16'h9e5;
17'hd777:	data_out=16'ha00;
17'hd778:	data_out=16'h8a00;
17'hd779:	data_out=16'h89fa;
17'hd77a:	data_out=16'h89c1;
17'hd77b:	data_out=16'ha00;
17'hd77c:	data_out=16'h89fd;
17'hd77d:	data_out=16'h9fe;
17'hd77e:	data_out=16'ha00;
17'hd77f:	data_out=16'h89ff;
17'hd780:	data_out=16'h8a00;
17'hd781:	data_out=16'h8a00;
17'hd782:	data_out=16'h899c;
17'hd783:	data_out=16'h898f;
17'hd784:	data_out=16'h61d;
17'hd785:	data_out=16'h9d9;
17'hd786:	data_out=16'h9e6;
17'hd787:	data_out=16'h9fb;
17'hd788:	data_out=16'h8a00;
17'hd789:	data_out=16'ha00;
17'hd78a:	data_out=16'h8a00;
17'hd78b:	data_out=16'h89b9;
17'hd78c:	data_out=16'h19d;
17'hd78d:	data_out=16'h89bb;
17'hd78e:	data_out=16'ha00;
17'hd78f:	data_out=16'h89af;
17'hd790:	data_out=16'h8867;
17'hd791:	data_out=16'h443;
17'hd792:	data_out=16'h8a00;
17'hd793:	data_out=16'h8a00;
17'hd794:	data_out=16'h89bf;
17'hd795:	data_out=16'h89f9;
17'hd796:	data_out=16'h89e0;
17'hd797:	data_out=16'h89b8;
17'hd798:	data_out=16'h89fd;
17'hd799:	data_out=16'h8a00;
17'hd79a:	data_out=16'h684;
17'hd79b:	data_out=16'h89c9;
17'hd79c:	data_out=16'h89ca;
17'hd79d:	data_out=16'h8a00;
17'hd79e:	data_out=16'h89dc;
17'hd79f:	data_out=16'h8153;
17'hd7a0:	data_out=16'h89f6;
17'hd7a1:	data_out=16'ha00;
17'hd7a2:	data_out=16'ha00;
17'hd7a3:	data_out=16'ha00;
17'hd7a4:	data_out=16'ha00;
17'hd7a5:	data_out=16'ha00;
17'hd7a6:	data_out=16'h89c0;
17'hd7a7:	data_out=16'h89f9;
17'hd7a8:	data_out=16'ha00;
17'hd7a9:	data_out=16'h89e7;
17'hd7aa:	data_out=16'h899c;
17'hd7ab:	data_out=16'h8a00;
17'hd7ac:	data_out=16'h89d5;
17'hd7ad:	data_out=16'h81b;
17'hd7ae:	data_out=16'h89d0;
17'hd7af:	data_out=16'h8a00;
17'hd7b0:	data_out=16'h9fc;
17'hd7b1:	data_out=16'h89fe;
17'hd7b2:	data_out=16'h8060;
17'hd7b3:	data_out=16'h89e6;
17'hd7b4:	data_out=16'h8a00;
17'hd7b5:	data_out=16'h89ef;
17'hd7b6:	data_out=16'h89ff;
17'hd7b7:	data_out=16'h89a4;
17'hd7b8:	data_out=16'h89ff;
17'hd7b9:	data_out=16'h89fb;
17'hd7ba:	data_out=16'h827b;
17'hd7bb:	data_out=16'ha00;
17'hd7bc:	data_out=16'h8a00;
17'hd7bd:	data_out=16'h89ea;
17'hd7be:	data_out=16'ha00;
17'hd7bf:	data_out=16'h9d9;
17'hd7c0:	data_out=16'h8729;
17'hd7c1:	data_out=16'h89e2;
17'hd7c2:	data_out=16'h4c4;
17'hd7c3:	data_out=16'h9fe;
17'hd7c4:	data_out=16'h81be;
17'hd7c5:	data_out=16'h89f9;
17'hd7c6:	data_out=16'h8a00;
17'hd7c7:	data_out=16'h89f8;
17'hd7c8:	data_out=16'h89e8;
17'hd7c9:	data_out=16'ha00;
17'hd7ca:	data_out=16'h89f6;
17'hd7cb:	data_out=16'h727;
17'hd7cc:	data_out=16'h9fd;
17'hd7cd:	data_out=16'h8c9;
17'hd7ce:	data_out=16'h8a00;
17'hd7cf:	data_out=16'ha00;
17'hd7d0:	data_out=16'h87f0;
17'hd7d1:	data_out=16'h8781;
17'hd7d2:	data_out=16'ha00;
17'hd7d3:	data_out=16'h89ff;
17'hd7d4:	data_out=16'h89fe;
17'hd7d5:	data_out=16'h895f;
17'hd7d6:	data_out=16'h89f8;
17'hd7d7:	data_out=16'h9c4;
17'hd7d8:	data_out=16'h8991;
17'hd7d9:	data_out=16'h71b;
17'hd7da:	data_out=16'h89de;
17'hd7db:	data_out=16'h89ec;
17'hd7dc:	data_out=16'h89f1;
17'hd7dd:	data_out=16'h89bd;
17'hd7de:	data_out=16'h88d4;
17'hd7df:	data_out=16'h8a00;
17'hd7e0:	data_out=16'h8986;
17'hd7e1:	data_out=16'h844;
17'hd7e2:	data_out=16'h89cb;
17'hd7e3:	data_out=16'h89ea;
17'hd7e4:	data_out=16'h8a00;
17'hd7e5:	data_out=16'h89fc;
17'hd7e6:	data_out=16'h9fe;
17'hd7e7:	data_out=16'h89e7;
17'hd7e8:	data_out=16'ha00;
17'hd7e9:	data_out=16'h8a00;
17'hd7ea:	data_out=16'ha00;
17'hd7eb:	data_out=16'h8931;
17'hd7ec:	data_out=16'h8a00;
17'hd7ed:	data_out=16'h89ec;
17'hd7ee:	data_out=16'ha00;
17'hd7ef:	data_out=16'h89a9;
17'hd7f0:	data_out=16'ha00;
17'hd7f1:	data_out=16'h89ec;
17'hd7f2:	data_out=16'h83bb;
17'hd7f3:	data_out=16'h8202;
17'hd7f4:	data_out=16'h9f0;
17'hd7f5:	data_out=16'h9fa;
17'hd7f6:	data_out=16'h854a;
17'hd7f7:	data_out=16'h86da;
17'hd7f8:	data_out=16'h7f5;
17'hd7f9:	data_out=16'h8a00;
17'hd7fa:	data_out=16'h89d5;
17'hd7fb:	data_out=16'ha00;
17'hd7fc:	data_out=16'h89fe;
17'hd7fd:	data_out=16'h9ff;
17'hd7fe:	data_out=16'ha00;
17'hd7ff:	data_out=16'h4f1;
17'hd800:	data_out=16'h89ff;
17'hd801:	data_out=16'h89ff;
17'hd802:	data_out=16'h899d;
17'hd803:	data_out=16'h8935;
17'hd804:	data_out=16'h9e5;
17'hd805:	data_out=16'ha00;
17'hd806:	data_out=16'h9dd;
17'hd807:	data_out=16'h8a00;
17'hd808:	data_out=16'h8a00;
17'hd809:	data_out=16'h87f5;
17'hd80a:	data_out=16'h8a00;
17'hd80b:	data_out=16'h89f0;
17'hd80c:	data_out=16'h8a00;
17'hd80d:	data_out=16'h8a00;
17'hd80e:	data_out=16'ha00;
17'hd80f:	data_out=16'h89ff;
17'hd810:	data_out=16'h88e1;
17'hd811:	data_out=16'h9c6;
17'hd812:	data_out=16'h8a00;
17'hd813:	data_out=16'h89e1;
17'hd814:	data_out=16'h89ac;
17'hd815:	data_out=16'h8946;
17'hd816:	data_out=16'h89df;
17'hd817:	data_out=16'h89b2;
17'hd818:	data_out=16'h89ff;
17'hd819:	data_out=16'h89fd;
17'hd81a:	data_out=16'ha00;
17'hd81b:	data_out=16'h89f0;
17'hd81c:	data_out=16'h552;
17'hd81d:	data_out=16'h8a00;
17'hd81e:	data_out=16'h899e;
17'hd81f:	data_out=16'h9fa;
17'hd820:	data_out=16'h89c4;
17'hd821:	data_out=16'ha00;
17'hd822:	data_out=16'ha00;
17'hd823:	data_out=16'h8590;
17'hd824:	data_out=16'h8587;
17'hd825:	data_out=16'ha00;
17'hd826:	data_out=16'h8a00;
17'hd827:	data_out=16'h89f8;
17'hd828:	data_out=16'ha00;
17'hd829:	data_out=16'h8a00;
17'hd82a:	data_out=16'h89fb;
17'hd82b:	data_out=16'h8a00;
17'hd82c:	data_out=16'h892c;
17'hd82d:	data_out=16'h70d;
17'hd82e:	data_out=16'h89e1;
17'hd82f:	data_out=16'h89ee;
17'hd830:	data_out=16'h9f0;
17'hd831:	data_out=16'h8787;
17'hd832:	data_out=16'h9e5;
17'hd833:	data_out=16'h89d0;
17'hd834:	data_out=16'h8a00;
17'hd835:	data_out=16'h89bc;
17'hd836:	data_out=16'h89ff;
17'hd837:	data_out=16'h899d;
17'hd838:	data_out=16'h9f8;
17'hd839:	data_out=16'h89e3;
17'hd83a:	data_out=16'h89fb;
17'hd83b:	data_out=16'h81b9;
17'hd83c:	data_out=16'h89fd;
17'hd83d:	data_out=16'h85bb;
17'hd83e:	data_out=16'ha00;
17'hd83f:	data_out=16'ha00;
17'hd840:	data_out=16'h9e8;
17'hd841:	data_out=16'h8a00;
17'hd842:	data_out=16'h89d3;
17'hd843:	data_out=16'ha00;
17'hd844:	data_out=16'h430;
17'hd845:	data_out=16'h894c;
17'hd846:	data_out=16'h8a00;
17'hd847:	data_out=16'h8a00;
17'hd848:	data_out=16'h89fc;
17'hd849:	data_out=16'ha00;
17'hd84a:	data_out=16'h8a00;
17'hd84b:	data_out=16'h89be;
17'hd84c:	data_out=16'h9f5;
17'hd84d:	data_out=16'ha00;
17'hd84e:	data_out=16'h8a00;
17'hd84f:	data_out=16'h85b4;
17'hd850:	data_out=16'h9fe;
17'hd851:	data_out=16'h9c4;
17'hd852:	data_out=16'h8544;
17'hd853:	data_out=16'h89e3;
17'hd854:	data_out=16'h89f0;
17'hd855:	data_out=16'h89a3;
17'hd856:	data_out=16'h89fd;
17'hd857:	data_out=16'h9da;
17'hd858:	data_out=16'h89ab;
17'hd859:	data_out=16'h9cb;
17'hd85a:	data_out=16'h89f4;
17'hd85b:	data_out=16'h9c1;
17'hd85c:	data_out=16'h897e;
17'hd85d:	data_out=16'h86fb;
17'hd85e:	data_out=16'h8677;
17'hd85f:	data_out=16'h89ff;
17'hd860:	data_out=16'h8a00;
17'hd861:	data_out=16'h9ff;
17'hd862:	data_out=16'h89db;
17'hd863:	data_out=16'h89d8;
17'hd864:	data_out=16'h8a00;
17'hd865:	data_out=16'h89f3;
17'hd866:	data_out=16'h89a7;
17'hd867:	data_out=16'h89b5;
17'hd868:	data_out=16'ha00;
17'hd869:	data_out=16'h8a00;
17'hd86a:	data_out=16'ha00;
17'hd86b:	data_out=16'ha00;
17'hd86c:	data_out=16'h89ff;
17'hd86d:	data_out=16'h89d9;
17'hd86e:	data_out=16'ha00;
17'hd86f:	data_out=16'h8e9;
17'hd870:	data_out=16'ha00;
17'hd871:	data_out=16'h8a00;
17'hd872:	data_out=16'h9d7;
17'hd873:	data_out=16'h9d5;
17'hd874:	data_out=16'h9e6;
17'hd875:	data_out=16'ha00;
17'hd876:	data_out=16'h89f5;
17'hd877:	data_out=16'h896b;
17'hd878:	data_out=16'ha00;
17'hd879:	data_out=16'h8a00;
17'hd87a:	data_out=16'h89cc;
17'hd87b:	data_out=16'ha00;
17'hd87c:	data_out=16'h89ff;
17'hd87d:	data_out=16'h9ff;
17'hd87e:	data_out=16'ha00;
17'hd87f:	data_out=16'ha00;
17'hd880:	data_out=16'h89fc;
17'hd881:	data_out=16'h89ed;
17'hd882:	data_out=16'h89e3;
17'hd883:	data_out=16'h81a5;
17'hd884:	data_out=16'h7eb;
17'hd885:	data_out=16'ha00;
17'hd886:	data_out=16'h9ca;
17'hd887:	data_out=16'h8a00;
17'hd888:	data_out=16'h8a00;
17'hd889:	data_out=16'h8a00;
17'hd88a:	data_out=16'h89c7;
17'hd88b:	data_out=16'h8a00;
17'hd88c:	data_out=16'h8a00;
17'hd88d:	data_out=16'h8a00;
17'hd88e:	data_out=16'ha00;
17'hd88f:	data_out=16'h8a00;
17'hd890:	data_out=16'h898a;
17'hd891:	data_out=16'h9eb;
17'hd892:	data_out=16'h8a00;
17'hd893:	data_out=16'h712;
17'hd894:	data_out=16'h9cf;
17'hd895:	data_out=16'h80e8;
17'hd896:	data_out=16'h862a;
17'hd897:	data_out=16'h494;
17'hd898:	data_out=16'h8a00;
17'hd899:	data_out=16'h89ff;
17'hd89a:	data_out=16'ha00;
17'hd89b:	data_out=16'h89ed;
17'hd89c:	data_out=16'h9fa;
17'hd89d:	data_out=16'h89fb;
17'hd89e:	data_out=16'h9c2;
17'hd89f:	data_out=16'h9fd;
17'hd8a0:	data_out=16'ha00;
17'hd8a1:	data_out=16'ha00;
17'hd8a2:	data_out=16'ha00;
17'hd8a3:	data_out=16'h8a00;
17'hd8a4:	data_out=16'h8a00;
17'hd8a5:	data_out=16'h9eb;
17'hd8a6:	data_out=16'h8a00;
17'hd8a7:	data_out=16'h89ff;
17'hd8a8:	data_out=16'ha00;
17'hd8a9:	data_out=16'h552;
17'hd8aa:	data_out=16'h89e0;
17'hd8ab:	data_out=16'h8a00;
17'hd8ac:	data_out=16'he3;
17'hd8ad:	data_out=16'h299;
17'hd8ae:	data_out=16'h983;
17'hd8af:	data_out=16'h118;
17'hd8b0:	data_out=16'h801;
17'hd8b1:	data_out=16'h8950;
17'hd8b2:	data_out=16'h9ea;
17'hd8b3:	data_out=16'h9f5;
17'hd8b4:	data_out=16'h8a00;
17'hd8b5:	data_out=16'h89ff;
17'hd8b6:	data_out=16'h89ff;
17'hd8b7:	data_out=16'h816a;
17'hd8b8:	data_out=16'ha00;
17'hd8b9:	data_out=16'h9dc;
17'hd8ba:	data_out=16'h8a00;
17'hd8bb:	data_out=16'h8a00;
17'hd8bc:	data_out=16'h9ec;
17'hd8bd:	data_out=16'ha00;
17'hd8be:	data_out=16'ha00;
17'hd8bf:	data_out=16'ha00;
17'hd8c0:	data_out=16'h9f3;
17'hd8c1:	data_out=16'h8a00;
17'hd8c2:	data_out=16'h8a00;
17'hd8c3:	data_out=16'ha00;
17'hd8c4:	data_out=16'h89e6;
17'hd8c5:	data_out=16'h80c2;
17'hd8c6:	data_out=16'h8a00;
17'hd8c7:	data_out=16'h8a00;
17'hd8c8:	data_out=16'h74c;
17'hd8c9:	data_out=16'h996;
17'hd8ca:	data_out=16'h8a00;
17'hd8cb:	data_out=16'h8a00;
17'hd8cc:	data_out=16'h813e;
17'hd8cd:	data_out=16'ha00;
17'hd8ce:	data_out=16'h8a00;
17'hd8cf:	data_out=16'h8a00;
17'hd8d0:	data_out=16'h9fb;
17'hd8d1:	data_out=16'h9a1;
17'hd8d2:	data_out=16'h8a00;
17'hd8d3:	data_out=16'h759;
17'hd8d4:	data_out=16'h391;
17'hd8d5:	data_out=16'h639;
17'hd8d6:	data_out=16'h8a00;
17'hd8d7:	data_out=16'h9dd;
17'hd8d8:	data_out=16'h83b8;
17'hd8d9:	data_out=16'ha00;
17'hd8da:	data_out=16'h89d6;
17'hd8db:	data_out=16'h9e5;
17'hd8dc:	data_out=16'ha00;
17'hd8dd:	data_out=16'h1fa;
17'hd8de:	data_out=16'h5cb;
17'hd8df:	data_out=16'h89fd;
17'hd8e0:	data_out=16'h8a00;
17'hd8e1:	data_out=16'ha00;
17'hd8e2:	data_out=16'h84b1;
17'hd8e3:	data_out=16'h9d6;
17'hd8e4:	data_out=16'h8a00;
17'hd8e5:	data_out=16'h8a00;
17'hd8e6:	data_out=16'h8a00;
17'hd8e7:	data_out=16'h9e4;
17'hd8e8:	data_out=16'ha00;
17'hd8e9:	data_out=16'h8a00;
17'hd8ea:	data_out=16'ha00;
17'hd8eb:	data_out=16'ha00;
17'hd8ec:	data_out=16'h89f7;
17'hd8ed:	data_out=16'h9db;
17'hd8ee:	data_out=16'ha00;
17'hd8ef:	data_out=16'h9d9;
17'hd8f0:	data_out=16'ha00;
17'hd8f1:	data_out=16'h8a00;
17'hd8f2:	data_out=16'ha00;
17'hd8f3:	data_out=16'ha00;
17'hd8f4:	data_out=16'h72f;
17'hd8f5:	data_out=16'ha00;
17'hd8f6:	data_out=16'h89fe;
17'hd8f7:	data_out=16'h8a00;
17'hd8f8:	data_out=16'ha00;
17'hd8f9:	data_out=16'h8a00;
17'hd8fa:	data_out=16'h9c9;
17'hd8fb:	data_out=16'ha00;
17'hd8fc:	data_out=16'h8a00;
17'hd8fd:	data_out=16'ha00;
17'hd8fe:	data_out=16'ha00;
17'hd8ff:	data_out=16'ha00;
17'hd900:	data_out=16'h8a00;
17'hd901:	data_out=16'h8a00;
17'hd902:	data_out=16'h8a00;
17'hd903:	data_out=16'h9be;
17'hd904:	data_out=16'h89a4;
17'hd905:	data_out=16'ha00;
17'hd906:	data_out=16'ha00;
17'hd907:	data_out=16'h8a00;
17'hd908:	data_out=16'h8a00;
17'hd909:	data_out=16'h8a00;
17'hd90a:	data_out=16'h8a00;
17'hd90b:	data_out=16'h8a00;
17'hd90c:	data_out=16'h8a00;
17'hd90d:	data_out=16'h89fd;
17'hd90e:	data_out=16'ha00;
17'hd90f:	data_out=16'h8a00;
17'hd910:	data_out=16'h89b6;
17'hd911:	data_out=16'h82a2;
17'hd912:	data_out=16'h87f6;
17'hd913:	data_out=16'h9ec;
17'hd914:	data_out=16'h9ff;
17'hd915:	data_out=16'h87b6;
17'hd916:	data_out=16'h8501;
17'hd917:	data_out=16'h9d8;
17'hd918:	data_out=16'h8a00;
17'hd919:	data_out=16'h8a00;
17'hd91a:	data_out=16'ha00;
17'hd91b:	data_out=16'h89fc;
17'hd91c:	data_out=16'h9eb;
17'hd91d:	data_out=16'h8a00;
17'hd91e:	data_out=16'h9e9;
17'hd91f:	data_out=16'h9fe;
17'hd920:	data_out=16'h9f6;
17'hd921:	data_out=16'ha00;
17'hd922:	data_out=16'h9fc;
17'hd923:	data_out=16'h8a00;
17'hd924:	data_out=16'h8a00;
17'hd925:	data_out=16'h8320;
17'hd926:	data_out=16'h8a00;
17'hd927:	data_out=16'h8a00;
17'hd928:	data_out=16'ha00;
17'hd929:	data_out=16'h8b1;
17'hd92a:	data_out=16'h89ff;
17'hd92b:	data_out=16'h8a00;
17'hd92c:	data_out=16'h1ae;
17'hd92d:	data_out=16'h8a00;
17'hd92e:	data_out=16'h9b0;
17'hd92f:	data_out=16'h9c8;
17'hd930:	data_out=16'h8a00;
17'hd931:	data_out=16'h8a00;
17'hd932:	data_out=16'h9b2;
17'hd933:	data_out=16'ha00;
17'hd934:	data_out=16'h8a00;
17'hd935:	data_out=16'h8a00;
17'hd936:	data_out=16'h8a00;
17'hd937:	data_out=16'h89ff;
17'hd938:	data_out=16'ha00;
17'hd939:	data_out=16'ha00;
17'hd93a:	data_out=16'h8a00;
17'hd93b:	data_out=16'h8a00;
17'hd93c:	data_out=16'h9bf;
17'hd93d:	data_out=16'h9d3;
17'hd93e:	data_out=16'ha00;
17'hd93f:	data_out=16'ha00;
17'hd940:	data_out=16'h9cd;
17'hd941:	data_out=16'h8a00;
17'hd942:	data_out=16'h8a00;
17'hd943:	data_out=16'ha00;
17'hd944:	data_out=16'h8a00;
17'hd945:	data_out=16'h876c;
17'hd946:	data_out=16'h8a00;
17'hd947:	data_out=16'h8a00;
17'hd948:	data_out=16'h94e;
17'hd949:	data_out=16'h89f5;
17'hd94a:	data_out=16'h8a00;
17'hd94b:	data_out=16'h8a00;
17'hd94c:	data_out=16'h87f4;
17'hd94d:	data_out=16'ha00;
17'hd94e:	data_out=16'h89f9;
17'hd94f:	data_out=16'h8a00;
17'hd950:	data_out=16'ha00;
17'hd951:	data_out=16'h9cf;
17'hd952:	data_out=16'h8a00;
17'hd953:	data_out=16'h89e5;
17'hd954:	data_out=16'h98b;
17'hd955:	data_out=16'h88e;
17'hd956:	data_out=16'h8a00;
17'hd957:	data_out=16'h8e6;
17'hd958:	data_out=16'h8427;
17'hd959:	data_out=16'h9e8;
17'hd95a:	data_out=16'h8101;
17'hd95b:	data_out=16'h89ee;
17'hd95c:	data_out=16'ha00;
17'hd95d:	data_out=16'h58d;
17'hd95e:	data_out=16'ha00;
17'hd95f:	data_out=16'h88c7;
17'hd960:	data_out=16'h8a00;
17'hd961:	data_out=16'h9f2;
17'hd962:	data_out=16'h2f0;
17'hd963:	data_out=16'ha00;
17'hd964:	data_out=16'h8a00;
17'hd965:	data_out=16'h8a00;
17'hd966:	data_out=16'h8a00;
17'hd967:	data_out=16'h9f2;
17'hd968:	data_out=16'ha00;
17'hd969:	data_out=16'h8a00;
17'hd96a:	data_out=16'ha00;
17'hd96b:	data_out=16'ha00;
17'hd96c:	data_out=16'h89fc;
17'hd96d:	data_out=16'ha00;
17'hd96e:	data_out=16'ha00;
17'hd96f:	data_out=16'h9da;
17'hd970:	data_out=16'ha00;
17'hd971:	data_out=16'h8a00;
17'hd972:	data_out=16'ha00;
17'hd973:	data_out=16'ha00;
17'hd974:	data_out=16'h8a00;
17'hd975:	data_out=16'ha00;
17'hd976:	data_out=16'h8a00;
17'hd977:	data_out=16'h8a00;
17'hd978:	data_out=16'ha00;
17'hd979:	data_out=16'h89e6;
17'hd97a:	data_out=16'h9fc;
17'hd97b:	data_out=16'ha00;
17'hd97c:	data_out=16'h8a00;
17'hd97d:	data_out=16'ha00;
17'hd97e:	data_out=16'h9fa;
17'hd97f:	data_out=16'ha00;
17'hd980:	data_out=16'h8a00;
17'hd981:	data_out=16'h8a00;
17'hd982:	data_out=16'h8a00;
17'hd983:	data_out=16'h9a1;
17'hd984:	data_out=16'h8a00;
17'hd985:	data_out=16'h9bd;
17'hd986:	data_out=16'ha00;
17'hd987:	data_out=16'h8a00;
17'hd988:	data_out=16'h8a00;
17'hd989:	data_out=16'h5cb;
17'hd98a:	data_out=16'h8a00;
17'hd98b:	data_out=16'h8a00;
17'hd98c:	data_out=16'h8a00;
17'hd98d:	data_out=16'h8937;
17'hd98e:	data_out=16'ha00;
17'hd98f:	data_out=16'h885d;
17'hd990:	data_out=16'h8f3;
17'hd991:	data_out=16'h8a00;
17'hd992:	data_out=16'h999;
17'hd993:	data_out=16'h9f3;
17'hd994:	data_out=16'h9da;
17'hd995:	data_out=16'h8a00;
17'hd996:	data_out=16'h8a00;
17'hd997:	data_out=16'h9c1;
17'hd998:	data_out=16'h89ff;
17'hd999:	data_out=16'h8a00;
17'hd99a:	data_out=16'h9d7;
17'hd99b:	data_out=16'h89fe;
17'hd99c:	data_out=16'h9a8;
17'hd99d:	data_out=16'h8a00;
17'hd99e:	data_out=16'h9d1;
17'hd99f:	data_out=16'h9e3;
17'hd9a0:	data_out=16'h8286;
17'hd9a1:	data_out=16'ha00;
17'hd9a2:	data_out=16'h9f6;
17'hd9a3:	data_out=16'h8a00;
17'hd9a4:	data_out=16'h8a00;
17'hd9a5:	data_out=16'h808e;
17'hd9a6:	data_out=16'h8a00;
17'hd9a7:	data_out=16'h8a00;
17'hd9a8:	data_out=16'ha00;
17'hd9a9:	data_out=16'h8298;
17'hd9aa:	data_out=16'h89ff;
17'hd9ab:	data_out=16'h8a00;
17'hd9ac:	data_out=16'h89ff;
17'hd9ad:	data_out=16'h8a00;
17'hd9ae:	data_out=16'h9c2;
17'hd9af:	data_out=16'h9d1;
17'hd9b0:	data_out=16'h8a00;
17'hd9b1:	data_out=16'h8a00;
17'hd9b2:	data_out=16'h8a00;
17'hd9b3:	data_out=16'ha00;
17'hd9b4:	data_out=16'h8a00;
17'hd9b5:	data_out=16'h8a00;
17'hd9b6:	data_out=16'h8a00;
17'hd9b7:	data_out=16'h89ff;
17'hd9b8:	data_out=16'ha00;
17'hd9b9:	data_out=16'ha00;
17'hd9ba:	data_out=16'h8a00;
17'hd9bb:	data_out=16'h8a00;
17'hd9bc:	data_out=16'h8406;
17'hd9bd:	data_out=16'h380;
17'hd9be:	data_out=16'ha00;
17'hd9bf:	data_out=16'h9bd;
17'hd9c0:	data_out=16'h850c;
17'hd9c1:	data_out=16'h8a00;
17'hd9c2:	data_out=16'h8a00;
17'hd9c3:	data_out=16'ha00;
17'hd9c4:	data_out=16'h8a00;
17'hd9c5:	data_out=16'h8a00;
17'hd9c6:	data_out=16'h8a00;
17'hd9c7:	data_out=16'h8a00;
17'hd9c8:	data_out=16'h9f0;
17'hd9c9:	data_out=16'h89fc;
17'hd9ca:	data_out=16'h8a00;
17'hd9cb:	data_out=16'h8a00;
17'hd9cc:	data_out=16'h8994;
17'hd9cd:	data_out=16'ha00;
17'hd9ce:	data_out=16'h3da;
17'hd9cf:	data_out=16'h8a00;
17'hd9d0:	data_out=16'h9fc;
17'hd9d1:	data_out=16'h9ab;
17'hd9d2:	data_out=16'h8a00;
17'hd9d3:	data_out=16'h8a00;
17'hd9d4:	data_out=16'h853a;
17'hd9d5:	data_out=16'h94a;
17'hd9d6:	data_out=16'h8a00;
17'hd9d7:	data_out=16'h7db;
17'hd9d8:	data_out=16'h85e8;
17'hd9d9:	data_out=16'h9c3;
17'hd9da:	data_out=16'h9bc;
17'hd9db:	data_out=16'h8a00;
17'hd9dc:	data_out=16'h9ac;
17'hd9dd:	data_out=16'h8191;
17'hd9de:	data_out=16'ha00;
17'hd9df:	data_out=16'h8456;
17'hd9e0:	data_out=16'h8a00;
17'hd9e1:	data_out=16'h89ff;
17'hd9e2:	data_out=16'h72;
17'hd9e3:	data_out=16'ha00;
17'hd9e4:	data_out=16'h8a00;
17'hd9e5:	data_out=16'h8a00;
17'hd9e6:	data_out=16'h8a00;
17'hd9e7:	data_out=16'h9cf;
17'hd9e8:	data_out=16'ha00;
17'hd9e9:	data_out=16'h8a00;
17'hd9ea:	data_out=16'ha00;
17'hd9eb:	data_out=16'h9eb;
17'hd9ec:	data_out=16'h8a00;
17'hd9ed:	data_out=16'ha00;
17'hd9ee:	data_out=16'ha00;
17'hd9ef:	data_out=16'h96c;
17'hd9f0:	data_out=16'ha00;
17'hd9f1:	data_out=16'h8a00;
17'hd9f2:	data_out=16'h9e1;
17'hd9f3:	data_out=16'h9a4;
17'hd9f4:	data_out=16'h8a00;
17'hd9f5:	data_out=16'h80a5;
17'hd9f6:	data_out=16'h8a00;
17'hd9f7:	data_out=16'h89d5;
17'hd9f8:	data_out=16'ha00;
17'hd9f9:	data_out=16'h89b9;
17'hd9fa:	data_out=16'h9ee;
17'hd9fb:	data_out=16'ha00;
17'hd9fc:	data_out=16'h89fe;
17'hd9fd:	data_out=16'ha00;
17'hd9fe:	data_out=16'h9fa;
17'hd9ff:	data_out=16'ha00;
17'hda00:	data_out=16'h8a00;
17'hda01:	data_out=16'h8a00;
17'hda02:	data_out=16'h84ae;
17'hda03:	data_out=16'h9ed;
17'hda04:	data_out=16'h8a00;
17'hda05:	data_out=16'h8a00;
17'hda06:	data_out=16'ha00;
17'hda07:	data_out=16'h8a00;
17'hda08:	data_out=16'h8a00;
17'hda09:	data_out=16'h978;
17'hda0a:	data_out=16'h8a00;
17'hda0b:	data_out=16'h8295;
17'hda0c:	data_out=16'h8a00;
17'hda0d:	data_out=16'h8662;
17'hda0e:	data_out=16'h9fe;
17'hda0f:	data_out=16'h9ae;
17'hda10:	data_out=16'h9df;
17'hda11:	data_out=16'h89eb;
17'hda12:	data_out=16'h9e0;
17'hda13:	data_out=16'ha00;
17'hda14:	data_out=16'h9ed;
17'hda15:	data_out=16'h8a00;
17'hda16:	data_out=16'h8a00;
17'hda17:	data_out=16'h9ea;
17'hda18:	data_out=16'h84ae;
17'hda19:	data_out=16'h8a00;
17'hda1a:	data_out=16'h8a00;
17'hda1b:	data_out=16'h83ed;
17'hda1c:	data_out=16'h9d5;
17'hda1d:	data_out=16'h8a00;
17'hda1e:	data_out=16'h9f5;
17'hda1f:	data_out=16'h9af;
17'hda20:	data_out=16'h89d8;
17'hda21:	data_out=16'ha00;
17'hda22:	data_out=16'h9ec;
17'hda23:	data_out=16'h8a00;
17'hda24:	data_out=16'h8a00;
17'hda25:	data_out=16'h986;
17'hda26:	data_out=16'h8a00;
17'hda27:	data_out=16'h8a00;
17'hda28:	data_out=16'ha00;
17'hda29:	data_out=16'h89ce;
17'hda2a:	data_out=16'h89fe;
17'hda2b:	data_out=16'h8a00;
17'hda2c:	data_out=16'h8a00;
17'hda2d:	data_out=16'h89fe;
17'hda2e:	data_out=16'h9a9;
17'hda2f:	data_out=16'h8895;
17'hda30:	data_out=16'h8a00;
17'hda31:	data_out=16'h8a00;
17'hda32:	data_out=16'h8a00;
17'hda33:	data_out=16'ha00;
17'hda34:	data_out=16'h8a00;
17'hda35:	data_out=16'h8a00;
17'hda36:	data_out=16'h8a00;
17'hda37:	data_out=16'h30a;
17'hda38:	data_out=16'ha00;
17'hda39:	data_out=16'ha00;
17'hda3a:	data_out=16'h6b7;
17'hda3b:	data_out=16'h8a00;
17'hda3c:	data_out=16'h89f8;
17'hda3d:	data_out=16'h89a6;
17'hda3e:	data_out=16'ha00;
17'hda3f:	data_out=16'h8a00;
17'hda40:	data_out=16'h8a00;
17'hda41:	data_out=16'h8a00;
17'hda42:	data_out=16'h8a00;
17'hda43:	data_out=16'h9fc;
17'hda44:	data_out=16'h8a00;
17'hda45:	data_out=16'h8a00;
17'hda46:	data_out=16'h8a00;
17'hda47:	data_out=16'h2ee;
17'hda48:	data_out=16'h9d9;
17'hda49:	data_out=16'h85e3;
17'hda4a:	data_out=16'h8a00;
17'hda4b:	data_out=16'h8a00;
17'hda4c:	data_out=16'h95e;
17'hda4d:	data_out=16'h9fd;
17'hda4e:	data_out=16'h9e2;
17'hda4f:	data_out=16'h89f0;
17'hda50:	data_out=16'h80b;
17'hda51:	data_out=16'h9d6;
17'hda52:	data_out=16'h8a00;
17'hda53:	data_out=16'h8a00;
17'hda54:	data_out=16'h89cb;
17'hda55:	data_out=16'h9aa;
17'hda56:	data_out=16'h8a00;
17'hda57:	data_out=16'h980;
17'hda58:	data_out=16'h84b3;
17'hda59:	data_out=16'h899c;
17'hda5a:	data_out=16'h9d6;
17'hda5b:	data_out=16'h8a00;
17'hda5c:	data_out=16'h89d5;
17'hda5d:	data_out=16'h88ac;
17'hda5e:	data_out=16'h84fe;
17'hda5f:	data_out=16'h49e;
17'hda60:	data_out=16'h8a00;
17'hda61:	data_out=16'h8a00;
17'hda62:	data_out=16'h9a2;
17'hda63:	data_out=16'h9ff;
17'hda64:	data_out=16'h8a00;
17'hda65:	data_out=16'h8a00;
17'hda66:	data_out=16'h8a00;
17'hda67:	data_out=16'h79f;
17'hda68:	data_out=16'ha00;
17'hda69:	data_out=16'h8a00;
17'hda6a:	data_out=16'h9fd;
17'hda6b:	data_out=16'h88f6;
17'hda6c:	data_out=16'h89ff;
17'hda6d:	data_out=16'ha00;
17'hda6e:	data_out=16'h9fd;
17'hda6f:	data_out=16'h8a00;
17'hda70:	data_out=16'h9fe;
17'hda71:	data_out=16'h5c7;
17'hda72:	data_out=16'h265;
17'hda73:	data_out=16'h8945;
17'hda74:	data_out=16'h8a00;
17'hda75:	data_out=16'h8a00;
17'hda76:	data_out=16'h8a00;
17'hda77:	data_out=16'h9b1;
17'hda78:	data_out=16'h8ab;
17'hda79:	data_out=16'h81a7;
17'hda7a:	data_out=16'h9fd;
17'hda7b:	data_out=16'ha00;
17'hda7c:	data_out=16'h8a00;
17'hda7d:	data_out=16'h9fb;
17'hda7e:	data_out=16'ha00;
17'hda7f:	data_out=16'ha00;
17'hda80:	data_out=16'h89d6;
17'hda81:	data_out=16'h89fb;
17'hda82:	data_out=16'ha00;
17'hda83:	data_out=16'h303;
17'hda84:	data_out=16'h89ff;
17'hda85:	data_out=16'h8a00;
17'hda86:	data_out=16'ha00;
17'hda87:	data_out=16'h1b7;
17'hda88:	data_out=16'h9ee;
17'hda89:	data_out=16'h9fb;
17'hda8a:	data_out=16'h89b7;
17'hda8b:	data_out=16'ha00;
17'hda8c:	data_out=16'h8845;
17'hda8d:	data_out=16'h89c7;
17'hda8e:	data_out=16'ha00;
17'hda8f:	data_out=16'ha00;
17'hda90:	data_out=16'ha00;
17'hda91:	data_out=16'h841c;
17'hda92:	data_out=16'ha00;
17'hda93:	data_out=16'h9ff;
17'hda94:	data_out=16'ha00;
17'hda95:	data_out=16'h89f9;
17'hda96:	data_out=16'h89e8;
17'hda97:	data_out=16'h9f6;
17'hda98:	data_out=16'h9f8;
17'hda99:	data_out=16'h9fe;
17'hda9a:	data_out=16'h8a00;
17'hda9b:	data_out=16'ha00;
17'hda9c:	data_out=16'h8898;
17'hda9d:	data_out=16'h89e7;
17'hda9e:	data_out=16'ha00;
17'hda9f:	data_out=16'h9c4;
17'hdaa0:	data_out=16'h89ae;
17'hdaa1:	data_out=16'ha00;
17'hdaa2:	data_out=16'ha00;
17'hdaa3:	data_out=16'h89d7;
17'hdaa4:	data_out=16'h89da;
17'hdaa5:	data_out=16'ha00;
17'hdaa6:	data_out=16'ha00;
17'hdaa7:	data_out=16'h89de;
17'hdaa8:	data_out=16'ha00;
17'hdaa9:	data_out=16'h8733;
17'hdaaa:	data_out=16'ha00;
17'hdaab:	data_out=16'h9e2;
17'hdaac:	data_out=16'h89fa;
17'hdaad:	data_out=16'h9e5;
17'hdaae:	data_out=16'h9e9;
17'hdaaf:	data_out=16'h8887;
17'hdab0:	data_out=16'h8844;
17'hdab1:	data_out=16'h8a00;
17'hdab2:	data_out=16'h8a00;
17'hdab3:	data_out=16'ha00;
17'hdab4:	data_out=16'h8a00;
17'hdab5:	data_out=16'h89d1;
17'hdab6:	data_out=16'h9fd;
17'hdab7:	data_out=16'ha00;
17'hdab8:	data_out=16'h869d;
17'hdab9:	data_out=16'ha00;
17'hdaba:	data_out=16'h9fc;
17'hdabb:	data_out=16'h8a00;
17'hdabc:	data_out=16'h894c;
17'hdabd:	data_out=16'h88fe;
17'hdabe:	data_out=16'ha00;
17'hdabf:	data_out=16'h8a00;
17'hdac0:	data_out=16'h89fc;
17'hdac1:	data_out=16'h8675;
17'hdac2:	data_out=16'h54c;
17'hdac3:	data_out=16'h859;
17'hdac4:	data_out=16'h89fe;
17'hdac5:	data_out=16'h89fa;
17'hdac6:	data_out=16'h9f7;
17'hdac7:	data_out=16'ha00;
17'hdac8:	data_out=16'h9e9;
17'hdac9:	data_out=16'ha00;
17'hdaca:	data_out=16'h89d5;
17'hdacb:	data_out=16'hbe;
17'hdacc:	data_out=16'h9fd;
17'hdacd:	data_out=16'ha00;
17'hdace:	data_out=16'h9fe;
17'hdacf:	data_out=16'ha00;
17'hdad0:	data_out=16'h89aa;
17'hdad1:	data_out=16'h8558;
17'hdad2:	data_out=16'h89d9;
17'hdad3:	data_out=16'h431;
17'hdad4:	data_out=16'h8692;
17'hdad5:	data_out=16'h9fe;
17'hdad6:	data_out=16'h9f6;
17'hdad7:	data_out=16'h9fb;
17'hdad8:	data_out=16'h8038;
17'hdad9:	data_out=16'h8978;
17'hdada:	data_out=16'h9f9;
17'hdadb:	data_out=16'h89fb;
17'hdadc:	data_out=16'h89ff;
17'hdadd:	data_out=16'h88eb;
17'hdade:	data_out=16'h8672;
17'hdadf:	data_out=16'h9ff;
17'hdae0:	data_out=16'h9f8;
17'hdae1:	data_out=16'h8a00;
17'hdae2:	data_out=16'h9ff;
17'hdae3:	data_out=16'ha00;
17'hdae4:	data_out=16'h89ff;
17'hdae5:	data_out=16'h89ea;
17'hdae6:	data_out=16'h9e0;
17'hdae7:	data_out=16'h9c0;
17'hdae8:	data_out=16'ha00;
17'hdae9:	data_out=16'ha00;
17'hdaea:	data_out=16'ha00;
17'hdaeb:	data_out=16'h89c2;
17'hdaec:	data_out=16'h897e;
17'hdaed:	data_out=16'ha00;
17'hdaee:	data_out=16'ha00;
17'hdaef:	data_out=16'h8a00;
17'hdaf0:	data_out=16'ha00;
17'hdaf1:	data_out=16'h9f6;
17'hdaf2:	data_out=16'h8971;
17'hdaf3:	data_out=16'h89b6;
17'hdaf4:	data_out=16'h89c2;
17'hdaf5:	data_out=16'h8a00;
17'hdaf6:	data_out=16'h9e6;
17'hdaf7:	data_out=16'ha00;
17'hdaf8:	data_out=16'h8a00;
17'hdaf9:	data_out=16'ha00;
17'hdafa:	data_out=16'ha00;
17'hdafb:	data_out=16'ha00;
17'hdafc:	data_out=16'h9ec;
17'hdafd:	data_out=16'ha3;
17'hdafe:	data_out=16'ha00;
17'hdaff:	data_out=16'h8a00;
17'hdb00:	data_out=16'h89d0;
17'hdb01:	data_out=16'h89fa;
17'hdb02:	data_out=16'ha00;
17'hdb03:	data_out=16'h8988;
17'hdb04:	data_out=16'h89fb;
17'hdb05:	data_out=16'h8a00;
17'hdb06:	data_out=16'h8148;
17'hdb07:	data_out=16'ha00;
17'hdb08:	data_out=16'ha00;
17'hdb09:	data_out=16'ha00;
17'hdb0a:	data_out=16'h8993;
17'hdb0b:	data_out=16'ha00;
17'hdb0c:	data_out=16'h9e1;
17'hdb0d:	data_out=16'h89f5;
17'hdb0e:	data_out=16'ha00;
17'hdb0f:	data_out=16'ha00;
17'hdb10:	data_out=16'h955;
17'hdb11:	data_out=16'h86fe;
17'hdb12:	data_out=16'h9fb;
17'hdb13:	data_out=16'h8901;
17'hdb14:	data_out=16'h9f2;
17'hdb15:	data_out=16'h8a00;
17'hdb16:	data_out=16'h89fd;
17'hdb17:	data_out=16'h51e;
17'hdb18:	data_out=16'h9fe;
17'hdb19:	data_out=16'ha00;
17'hdb1a:	data_out=16'h8a00;
17'hdb1b:	data_out=16'ha00;
17'hdb1c:	data_out=16'h89f2;
17'hdb1d:	data_out=16'h89be;
17'hdb1e:	data_out=16'h9ff;
17'hdb1f:	data_out=16'h993;
17'hdb20:	data_out=16'h89ca;
17'hdb21:	data_out=16'ha00;
17'hdb22:	data_out=16'h9b1;
17'hdb23:	data_out=16'ha00;
17'hdb24:	data_out=16'ha00;
17'hdb25:	data_out=16'h9f4;
17'hdb26:	data_out=16'ha00;
17'hdb27:	data_out=16'h77;
17'hdb28:	data_out=16'ha00;
17'hdb29:	data_out=16'h87db;
17'hdb2a:	data_out=16'ha00;
17'hdb2b:	data_out=16'ha00;
17'hdb2c:	data_out=16'h8a00;
17'hdb2d:	data_out=16'h84b5;
17'hdb2e:	data_out=16'h9f0;
17'hdb2f:	data_out=16'h8953;
17'hdb30:	data_out=16'h83e1;
17'hdb31:	data_out=16'h89fd;
17'hdb32:	data_out=16'h89f3;
17'hdb33:	data_out=16'h9fb;
17'hdb34:	data_out=16'h89ee;
17'hdb35:	data_out=16'h8934;
17'hdb36:	data_out=16'ha00;
17'hdb37:	data_out=16'ha00;
17'hdb38:	data_out=16'h8a00;
17'hdb39:	data_out=16'h9fb;
17'hdb3a:	data_out=16'ha00;
17'hdb3b:	data_out=16'h89a0;
17'hdb3c:	data_out=16'h88ea;
17'hdb3d:	data_out=16'h8972;
17'hdb3e:	data_out=16'ha00;
17'hdb3f:	data_out=16'h8a00;
17'hdb40:	data_out=16'h89ff;
17'hdb41:	data_out=16'h7e2;
17'hdb42:	data_out=16'h8a8;
17'hdb43:	data_out=16'h89c8;
17'hdb44:	data_out=16'h89f3;
17'hdb45:	data_out=16'h8a00;
17'hdb46:	data_out=16'h9fb;
17'hdb47:	data_out=16'ha00;
17'hdb48:	data_out=16'h989;
17'hdb49:	data_out=16'h6bd;
17'hdb4a:	data_out=16'h9d7;
17'hdb4b:	data_out=16'h99d;
17'hdb4c:	data_out=16'h9f2;
17'hdb4d:	data_out=16'h9eb;
17'hdb4e:	data_out=16'ha00;
17'hdb4f:	data_out=16'ha00;
17'hdb50:	data_out=16'h89ff;
17'hdb51:	data_out=16'h89a8;
17'hdb52:	data_out=16'h268;
17'hdb53:	data_out=16'h9ae;
17'hdb54:	data_out=16'h36;
17'hdb55:	data_out=16'h9f6;
17'hdb56:	data_out=16'h9f4;
17'hdb57:	data_out=16'h2ff;
17'hdb58:	data_out=16'hec;
17'hdb59:	data_out=16'h89c8;
17'hdb5a:	data_out=16'h9ee;
17'hdb5b:	data_out=16'h89c4;
17'hdb5c:	data_out=16'h8a00;
17'hdb5d:	data_out=16'h89b0;
17'hdb5e:	data_out=16'h89b7;
17'hdb5f:	data_out=16'ha00;
17'hdb60:	data_out=16'h632;
17'hdb61:	data_out=16'h8a00;
17'hdb62:	data_out=16'h9f4;
17'hdb63:	data_out=16'h9f9;
17'hdb64:	data_out=16'h89ff;
17'hdb65:	data_out=16'h899e;
17'hdb66:	data_out=16'ha00;
17'hdb67:	data_out=16'h9ff;
17'hdb68:	data_out=16'ha00;
17'hdb69:	data_out=16'ha00;
17'hdb6a:	data_out=16'ha00;
17'hdb6b:	data_out=16'h89fd;
17'hdb6c:	data_out=16'h899f;
17'hdb6d:	data_out=16'h9fc;
17'hdb6e:	data_out=16'ha00;
17'hdb6f:	data_out=16'h89ff;
17'hdb70:	data_out=16'ha00;
17'hdb71:	data_out=16'ha00;
17'hdb72:	data_out=16'h8a00;
17'hdb73:	data_out=16'h8a00;
17'hdb74:	data_out=16'h845e;
17'hdb75:	data_out=16'h8a00;
17'hdb76:	data_out=16'ha00;
17'hdb77:	data_out=16'h9f6;
17'hdb78:	data_out=16'h8a00;
17'hdb79:	data_out=16'ha00;
17'hdb7a:	data_out=16'h9fb;
17'hdb7b:	data_out=16'ha00;
17'hdb7c:	data_out=16'h9f9;
17'hdb7d:	data_out=16'h891d;
17'hdb7e:	data_out=16'h83c7;
17'hdb7f:	data_out=16'h8a00;
17'hdb80:	data_out=16'h8a00;
17'hdb81:	data_out=16'h8a00;
17'hdb82:	data_out=16'h9c8;
17'hdb83:	data_out=16'h89fc;
17'hdb84:	data_out=16'h89ff;
17'hdb85:	data_out=16'h8a00;
17'hdb86:	data_out=16'h892a;
17'hdb87:	data_out=16'ha00;
17'hdb88:	data_out=16'h9d0;
17'hdb89:	data_out=16'h9f1;
17'hdb8a:	data_out=16'h8a00;
17'hdb8b:	data_out=16'ha00;
17'hdb8c:	data_out=16'ha00;
17'hdb8d:	data_out=16'h89fd;
17'hdb8e:	data_out=16'h89b0;
17'hdb8f:	data_out=16'h9f4;
17'hdb90:	data_out=16'h7fe;
17'hdb91:	data_out=16'h89ed;
17'hdb92:	data_out=16'h99f;
17'hdb93:	data_out=16'h89f9;
17'hdb94:	data_out=16'h889e;
17'hdb95:	data_out=16'h8a00;
17'hdb96:	data_out=16'h8a00;
17'hdb97:	data_out=16'h8928;
17'hdb98:	data_out=16'h9df;
17'hdb99:	data_out=16'ha00;
17'hdb9a:	data_out=16'h8a00;
17'hdb9b:	data_out=16'h9e9;
17'hdb9c:	data_out=16'h8a00;
17'hdb9d:	data_out=16'h89e8;
17'hdb9e:	data_out=16'h8962;
17'hdb9f:	data_out=16'h89de;
17'hdba0:	data_out=16'h89fa;
17'hdba1:	data_out=16'h89ab;
17'hdba2:	data_out=16'h8922;
17'hdba3:	data_out=16'ha00;
17'hdba4:	data_out=16'ha00;
17'hdba5:	data_out=16'h89b4;
17'hdba6:	data_out=16'h828f;
17'hdba7:	data_out=16'h145;
17'hdba8:	data_out=16'h86f9;
17'hdba9:	data_out=16'h8871;
17'hdbaa:	data_out=16'ha00;
17'hdbab:	data_out=16'ha00;
17'hdbac:	data_out=16'h8a00;
17'hdbad:	data_out=16'h8986;
17'hdbae:	data_out=16'h9a3;
17'hdbaf:	data_out=16'h8818;
17'hdbb0:	data_out=16'h87e0;
17'hdbb1:	data_out=16'h89ff;
17'hdbb2:	data_out=16'h89fd;
17'hdbb3:	data_out=16'h726;
17'hdbb4:	data_out=16'h89fb;
17'hdbb5:	data_out=16'h89f8;
17'hdbb6:	data_out=16'h9fc;
17'hdbb7:	data_out=16'h9dc;
17'hdbb8:	data_out=16'h8a00;
17'hdbb9:	data_out=16'h37;
17'hdbba:	data_out=16'h9f8;
17'hdbbb:	data_out=16'h85ee;
17'hdbbc:	data_out=16'h8982;
17'hdbbd:	data_out=16'h89fb;
17'hdbbe:	data_out=16'h86f1;
17'hdbbf:	data_out=16'h8a00;
17'hdbc0:	data_out=16'h89fd;
17'hdbc1:	data_out=16'h995;
17'hdbc2:	data_out=16'h82cf;
17'hdbc3:	data_out=16'h8854;
17'hdbc4:	data_out=16'h89ec;
17'hdbc5:	data_out=16'h8a00;
17'hdbc6:	data_out=16'h881a;
17'hdbc7:	data_out=16'ha00;
17'hdbc8:	data_out=16'h816;
17'hdbc9:	data_out=16'h89ac;
17'hdbca:	data_out=16'ha00;
17'hdbcb:	data_out=16'h974;
17'hdbcc:	data_out=16'h81e8;
17'hdbcd:	data_out=16'h86bb;
17'hdbce:	data_out=16'ha00;
17'hdbcf:	data_out=16'h9f4;
17'hdbd0:	data_out=16'h89fc;
17'hdbd1:	data_out=16'h89f7;
17'hdbd2:	data_out=16'h82e2;
17'hdbd3:	data_out=16'h980;
17'hdbd4:	data_out=16'h81b4;
17'hdbd5:	data_out=16'h86f0;
17'hdbd6:	data_out=16'h8929;
17'hdbd7:	data_out=16'h89a9;
17'hdbd8:	data_out=16'h8876;
17'hdbd9:	data_out=16'h89f7;
17'hdbda:	data_out=16'h9b2;
17'hdbdb:	data_out=16'h89f2;
17'hdbdc:	data_out=16'h8a00;
17'hdbdd:	data_out=16'h89fd;
17'hdbde:	data_out=16'h891e;
17'hdbdf:	data_out=16'h9dd;
17'hdbe0:	data_out=16'h8967;
17'hdbe1:	data_out=16'h8a00;
17'hdbe2:	data_out=16'h754;
17'hdbe3:	data_out=16'h987;
17'hdbe4:	data_out=16'h89ec;
17'hdbe5:	data_out=16'h88df;
17'hdbe6:	data_out=16'ha00;
17'hdbe7:	data_out=16'ha00;
17'hdbe8:	data_out=16'h88ac;
17'hdbe9:	data_out=16'h9d2;
17'hdbea:	data_out=16'h89b2;
17'hdbeb:	data_out=16'h89ff;
17'hdbec:	data_out=16'h8a00;
17'hdbed:	data_out=16'h8dc;
17'hdbee:	data_out=16'h89b2;
17'hdbef:	data_out=16'h89fe;
17'hdbf0:	data_out=16'h89b0;
17'hdbf1:	data_out=16'h9cd;
17'hdbf2:	data_out=16'h8a00;
17'hdbf3:	data_out=16'h8a00;
17'hdbf4:	data_out=16'h87d1;
17'hdbf5:	data_out=16'h8a00;
17'hdbf6:	data_out=16'ha00;
17'hdbf7:	data_out=16'h9cf;
17'hdbf8:	data_out=16'h8a00;
17'hdbf9:	data_out=16'h9cb;
17'hdbfa:	data_out=16'h5e0;
17'hdbfb:	data_out=16'h86eb;
17'hdbfc:	data_out=16'h9de;
17'hdbfd:	data_out=16'h89d4;
17'hdbfe:	data_out=16'h8a00;
17'hdbff:	data_out=16'h8a00;
17'hdc00:	data_out=16'h89fe;
17'hdc01:	data_out=16'h8a00;
17'hdc02:	data_out=16'h87be;
17'hdc03:	data_out=16'h89fb;
17'hdc04:	data_out=16'h89f5;
17'hdc05:	data_out=16'h8a00;
17'hdc06:	data_out=16'h89f2;
17'hdc07:	data_out=16'ha00;
17'hdc08:	data_out=16'h9ce;
17'hdc09:	data_out=16'h9ed;
17'hdc0a:	data_out=16'h8a00;
17'hdc0b:	data_out=16'ha00;
17'hdc0c:	data_out=16'ha00;
17'hdc0d:	data_out=16'h89fb;
17'hdc0e:	data_out=16'h8a00;
17'hdc0f:	data_out=16'h9c0;
17'hdc10:	data_out=16'h4cb;
17'hdc11:	data_out=16'h89f8;
17'hdc12:	data_out=16'h265;
17'hdc13:	data_out=16'h89f6;
17'hdc14:	data_out=16'h89e0;
17'hdc15:	data_out=16'h89ff;
17'hdc16:	data_out=16'h89fd;
17'hdc17:	data_out=16'h89d3;
17'hdc18:	data_out=16'h82d7;
17'hdc19:	data_out=16'ha00;
17'hdc1a:	data_out=16'h8a00;
17'hdc1b:	data_out=16'h7cf;
17'hdc1c:	data_out=16'h8a00;
17'hdc1d:	data_out=16'h89ee;
17'hdc1e:	data_out=16'h89f5;
17'hdc1f:	data_out=16'h89f7;
17'hdc20:	data_out=16'h89f9;
17'hdc21:	data_out=16'h8a00;
17'hdc22:	data_out=16'h89de;
17'hdc23:	data_out=16'ha00;
17'hdc24:	data_out=16'ha00;
17'hdc25:	data_out=16'h89eb;
17'hdc26:	data_out=16'h8615;
17'hdc27:	data_out=16'hc8;
17'hdc28:	data_out=16'h8a00;
17'hdc29:	data_out=16'h89f8;
17'hdc2a:	data_out=16'h9e4;
17'hdc2b:	data_out=16'ha00;
17'hdc2c:	data_out=16'h89fe;
17'hdc2d:	data_out=16'h89ca;
17'hdc2e:	data_out=16'h65e;
17'hdc2f:	data_out=16'h85cc;
17'hdc30:	data_out=16'h899c;
17'hdc31:	data_out=16'h89ff;
17'hdc32:	data_out=16'h87fb;
17'hdc33:	data_out=16'h89f8;
17'hdc34:	data_out=16'h89ef;
17'hdc35:	data_out=16'h89e9;
17'hdc36:	data_out=16'h9e3;
17'hdc37:	data_out=16'h86a6;
17'hdc38:	data_out=16'h8a00;
17'hdc39:	data_out=16'h89f9;
17'hdc3a:	data_out=16'h9ed;
17'hdc3b:	data_out=16'h918;
17'hdc3c:	data_out=16'h89f5;
17'hdc3d:	data_out=16'h89f9;
17'hdc3e:	data_out=16'h8a00;
17'hdc3f:	data_out=16'h8a00;
17'hdc40:	data_out=16'h89f7;
17'hdc41:	data_out=16'h9ba;
17'hdc42:	data_out=16'h9ec;
17'hdc43:	data_out=16'h80a4;
17'hdc44:	data_out=16'h89e1;
17'hdc45:	data_out=16'h89ff;
17'hdc46:	data_out=16'h89ed;
17'hdc47:	data_out=16'h9fb;
17'hdc48:	data_out=16'h6dc;
17'hdc49:	data_out=16'h89d1;
17'hdc4a:	data_out=16'ha00;
17'hdc4b:	data_out=16'h9f5;
17'hdc4c:	data_out=16'h500;
17'hdc4d:	data_out=16'h89e4;
17'hdc4e:	data_out=16'h9ff;
17'hdc4f:	data_out=16'h9e3;
17'hdc50:	data_out=16'h89f7;
17'hdc51:	data_out=16'h89ff;
17'hdc52:	data_out=16'h846f;
17'hdc53:	data_out=16'h9a3;
17'hdc54:	data_out=16'h85cf;
17'hdc55:	data_out=16'h88f8;
17'hdc56:	data_out=16'h89a4;
17'hdc57:	data_out=16'h89f9;
17'hdc58:	data_out=16'h89ff;
17'hdc59:	data_out=16'h89f5;
17'hdc5a:	data_out=16'h88ed;
17'hdc5b:	data_out=16'h89e8;
17'hdc5c:	data_out=16'h8a00;
17'hdc5d:	data_out=16'h877a;
17'hdc5e:	data_out=16'h8564;
17'hdc5f:	data_out=16'h709;
17'hdc60:	data_out=16'h89c5;
17'hdc61:	data_out=16'h8a00;
17'hdc62:	data_out=16'hb0;
17'hdc63:	data_out=16'h89f0;
17'hdc64:	data_out=16'h89e4;
17'hdc65:	data_out=16'h85f6;
17'hdc66:	data_out=16'ha00;
17'hdc67:	data_out=16'ha00;
17'hdc68:	data_out=16'h8a00;
17'hdc69:	data_out=16'h9db;
17'hdc6a:	data_out=16'h8a00;
17'hdc6b:	data_out=16'h89fb;
17'hdc6c:	data_out=16'h89fe;
17'hdc6d:	data_out=16'h89f2;
17'hdc6e:	data_out=16'h8a00;
17'hdc6f:	data_out=16'h89f9;
17'hdc70:	data_out=16'h8a00;
17'hdc71:	data_out=16'h9b6;
17'hdc72:	data_out=16'h8a00;
17'hdc73:	data_out=16'h8a00;
17'hdc74:	data_out=16'h89c7;
17'hdc75:	data_out=16'h8a00;
17'hdc76:	data_out=16'ha00;
17'hdc77:	data_out=16'h9a6;
17'hdc78:	data_out=16'h89ff;
17'hdc79:	data_out=16'h983;
17'hdc7a:	data_out=16'h89e7;
17'hdc7b:	data_out=16'h8a00;
17'hdc7c:	data_out=16'h9a2;
17'hdc7d:	data_out=16'h89f2;
17'hdc7e:	data_out=16'h8a00;
17'hdc7f:	data_out=16'h8a00;
17'hdc80:	data_out=16'h89fc;
17'hdc81:	data_out=16'h8a00;
17'hdc82:	data_out=16'h884d;
17'hdc83:	data_out=16'h8896;
17'hdc84:	data_out=16'h87c1;
17'hdc85:	data_out=16'h8a00;
17'hdc86:	data_out=16'h89e1;
17'hdc87:	data_out=16'ha00;
17'hdc88:	data_out=16'h9ba;
17'hdc89:	data_out=16'ha00;
17'hdc8a:	data_out=16'h8a00;
17'hdc8b:	data_out=16'ha00;
17'hdc8c:	data_out=16'ha00;
17'hdc8d:	data_out=16'h89d6;
17'hdc8e:	data_out=16'h8a00;
17'hdc8f:	data_out=16'h9fc;
17'hdc90:	data_out=16'h695;
17'hdc91:	data_out=16'h8a00;
17'hdc92:	data_out=16'h8198;
17'hdc93:	data_out=16'h8858;
17'hdc94:	data_out=16'h89e7;
17'hdc95:	data_out=16'h89fe;
17'hdc96:	data_out=16'h8885;
17'hdc97:	data_out=16'h87db;
17'hdc98:	data_out=16'h89fe;
17'hdc99:	data_out=16'ha00;
17'hdc9a:	data_out=16'h8a00;
17'hdc9b:	data_out=16'h8356;
17'hdc9c:	data_out=16'h8a00;
17'hdc9d:	data_out=16'h89f3;
17'hdc9e:	data_out=16'h89f5;
17'hdc9f:	data_out=16'h89d8;
17'hdca0:	data_out=16'h89fa;
17'hdca1:	data_out=16'h8a00;
17'hdca2:	data_out=16'h890a;
17'hdca3:	data_out=16'h9fd;
17'hdca4:	data_out=16'h9fd;
17'hdca5:	data_out=16'h89f3;
17'hdca6:	data_out=16'h9e0;
17'hdca7:	data_out=16'h9c8;
17'hdca8:	data_out=16'h8a00;
17'hdca9:	data_out=16'h8a00;
17'hdcaa:	data_out=16'ha00;
17'hdcab:	data_out=16'ha00;
17'hdcac:	data_out=16'h89a4;
17'hdcad:	data_out=16'h84ba;
17'hdcae:	data_out=16'ha00;
17'hdcaf:	data_out=16'h698;
17'hdcb0:	data_out=16'h89dd;
17'hdcb1:	data_out=16'h8a00;
17'hdcb2:	data_out=16'h8540;
17'hdcb3:	data_out=16'h89f8;
17'hdcb4:	data_out=16'h89d7;
17'hdcb5:	data_out=16'h8877;
17'hdcb6:	data_out=16'h9db;
17'hdcb7:	data_out=16'h865b;
17'hdcb8:	data_out=16'h8a00;
17'hdcb9:	data_out=16'h89fd;
17'hdcba:	data_out=16'h9f0;
17'hdcbb:	data_out=16'ha00;
17'hdcbc:	data_out=16'h8a00;
17'hdcbd:	data_out=16'h89f9;
17'hdcbe:	data_out=16'h8a00;
17'hdcbf:	data_out=16'h8a00;
17'hdcc0:	data_out=16'h884c;
17'hdcc1:	data_out=16'h982;
17'hdcc2:	data_out=16'ha00;
17'hdcc3:	data_out=16'h828;
17'hdcc4:	data_out=16'h895c;
17'hdcc5:	data_out=16'h89fe;
17'hdcc6:	data_out=16'h8a00;
17'hdcc7:	data_out=16'ha00;
17'hdcc8:	data_out=16'h9d6;
17'hdcc9:	data_out=16'h89db;
17'hdcca:	data_out=16'ha00;
17'hdccb:	data_out=16'ha00;
17'hdccc:	data_out=16'h9af;
17'hdccd:	data_out=16'h89f2;
17'hdcce:	data_out=16'h9f6;
17'hdccf:	data_out=16'h9ef;
17'hdcd0:	data_out=16'h893c;
17'hdcd1:	data_out=16'h8a00;
17'hdcd2:	data_out=16'h85d7;
17'hdcd3:	data_out=16'h9e1;
17'hdcd4:	data_out=16'h8861;
17'hdcd5:	data_out=16'h8843;
17'hdcd6:	data_out=16'h89ba;
17'hdcd7:	data_out=16'h89fe;
17'hdcd8:	data_out=16'h8a00;
17'hdcd9:	data_out=16'h89f1;
17'hdcda:	data_out=16'h89d7;
17'hdcdb:	data_out=16'h89ec;
17'hdcdc:	data_out=16'h8a00;
17'hdcdd:	data_out=16'h7e2;
17'hdcde:	data_out=16'h9ae;
17'hdcdf:	data_out=16'h86f8;
17'hdce0:	data_out=16'h84a0;
17'hdce1:	data_out=16'h8a00;
17'hdce2:	data_out=16'h9fe;
17'hdce3:	data_out=16'h89ec;
17'hdce4:	data_out=16'h89c4;
17'hdce5:	data_out=16'h689;
17'hdce6:	data_out=16'ha00;
17'hdce7:	data_out=16'ha00;
17'hdce8:	data_out=16'h8a00;
17'hdce9:	data_out=16'h9d2;
17'hdcea:	data_out=16'h8a00;
17'hdceb:	data_out=16'h89fb;
17'hdcec:	data_out=16'h886c;
17'hdced:	data_out=16'h89ee;
17'hdcee:	data_out=16'h8a00;
17'hdcef:	data_out=16'h8101;
17'hdcf0:	data_out=16'h8a00;
17'hdcf1:	data_out=16'h9ff;
17'hdcf2:	data_out=16'h8a00;
17'hdcf3:	data_out=16'h8a00;
17'hdcf4:	data_out=16'h89f0;
17'hdcf5:	data_out=16'h8a00;
17'hdcf6:	data_out=16'ha00;
17'hdcf7:	data_out=16'h9f4;
17'hdcf8:	data_out=16'h367;
17'hdcf9:	data_out=16'h86b;
17'hdcfa:	data_out=16'h89e5;
17'hdcfb:	data_out=16'h8a00;
17'hdcfc:	data_out=16'h89fe;
17'hdcfd:	data_out=16'h89e8;
17'hdcfe:	data_out=16'h8a00;
17'hdcff:	data_out=16'h8a00;
17'hdd00:	data_out=16'h89fd;
17'hdd01:	data_out=16'h8a00;
17'hdd02:	data_out=16'h89e7;
17'hdd03:	data_out=16'h8984;
17'hdd04:	data_out=16'h888b;
17'hdd05:	data_out=16'h89f7;
17'hdd06:	data_out=16'h89e8;
17'hdd07:	data_out=16'ha00;
17'hdd08:	data_out=16'h9cd;
17'hdd09:	data_out=16'h9f4;
17'hdd0a:	data_out=16'h8a00;
17'hdd0b:	data_out=16'ha00;
17'hdd0c:	data_out=16'ha00;
17'hdd0d:	data_out=16'h89eb;
17'hdd0e:	data_out=16'h8a00;
17'hdd0f:	data_out=16'ha00;
17'hdd10:	data_out=16'h89ff;
17'hdd11:	data_out=16'h8a00;
17'hdd12:	data_out=16'h99f;
17'hdd13:	data_out=16'h79;
17'hdd14:	data_out=16'h89ee;
17'hdd15:	data_out=16'h8a00;
17'hdd16:	data_out=16'h897e;
17'hdd17:	data_out=16'h12a;
17'hdd18:	data_out=16'h8a00;
17'hdd19:	data_out=16'ha00;
17'hdd1a:	data_out=16'h89cc;
17'hdd1b:	data_out=16'h87f8;
17'hdd1c:	data_out=16'h8a00;
17'hdd1d:	data_out=16'h89c6;
17'hdd1e:	data_out=16'h89f9;
17'hdd1f:	data_out=16'h89f1;
17'hdd20:	data_out=16'h8a00;
17'hdd21:	data_out=16'h8a00;
17'hdd22:	data_out=16'h27;
17'hdd23:	data_out=16'h7a2;
17'hdd24:	data_out=16'h7b8;
17'hdd25:	data_out=16'h89da;
17'hdd26:	data_out=16'h9dc;
17'hdd27:	data_out=16'h82a4;
17'hdd28:	data_out=16'h89ff;
17'hdd29:	data_out=16'h8a00;
17'hdd2a:	data_out=16'ha00;
17'hdd2b:	data_out=16'ha00;
17'hdd2c:	data_out=16'h89fc;
17'hdd2d:	data_out=16'h9c7;
17'hdd2e:	data_out=16'ha00;
17'hdd2f:	data_out=16'h8703;
17'hdd30:	data_out=16'h3d9;
17'hdd31:	data_out=16'h8a00;
17'hdd32:	data_out=16'h301;
17'hdd33:	data_out=16'h89ff;
17'hdd34:	data_out=16'h89be;
17'hdd35:	data_out=16'h89dd;
17'hdd36:	data_out=16'h18d;
17'hdd37:	data_out=16'h8750;
17'hdd38:	data_out=16'h8a00;
17'hdd39:	data_out=16'h8a00;
17'hdd3a:	data_out=16'h9b1;
17'hdd3b:	data_out=16'ha00;
17'hdd3c:	data_out=16'h8a00;
17'hdd3d:	data_out=16'h8a00;
17'hdd3e:	data_out=16'h89ff;
17'hdd3f:	data_out=16'h89f9;
17'hdd40:	data_out=16'h8917;
17'hdd41:	data_out=16'h5b8;
17'hdd42:	data_out=16'ha00;
17'hdd43:	data_out=16'h3c8;
17'hdd44:	data_out=16'h89fd;
17'hdd45:	data_out=16'h8a00;
17'hdd46:	data_out=16'h89ff;
17'hdd47:	data_out=16'ha00;
17'hdd48:	data_out=16'h9f6;
17'hdd49:	data_out=16'h89fc;
17'hdd4a:	data_out=16'ha00;
17'hdd4b:	data_out=16'ha00;
17'hdd4c:	data_out=16'h960;
17'hdd4d:	data_out=16'h866b;
17'hdd4e:	data_out=16'ha00;
17'hdd4f:	data_out=16'h9e9;
17'hdd50:	data_out=16'h89c0;
17'hdd51:	data_out=16'h8a00;
17'hdd52:	data_out=16'h82a8;
17'hdd53:	data_out=16'h9eb;
17'hdd54:	data_out=16'h89fb;
17'hdd55:	data_out=16'h8944;
17'hdd56:	data_out=16'h89fc;
17'hdd57:	data_out=16'h8a00;
17'hdd58:	data_out=16'h8a00;
17'hdd59:	data_out=16'h89ea;
17'hdd5a:	data_out=16'h8348;
17'hdd5b:	data_out=16'h89fd;
17'hdd5c:	data_out=16'h8a00;
17'hdd5d:	data_out=16'h8231;
17'hdd5e:	data_out=16'h80ba;
17'hdd5f:	data_out=16'h891c;
17'hdd60:	data_out=16'h9d0;
17'hdd61:	data_out=16'h89fe;
17'hdd62:	data_out=16'ha00;
17'hdd63:	data_out=16'h89f7;
17'hdd64:	data_out=16'h89de;
17'hdd65:	data_out=16'h9c1;
17'hdd66:	data_out=16'ha00;
17'hdd67:	data_out=16'ha00;
17'hdd68:	data_out=16'h89ff;
17'hdd69:	data_out=16'h9d7;
17'hdd6a:	data_out=16'h8a00;
17'hdd6b:	data_out=16'h8a00;
17'hdd6c:	data_out=16'h89fc;
17'hdd6d:	data_out=16'h89f9;
17'hdd6e:	data_out=16'h8a00;
17'hdd6f:	data_out=16'h9fe;
17'hdd70:	data_out=16'h8a00;
17'hdd71:	data_out=16'ha00;
17'hdd72:	data_out=16'h8a00;
17'hdd73:	data_out=16'h8a00;
17'hdd74:	data_out=16'h363;
17'hdd75:	data_out=16'h8a00;
17'hdd76:	data_out=16'ha00;
17'hdd77:	data_out=16'h85d;
17'hdd78:	data_out=16'h82f2;
17'hdd79:	data_out=16'h809;
17'hdd7a:	data_out=16'h89df;
17'hdd7b:	data_out=16'h89ff;
17'hdd7c:	data_out=16'h89ff;
17'hdd7d:	data_out=16'h89ff;
17'hdd7e:	data_out=16'h889b;
17'hdd7f:	data_out=16'h8a00;
17'hdd80:	data_out=16'h89fd;
17'hdd81:	data_out=16'h85a0;
17'hdd82:	data_out=16'h89ff;
17'hdd83:	data_out=16'h89f5;
17'hdd84:	data_out=16'ha00;
17'hdd85:	data_out=16'h89e7;
17'hdd86:	data_out=16'h818e;
17'hdd87:	data_out=16'ha00;
17'hdd88:	data_out=16'h783;
17'hdd89:	data_out=16'h9fd;
17'hdd8a:	data_out=16'h899b;
17'hdd8b:	data_out=16'ha00;
17'hdd8c:	data_out=16'ha00;
17'hdd8d:	data_out=16'h89fd;
17'hdd8e:	data_out=16'h89ff;
17'hdd8f:	data_out=16'h175;
17'hdd90:	data_out=16'h8923;
17'hdd91:	data_out=16'h9b8;
17'hdd92:	data_out=16'h744;
17'hdd93:	data_out=16'h62a;
17'hdd94:	data_out=16'h89f1;
17'hdd95:	data_out=16'h8a00;
17'hdd96:	data_out=16'h89ae;
17'hdd97:	data_out=16'h83c0;
17'hdd98:	data_out=16'h8a00;
17'hdd99:	data_out=16'ha00;
17'hdd9a:	data_out=16'h834e;
17'hdd9b:	data_out=16'h89f5;
17'hdd9c:	data_out=16'h8a00;
17'hdd9d:	data_out=16'h9c9;
17'hdd9e:	data_out=16'h89ff;
17'hdd9f:	data_out=16'h8648;
17'hdda0:	data_out=16'h8a00;
17'hdda1:	data_out=16'h89ff;
17'hdda2:	data_out=16'h2a1;
17'hdda3:	data_out=16'h896;
17'hdda4:	data_out=16'h89e;
17'hdda5:	data_out=16'hb2;
17'hdda6:	data_out=16'h9ea;
17'hdda7:	data_out=16'h9eb;
17'hdda8:	data_out=16'h89fe;
17'hdda9:	data_out=16'h8a00;
17'hddaa:	data_out=16'ha00;
17'hddab:	data_out=16'ha00;
17'hddac:	data_out=16'h89fb;
17'hddad:	data_out=16'h9e9;
17'hddae:	data_out=16'ha00;
17'hddaf:	data_out=16'h8948;
17'hddb0:	data_out=16'h3f0;
17'hddb1:	data_out=16'h89fe;
17'hddb2:	data_out=16'h5b7;
17'hddb3:	data_out=16'h8a00;
17'hddb4:	data_out=16'h9be;
17'hddb5:	data_out=16'h74e;
17'hddb6:	data_out=16'h8867;
17'hddb7:	data_out=16'h89f6;
17'hddb8:	data_out=16'h8a00;
17'hddb9:	data_out=16'h8a00;
17'hddba:	data_out=16'h98d;
17'hddbb:	data_out=16'ha00;
17'hddbc:	data_out=16'h89fd;
17'hddbd:	data_out=16'h8a00;
17'hddbe:	data_out=16'h89fe;
17'hddbf:	data_out=16'h89e8;
17'hddc0:	data_out=16'h2e0;
17'hddc1:	data_out=16'h89ee;
17'hddc2:	data_out=16'ha00;
17'hddc3:	data_out=16'h81a9;
17'hddc4:	data_out=16'h88c2;
17'hddc5:	data_out=16'h8a00;
17'hddc6:	data_out=16'h8a00;
17'hddc7:	data_out=16'h9fc;
17'hddc8:	data_out=16'h9fa;
17'hddc9:	data_out=16'h858f;
17'hddca:	data_out=16'ha00;
17'hddcb:	data_out=16'ha00;
17'hddcc:	data_out=16'h92c;
17'hddcd:	data_out=16'h842e;
17'hddce:	data_out=16'ha00;
17'hddcf:	data_out=16'h9f2;
17'hddd0:	data_out=16'h89d9;
17'hddd1:	data_out=16'h8a00;
17'hddd2:	data_out=16'h893;
17'hddd3:	data_out=16'ha00;
17'hddd4:	data_out=16'h89fe;
17'hddd5:	data_out=16'h8975;
17'hddd6:	data_out=16'h89ff;
17'hddd7:	data_out=16'h8a00;
17'hddd8:	data_out=16'h8a00;
17'hddd9:	data_out=16'h89e5;
17'hddda:	data_out=16'h89f0;
17'hdddb:	data_out=16'h8860;
17'hdddc:	data_out=16'h89f2;
17'hdddd:	data_out=16'h8633;
17'hddde:	data_out=16'h8475;
17'hdddf:	data_out=16'h89ab;
17'hdde0:	data_out=16'h9f3;
17'hdde1:	data_out=16'h89e6;
17'hdde2:	data_out=16'ha00;
17'hdde3:	data_out=16'h89f9;
17'hdde4:	data_out=16'h9c8;
17'hdde5:	data_out=16'h9f2;
17'hdde6:	data_out=16'ha00;
17'hdde7:	data_out=16'h9ff;
17'hdde8:	data_out=16'h89fe;
17'hdde9:	data_out=16'h9da;
17'hddea:	data_out=16'h8a00;
17'hddeb:	data_out=16'h89f5;
17'hddec:	data_out=16'h89fc;
17'hdded:	data_out=16'h89fc;
17'hddee:	data_out=16'h8a00;
17'hddef:	data_out=16'h9fd;
17'hddf0:	data_out=16'h89ff;
17'hddf1:	data_out=16'h840;
17'hddf2:	data_out=16'h89fc;
17'hddf3:	data_out=16'h89e4;
17'hddf4:	data_out=16'h2aa;
17'hddf5:	data_out=16'h89f9;
17'hddf6:	data_out=16'ha00;
17'hddf7:	data_out=16'h804a;
17'hddf8:	data_out=16'h89c6;
17'hddf9:	data_out=16'h76c;
17'hddfa:	data_out=16'h89f2;
17'hddfb:	data_out=16'h89fe;
17'hddfc:	data_out=16'h8a00;
17'hddfd:	data_out=16'h8679;
17'hddfe:	data_out=16'h56c;
17'hddff:	data_out=16'h8a00;
17'hde00:	data_out=16'h9df;
17'hde01:	data_out=16'h9f9;
17'hde02:	data_out=16'h8a00;
17'hde03:	data_out=16'h89f1;
17'hde04:	data_out=16'ha00;
17'hde05:	data_out=16'h875b;
17'hde06:	data_out=16'h80cd;
17'hde07:	data_out=16'ha00;
17'hde08:	data_out=16'h8a00;
17'hde09:	data_out=16'ha00;
17'hde0a:	data_out=16'h9ff;
17'hde0b:	data_out=16'ha00;
17'hde0c:	data_out=16'ha00;
17'hde0d:	data_out=16'h8a00;
17'hde0e:	data_out=16'h8981;
17'hde0f:	data_out=16'h89e8;
17'hde10:	data_out=16'h913;
17'hde11:	data_out=16'ha00;
17'hde12:	data_out=16'h8a00;
17'hde13:	data_out=16'h8764;
17'hde14:	data_out=16'h89f2;
17'hde15:	data_out=16'h8a00;
17'hde16:	data_out=16'h89f8;
17'hde17:	data_out=16'h89e6;
17'hde18:	data_out=16'h8a00;
17'hde19:	data_out=16'ha00;
17'hde1a:	data_out=16'h9fe;
17'hde1b:	data_out=16'h89fb;
17'hde1c:	data_out=16'h8a00;
17'hde1d:	data_out=16'h9fc;
17'hde1e:	data_out=16'h89f7;
17'hde1f:	data_out=16'h89e8;
17'hde20:	data_out=16'h9f3;
17'hde21:	data_out=16'h8986;
17'hde22:	data_out=16'h9c1;
17'hde23:	data_out=16'h25;
17'hde24:	data_out=16'h29;
17'hde25:	data_out=16'h904;
17'hde26:	data_out=16'h49d;
17'hde27:	data_out=16'h9fe;
17'hde28:	data_out=16'h89fe;
17'hde29:	data_out=16'h8a00;
17'hde2a:	data_out=16'h84b4;
17'hde2b:	data_out=16'ha00;
17'hde2c:	data_out=16'h89f2;
17'hde2d:	data_out=16'h9fd;
17'hde2e:	data_out=16'h87c0;
17'hde2f:	data_out=16'h9fd;
17'hde30:	data_out=16'h7c7;
17'hde31:	data_out=16'h9ed;
17'hde32:	data_out=16'h9fd;
17'hde33:	data_out=16'h89fc;
17'hde34:	data_out=16'h9f1;
17'hde35:	data_out=16'h9f4;
17'hde36:	data_out=16'h89f5;
17'hde37:	data_out=16'h89f8;
17'hde38:	data_out=16'h96c;
17'hde39:	data_out=16'h8a00;
17'hde3a:	data_out=16'h9f3;
17'hde3b:	data_out=16'h9ff;
17'hde3c:	data_out=16'h89ee;
17'hde3d:	data_out=16'h96b;
17'hde3e:	data_out=16'h89fe;
17'hde3f:	data_out=16'h8758;
17'hde40:	data_out=16'ha00;
17'hde41:	data_out=16'h8a00;
17'hde42:	data_out=16'ha00;
17'hde43:	data_out=16'h861e;
17'hde44:	data_out=16'h9f6;
17'hde45:	data_out=16'h8a00;
17'hde46:	data_out=16'h8a00;
17'hde47:	data_out=16'h9fd;
17'hde48:	data_out=16'h9d6;
17'hde49:	data_out=16'h855;
17'hde4a:	data_out=16'ha00;
17'hde4b:	data_out=16'ha00;
17'hde4c:	data_out=16'h9e3;
17'hde4d:	data_out=16'h97f;
17'hde4e:	data_out=16'h203;
17'hde4f:	data_out=16'ha00;
17'hde50:	data_out=16'h8682;
17'hde51:	data_out=16'h8a00;
17'hde52:	data_out=16'h489;
17'hde53:	data_out=16'h9fc;
17'hde54:	data_out=16'h9f9;
17'hde55:	data_out=16'h89f5;
17'hde56:	data_out=16'h8a00;
17'hde57:	data_out=16'h8a00;
17'hde58:	data_out=16'h8a00;
17'hde59:	data_out=16'ha00;
17'hde5a:	data_out=16'h89fc;
17'hde5b:	data_out=16'h459;
17'hde5c:	data_out=16'h8152;
17'hde5d:	data_out=16'h80a6;
17'hde5e:	data_out=16'h9fe;
17'hde5f:	data_out=16'h86fe;
17'hde60:	data_out=16'h2ea;
17'hde61:	data_out=16'h9fb;
17'hde62:	data_out=16'h869e;
17'hde63:	data_out=16'h89f5;
17'hde64:	data_out=16'h9f6;
17'hde65:	data_out=16'ha00;
17'hde66:	data_out=16'ha00;
17'hde67:	data_out=16'ha00;
17'hde68:	data_out=16'h89a5;
17'hde69:	data_out=16'h8477;
17'hde6a:	data_out=16'h89fe;
17'hde6b:	data_out=16'h9ff;
17'hde6c:	data_out=16'h9e9;
17'hde6d:	data_out=16'h89f6;
17'hde6e:	data_out=16'h89fe;
17'hde6f:	data_out=16'h9fe;
17'hde70:	data_out=16'h8997;
17'hde71:	data_out=16'h89ea;
17'hde72:	data_out=16'h9ff;
17'hde73:	data_out=16'ha00;
17'hde74:	data_out=16'h56e;
17'hde75:	data_out=16'h89f6;
17'hde76:	data_out=16'ha00;
17'hde77:	data_out=16'h85d0;
17'hde78:	data_out=16'h89da;
17'hde79:	data_out=16'h888b;
17'hde7a:	data_out=16'h89f1;
17'hde7b:	data_out=16'h89fe;
17'hde7c:	data_out=16'h8a00;
17'hde7d:	data_out=16'h83a1;
17'hde7e:	data_out=16'h901;
17'hde7f:	data_out=16'h871b;
17'hde80:	data_out=16'ha00;
17'hde81:	data_out=16'ha00;
17'hde82:	data_out=16'h89fc;
17'hde83:	data_out=16'h2f0;
17'hde84:	data_out=16'ha00;
17'hde85:	data_out=16'ha00;
17'hde86:	data_out=16'h3ba;
17'hde87:	data_out=16'h821c;
17'hde88:	data_out=16'h89fe;
17'hde89:	data_out=16'h9ff;
17'hde8a:	data_out=16'ha00;
17'hde8b:	data_out=16'h87b0;
17'hde8c:	data_out=16'h8a00;
17'hde8d:	data_out=16'h8a00;
17'hde8e:	data_out=16'h8401;
17'hde8f:	data_out=16'h89f8;
17'hde90:	data_out=16'h99e;
17'hde91:	data_out=16'ha00;
17'hde92:	data_out=16'h8a00;
17'hde93:	data_out=16'h89f9;
17'hde94:	data_out=16'h89f6;
17'hde95:	data_out=16'h9bb;
17'hde96:	data_out=16'h89fa;
17'hde97:	data_out=16'h89f5;
17'hde98:	data_out=16'h8903;
17'hde99:	data_out=16'ha00;
17'hde9a:	data_out=16'ha00;
17'hde9b:	data_out=16'h89fa;
17'hde9c:	data_out=16'h830;
17'hde9d:	data_out=16'ha00;
17'hde9e:	data_out=16'h88b3;
17'hde9f:	data_out=16'h65d;
17'hdea0:	data_out=16'ha00;
17'hdea1:	data_out=16'h8418;
17'hdea2:	data_out=16'ha00;
17'hdea3:	data_out=16'h8a00;
17'hdea4:	data_out=16'h8a00;
17'hdea5:	data_out=16'ha00;
17'hdea6:	data_out=16'h89fa;
17'hdea7:	data_out=16'ha00;
17'hdea8:	data_out=16'h844c;
17'hdea9:	data_out=16'h8a00;
17'hdeaa:	data_out=16'h89f3;
17'hdeab:	data_out=16'ha00;
17'hdeac:	data_out=16'h82fc;
17'hdead:	data_out=16'h821e;
17'hdeae:	data_out=16'h89f4;
17'hdeaf:	data_out=16'ha00;
17'hdeb0:	data_out=16'h8730;
17'hdeb1:	data_out=16'ha00;
17'hdeb2:	data_out=16'h80a5;
17'hdeb3:	data_out=16'h8618;
17'hdeb4:	data_out=16'ha00;
17'hdeb5:	data_out=16'ha00;
17'hdeb6:	data_out=16'h89f9;
17'hdeb7:	data_out=16'h89fa;
17'hdeb8:	data_out=16'ha00;
17'hdeb9:	data_out=16'h8488;
17'hdeba:	data_out=16'h9fb;
17'hdebb:	data_out=16'h40f;
17'hdebc:	data_out=16'h89ee;
17'hdebd:	data_out=16'ha00;
17'hdebe:	data_out=16'h8450;
17'hdebf:	data_out=16'ha00;
17'hdec0:	data_out=16'ha00;
17'hdec1:	data_out=16'h89fd;
17'hdec2:	data_out=16'h586;
17'hdec3:	data_out=16'h806e;
17'hdec4:	data_out=16'ha00;
17'hdec5:	data_out=16'h953;
17'hdec6:	data_out=16'h89fb;
17'hdec7:	data_out=16'h9fc;
17'hdec8:	data_out=16'h8151;
17'hdec9:	data_out=16'ha00;
17'hdeca:	data_out=16'h1a9;
17'hdecb:	data_out=16'h879e;
17'hdecc:	data_out=16'h8d5;
17'hdecd:	data_out=16'ha00;
17'hdece:	data_out=16'h88b1;
17'hdecf:	data_out=16'h9ea;
17'hded0:	data_out=16'ha00;
17'hded1:	data_out=16'h8a00;
17'hded2:	data_out=16'h8764;
17'hded3:	data_out=16'h83b;
17'hded4:	data_out=16'ha00;
17'hded5:	data_out=16'h89fa;
17'hded6:	data_out=16'h901;
17'hded7:	data_out=16'ha00;
17'hded8:	data_out=16'h89ff;
17'hded9:	data_out=16'ha00;
17'hdeda:	data_out=16'h89ff;
17'hdedb:	data_out=16'ha00;
17'hdedc:	data_out=16'h720;
17'hdedd:	data_out=16'h82a4;
17'hdede:	data_out=16'ha00;
17'hdedf:	data_out=16'h1e6;
17'hdee0:	data_out=16'h89fc;
17'hdee1:	data_out=16'ha00;
17'hdee2:	data_out=16'h89f0;
17'hdee3:	data_out=16'h875c;
17'hdee4:	data_out=16'ha00;
17'hdee5:	data_out=16'ha00;
17'hdee6:	data_out=16'ha00;
17'hdee7:	data_out=16'h305;
17'hdee8:	data_out=16'h8421;
17'hdee9:	data_out=16'h8a00;
17'hdeea:	data_out=16'h83e5;
17'hdeeb:	data_out=16'ha00;
17'hdeec:	data_out=16'h831a;
17'hdeed:	data_out=16'h86ad;
17'hdeee:	data_out=16'h83e7;
17'hdeef:	data_out=16'h8f6;
17'hdef0:	data_out=16'h83ff;
17'hdef1:	data_out=16'h89fa;
17'hdef2:	data_out=16'ha00;
17'hdef3:	data_out=16'ha00;
17'hdef4:	data_out=16'h897f;
17'hdef5:	data_out=16'h89f7;
17'hdef6:	data_out=16'ha00;
17'hdef7:	data_out=16'ha00;
17'hdef8:	data_out=16'h81b9;
17'hdef9:	data_out=16'h89fd;
17'hdefa:	data_out=16'h89f7;
17'hdefb:	data_out=16'h8453;
17'hdefc:	data_out=16'h83e0;
17'hdefd:	data_out=16'h41d;
17'hdefe:	data_out=16'ha00;
17'hdeff:	data_out=16'ha00;
17'hdf00:	data_out=16'ha00;
17'hdf01:	data_out=16'h881;
17'hdf02:	data_out=16'h8a00;
17'hdf03:	data_out=16'h3c1;
17'hdf04:	data_out=16'ha00;
17'hdf05:	data_out=16'h7e7;
17'hdf06:	data_out=16'h1ac;
17'hdf07:	data_out=16'h81af;
17'hdf08:	data_out=16'h89ff;
17'hdf09:	data_out=16'ha00;
17'hdf0a:	data_out=16'h6c9;
17'hdf0b:	data_out=16'h8876;
17'hdf0c:	data_out=16'h8a00;
17'hdf0d:	data_out=16'h89b2;
17'hdf0e:	data_out=16'h8161;
17'hdf0f:	data_out=16'h89ff;
17'hdf10:	data_out=16'h577;
17'hdf11:	data_out=16'ha00;
17'hdf12:	data_out=16'h858b;
17'hdf13:	data_out=16'h838a;
17'hdf14:	data_out=16'h55e;
17'hdf15:	data_out=16'h590;
17'hdf16:	data_out=16'h8405;
17'hdf17:	data_out=16'h82cc;
17'hdf18:	data_out=16'h8048;
17'hdf19:	data_out=16'h751;
17'hdf1a:	data_out=16'h4f9;
17'hdf1b:	data_out=16'h8596;
17'hdf1c:	data_out=16'h9ab;
17'hdf1d:	data_out=16'ha00;
17'hdf1e:	data_out=16'h394;
17'hdf1f:	data_out=16'ha00;
17'hdf20:	data_out=16'ha00;
17'hdf21:	data_out=16'h816c;
17'hdf22:	data_out=16'ha00;
17'hdf23:	data_out=16'h86d0;
17'hdf24:	data_out=16'h86cd;
17'hdf25:	data_out=16'hfd;
17'hdf26:	data_out=16'h8719;
17'hdf27:	data_out=16'ha00;
17'hdf28:	data_out=16'h8179;
17'hdf29:	data_out=16'h88;
17'hdf2a:	data_out=16'h89ff;
17'hdf2b:	data_out=16'ha00;
17'hdf2c:	data_out=16'h8076;
17'hdf2d:	data_out=16'h867b;
17'hdf2e:	data_out=16'h89ff;
17'hdf2f:	data_out=16'h8fd;
17'hdf30:	data_out=16'h8a00;
17'hdf31:	data_out=16'ha00;
17'hdf32:	data_out=16'h8a00;
17'hdf33:	data_out=16'ha00;
17'hdf34:	data_out=16'h9fd;
17'hdf35:	data_out=16'h85ad;
17'hdf36:	data_out=16'h85a3;
17'hdf37:	data_out=16'h8a00;
17'hdf38:	data_out=16'ha00;
17'hdf39:	data_out=16'ha00;
17'hdf3a:	data_out=16'h9e5;
17'hdf3b:	data_out=16'hf;
17'hdf3c:	data_out=16'h8a00;
17'hdf3d:	data_out=16'ha00;
17'hdf3e:	data_out=16'h817a;
17'hdf3f:	data_out=16'h781;
17'hdf40:	data_out=16'h4a1;
17'hdf41:	data_out=16'h8a00;
17'hdf42:	data_out=16'h8a00;
17'hdf43:	data_out=16'h11d;
17'hdf44:	data_out=16'ha00;
17'hdf45:	data_out=16'h55c;
17'hdf46:	data_out=16'h8a00;
17'hdf47:	data_out=16'h535;
17'hdf48:	data_out=16'h5e;
17'hdf49:	data_out=16'h1a5;
17'hdf4a:	data_out=16'h85cf;
17'hdf4b:	data_out=16'h8a00;
17'hdf4c:	data_out=16'h83dd;
17'hdf4d:	data_out=16'ha00;
17'hdf4e:	data_out=16'h89ff;
17'hdf4f:	data_out=16'h812e;
17'hdf50:	data_out=16'h4f8;
17'hdf51:	data_out=16'h8a00;
17'hdf52:	data_out=16'h8527;
17'hdf53:	data_out=16'h935;
17'hdf54:	data_out=16'ha00;
17'hdf55:	data_out=16'h89ff;
17'hdf56:	data_out=16'h7ba;
17'hdf57:	data_out=16'ha00;
17'hdf58:	data_out=16'h8a00;
17'hdf59:	data_out=16'h65e;
17'hdf5a:	data_out=16'h8a00;
17'hdf5b:	data_out=16'ha00;
17'hdf5c:	data_out=16'h93c;
17'hdf5d:	data_out=16'h84d1;
17'hdf5e:	data_out=16'h721;
17'hdf5f:	data_out=16'h205;
17'hdf60:	data_out=16'h8976;
17'hdf61:	data_out=16'h9e7;
17'hdf62:	data_out=16'h8a00;
17'hdf63:	data_out=16'h9fa;
17'hdf64:	data_out=16'ha00;
17'hdf65:	data_out=16'h745;
17'hdf66:	data_out=16'h77a;
17'hdf67:	data_out=16'h260;
17'hdf68:	data_out=16'h816e;
17'hdf69:	data_out=16'h89ff;
17'hdf6a:	data_out=16'h8156;
17'hdf6b:	data_out=16'ha00;
17'hdf6c:	data_out=16'h8444;
17'hdf6d:	data_out=16'ha00;
17'hdf6e:	data_out=16'h8157;
17'hdf6f:	data_out=16'h8589;
17'hdf70:	data_out=16'h815f;
17'hdf71:	data_out=16'h87fe;
17'hdf72:	data_out=16'ha00;
17'hdf73:	data_out=16'ha00;
17'hdf74:	data_out=16'h8a00;
17'hdf75:	data_out=16'h8a00;
17'hdf76:	data_out=16'ha00;
17'hdf77:	data_out=16'h441;
17'hdf78:	data_out=16'h80cb;
17'hdf79:	data_out=16'h89ff;
17'hdf7a:	data_out=16'h6b9;
17'hdf7b:	data_out=16'h817c;
17'hdf7c:	data_out=16'hfc;
17'hdf7d:	data_out=16'h577;
17'hdf7e:	data_out=16'ha00;
17'hdf7f:	data_out=16'h859;
17'hdf80:	data_out=16'h457;
17'hdf81:	data_out=16'h1e1;
17'hdf82:	data_out=16'h82e9;
17'hdf83:	data_out=16'h30;
17'hdf84:	data_out=16'hb4;
17'hdf85:	data_out=16'hdc;
17'hdf86:	data_out=16'h8100;
17'hdf87:	data_out=16'h80c1;
17'hdf88:	data_out=16'h8164;
17'hdf89:	data_out=16'h234;
17'hdf8a:	data_out=16'h100;
17'hdf8b:	data_out=16'h81c5;
17'hdf8c:	data_out=16'h8497;
17'hdf8d:	data_out=16'h80aa;
17'hdf8e:	data_out=16'h805a;
17'hdf8f:	data_out=16'h815e;
17'hdf90:	data_out=16'h5b;
17'hdf91:	data_out=16'h245;
17'hdf92:	data_out=16'h8296;
17'hdf93:	data_out=16'h50;
17'hdf94:	data_out=16'h8092;
17'hdf95:	data_out=16'h1a0;
17'hdf96:	data_out=16'h6f;
17'hdf97:	data_out=16'h8197;
17'hdf98:	data_out=16'h8031;
17'hdf99:	data_out=16'h24d;
17'hdf9a:	data_out=16'h3b;
17'hdf9b:	data_out=16'h1a;
17'hdf9c:	data_out=16'h363;
17'hdf9d:	data_out=16'h164;
17'hdf9e:	data_out=16'h91;
17'hdf9f:	data_out=16'h8065;
17'hdfa0:	data_out=16'h482;
17'hdfa1:	data_out=16'h805d;
17'hdfa2:	data_out=16'h152;
17'hdfa3:	data_out=16'h81da;
17'hdfa4:	data_out=16'h81d8;
17'hdfa5:	data_out=16'h802c;
17'hdfa6:	data_out=16'h8067;
17'hdfa7:	data_out=16'h19e;
17'hdfa8:	data_out=16'h8057;
17'hdfa9:	data_out=16'he;
17'hdfaa:	data_out=16'h8269;
17'hdfab:	data_out=16'h69c;
17'hdfac:	data_out=16'h14;
17'hdfad:	data_out=16'h80d6;
17'hdfae:	data_out=16'h82ee;
17'hdfaf:	data_out=16'h201;
17'hdfb0:	data_out=16'h8203;
17'hdfb1:	data_out=16'h44e;
17'hdfb2:	data_out=16'h81aa;
17'hdfb3:	data_out=16'h9b;
17'hdfb4:	data_out=16'h44a;
17'hdfb5:	data_out=16'h8192;
17'hdfb6:	data_out=16'h81d8;
17'hdfb7:	data_out=16'h82ed;
17'hdfb8:	data_out=16'h637;
17'hdfb9:	data_out=16'h1c4;
17'hdfba:	data_out=16'h801e;
17'hdfbb:	data_out=16'h173;
17'hdfbc:	data_out=16'h8325;
17'hdfbd:	data_out=16'h663;
17'hdfbe:	data_out=16'h8059;
17'hdfbf:	data_out=16'h107;
17'hdfc0:	data_out=16'h5;
17'hdfc1:	data_out=16'h8283;
17'hdfc2:	data_out=16'h81d7;
17'hdfc3:	data_out=16'h810d;
17'hdfc4:	data_out=16'h1de;
17'hdfc5:	data_out=16'h199;
17'hdfc6:	data_out=16'h818b;
17'hdfc7:	data_out=16'h80f6;
17'hdfc8:	data_out=16'h819f;
17'hdfc9:	data_out=16'h1;
17'hdfca:	data_out=16'h8218;
17'hdfcb:	data_out=16'h8450;
17'hdfcc:	data_out=16'h8180;
17'hdfcd:	data_out=16'h249;
17'hdfce:	data_out=16'h8187;
17'hdfcf:	data_out=16'h812f;
17'hdfd0:	data_out=16'h8034;
17'hdfd1:	data_out=16'h80e0;
17'hdfd2:	data_out=16'h814b;
17'hdfd3:	data_out=16'h118;
17'hdfd4:	data_out=16'h26e;
17'hdfd5:	data_out=16'h834e;
17'hdfd6:	data_out=16'h8064;
17'hdfd7:	data_out=16'h8016;
17'hdfd8:	data_out=16'h838e;
17'hdfd9:	data_out=16'h8001;
17'hdfda:	data_out=16'h8287;
17'hdfdb:	data_out=16'hff;
17'hdfdc:	data_out=16'hb9;
17'hdfdd:	data_out=16'h8065;
17'hdfde:	data_out=16'h110;
17'hdfdf:	data_out=16'h3f;
17'hdfe0:	data_out=16'h80c8;
17'hdfe1:	data_out=16'h2a5;
17'hdfe2:	data_out=16'h82e0;
17'hdfe3:	data_out=16'h43;
17'hdfe4:	data_out=16'h518;
17'hdfe5:	data_out=16'h11b;
17'hdfe6:	data_out=16'h1a2;
17'hdfe7:	data_out=16'h80e4;
17'hdfe8:	data_out=16'h805e;
17'hdfe9:	data_out=16'h833f;
17'hdfea:	data_out=16'h806c;
17'hdfeb:	data_out=16'h345;
17'hdfec:	data_out=16'h8076;
17'hdfed:	data_out=16'hae;
17'hdfee:	data_out=16'h8067;
17'hdfef:	data_out=16'h8071;
17'hdff0:	data_out=16'h8067;
17'hdff1:	data_out=16'h82e4;
17'hdff2:	data_out=16'h18e;
17'hdff3:	data_out=16'h319;
17'hdff4:	data_out=16'h821e;
17'hdff5:	data_out=16'h821d;
17'hdff6:	data_out=16'h414;
17'hdff7:	data_out=16'h8075;
17'hdff8:	data_out=16'h98;
17'hdff9:	data_out=16'h83af;
17'hdffa:	data_out=16'h8067;
17'hdffb:	data_out=16'h8055;
17'hdffc:	data_out=16'h80d5;
17'hdffd:	data_out=16'h80c7;
17'hdffe:	data_out=16'h237;
17'hdfff:	data_out=16'h35;
17'he000:	data_out=16'h8023;
17'he001:	data_out=16'h800c;
17'he002:	data_out=16'h8;
17'he003:	data_out=16'hd;
17'he004:	data_out=16'h800c;
17'he005:	data_out=16'h800c;
17'he006:	data_out=16'h6;
17'he007:	data_out=16'h2;
17'he008:	data_out=16'h801a;
17'he009:	data_out=16'h8016;
17'he00a:	data_out=16'h8012;
17'he00b:	data_out=16'h8009;
17'he00c:	data_out=16'h8006;
17'he00d:	data_out=16'h8009;
17'he00e:	data_out=16'h8006;
17'he00f:	data_out=16'h8005;
17'he010:	data_out=16'h0;
17'he011:	data_out=16'h8005;
17'he012:	data_out=16'h24;
17'he013:	data_out=16'h800b;
17'he014:	data_out=16'h3c;
17'he015:	data_out=16'h801f;
17'he016:	data_out=16'h8015;
17'he017:	data_out=16'h43;
17'he018:	data_out=16'h8019;
17'he019:	data_out=16'h8012;
17'he01a:	data_out=16'h8019;
17'he01b:	data_out=16'he;
17'he01c:	data_out=16'h15;
17'he01d:	data_out=16'h1d;
17'he01e:	data_out=16'h26;
17'he01f:	data_out=16'h8010;
17'he020:	data_out=16'h4;
17'he021:	data_out=16'h800e;
17'he022:	data_out=16'h2d;
17'he023:	data_out=16'h8012;
17'he024:	data_out=16'h8019;
17'he025:	data_out=16'he;
17'he026:	data_out=16'h800f;
17'he027:	data_out=16'he;
17'he028:	data_out=16'h8006;
17'he029:	data_out=16'h5;
17'he02a:	data_out=16'h8003;
17'he02b:	data_out=16'h14;
17'he02c:	data_out=16'h801d;
17'he02d:	data_out=16'h9;
17'he02e:	data_out=16'h8;
17'he02f:	data_out=16'h14;
17'he030:	data_out=16'h8014;
17'he031:	data_out=16'h8007;
17'he032:	data_out=16'h8014;
17'he033:	data_out=16'h36;
17'he034:	data_out=16'h8009;
17'he035:	data_out=16'h802d;
17'he036:	data_out=16'h8018;
17'he037:	data_out=16'h1a;
17'he038:	data_out=16'h800e;
17'he039:	data_out=16'h3;
17'he03a:	data_out=16'h12;
17'he03b:	data_out=16'h802a;
17'he03c:	data_out=16'h12;
17'he03d:	data_out=16'h801d;
17'he03e:	data_out=16'h8004;
17'he03f:	data_out=16'h801b;
17'he040:	data_out=16'h13;
17'he041:	data_out=16'h16;
17'he042:	data_out=16'h8005;
17'he043:	data_out=16'h8007;
17'he044:	data_out=16'h801a;
17'he045:	data_out=16'h801e;
17'he046:	data_out=16'h16;
17'he047:	data_out=16'hf;
17'he048:	data_out=16'h1b;
17'he049:	data_out=16'hd;
17'he04a:	data_out=16'h800a;
17'he04b:	data_out=16'hb;
17'he04c:	data_out=16'h1;
17'he04d:	data_out=16'h28;
17'he04e:	data_out=16'h8010;
17'he04f:	data_out=16'h8008;
17'he050:	data_out=16'h16;
17'he051:	data_out=16'h802b;
17'he052:	data_out=16'h8029;
17'he053:	data_out=16'h3f;
17'he054:	data_out=16'h8002;
17'he055:	data_out=16'h8004;
17'he056:	data_out=16'h14;
17'he057:	data_out=16'h0;
17'he058:	data_out=16'he;
17'he059:	data_out=16'h3;
17'he05a:	data_out=16'h15;
17'he05b:	data_out=16'h8039;
17'he05c:	data_out=16'h8003;
17'he05d:	data_out=16'h1;
17'he05e:	data_out=16'h4;
17'he05f:	data_out=16'h8005;
17'he060:	data_out=16'h800f;
17'he061:	data_out=16'h8030;
17'he062:	data_out=16'he;
17'he063:	data_out=16'h2c;
17'he064:	data_out=16'h4;
17'he065:	data_out=16'h10;
17'he066:	data_out=16'h8007;
17'he067:	data_out=16'h13;
17'he068:	data_out=16'h800c;
17'he069:	data_out=16'h8005;
17'he06a:	data_out=16'h8004;
17'he06b:	data_out=16'h800a;
17'he06c:	data_out=16'h19;
17'he06d:	data_out=16'h30;
17'he06e:	data_out=16'h800a;
17'he06f:	data_out=16'h23;
17'he070:	data_out=16'h800b;
17'he071:	data_out=16'h8009;
17'he072:	data_out=16'h800d;
17'he073:	data_out=16'h8005;
17'he074:	data_out=16'h8019;
17'he075:	data_out=16'h8005;
17'he076:	data_out=16'h8009;
17'he077:	data_out=16'h800a;
17'he078:	data_out=16'h8004;
17'he079:	data_out=16'h8002;
17'he07a:	data_out=16'h3d;
17'he07b:	data_out=16'h8010;
17'he07c:	data_out=16'h8018;
17'he07d:	data_out=16'h800a;
17'he07e:	data_out=16'h8005;
17'he07f:	data_out=16'h801e;
17'he080:	data_out=16'h814d;
17'he081:	data_out=16'h800e;
17'he082:	data_out=16'h8067;
17'he083:	data_out=16'h80a3;
17'he084:	data_out=16'h8081;
17'he085:	data_out=16'h84;
17'he086:	data_out=16'h19;
17'he087:	data_out=16'h80cd;
17'he088:	data_out=16'h18;
17'he089:	data_out=16'h8162;
17'he08a:	data_out=16'h808e;
17'he08b:	data_out=16'h92;
17'he08c:	data_out=16'h6f;
17'he08d:	data_out=16'h8093;
17'he08e:	data_out=16'h8022;
17'he08f:	data_out=16'h805b;
17'he090:	data_out=16'h816e;
17'he091:	data_out=16'h802f;
17'he092:	data_out=16'h8092;
17'he093:	data_out=16'h8122;
17'he094:	data_out=16'h8025;
17'he095:	data_out=16'h80b4;
17'he096:	data_out=16'h80dd;
17'he097:	data_out=16'h800c;
17'he098:	data_out=16'h8079;
17'he099:	data_out=16'h3;
17'he09a:	data_out=16'h807a;
17'he09b:	data_out=16'h98;
17'he09c:	data_out=16'h7b;
17'he09d:	data_out=16'h8011;
17'he09e:	data_out=16'h8024;
17'he09f:	data_out=16'h8027;
17'he0a0:	data_out=16'h36;
17'he0a1:	data_out=16'h8021;
17'he0a2:	data_out=16'h8166;
17'he0a3:	data_out=16'h8077;
17'he0a4:	data_out=16'h8076;
17'he0a5:	data_out=16'h8132;
17'he0a6:	data_out=16'h80f1;
17'he0a7:	data_out=16'h4f;
17'he0a8:	data_out=16'h8012;
17'he0a9:	data_out=16'h80c7;
17'he0aa:	data_out=16'h812d;
17'he0ab:	data_out=16'h24;
17'he0ac:	data_out=16'h8094;
17'he0ad:	data_out=16'h81bb;
17'he0ae:	data_out=16'h80e4;
17'he0af:	data_out=16'h800f;
17'he0b0:	data_out=16'h8039;
17'he0b1:	data_out=16'h1a;
17'he0b2:	data_out=16'h803b;
17'he0b3:	data_out=16'h801d;
17'he0b4:	data_out=16'h8057;
17'he0b5:	data_out=16'h87;
17'he0b6:	data_out=16'h1d;
17'he0b7:	data_out=16'h8055;
17'he0b8:	data_out=16'h4f;
17'he0b9:	data_out=16'h8016;
17'he0ba:	data_out=16'h81d9;
17'he0bb:	data_out=16'h19;
17'he0bc:	data_out=16'h38;
17'he0bd:	data_out=16'h8149;
17'he0be:	data_out=16'h8018;
17'he0bf:	data_out=16'h1c;
17'he0c0:	data_out=16'h81a1;
17'he0c1:	data_out=16'ha9;
17'he0c2:	data_out=16'h8140;
17'he0c3:	data_out=16'h49;
17'he0c4:	data_out=16'h805d;
17'he0c5:	data_out=16'h80d1;
17'he0c6:	data_out=16'h2f;
17'he0c7:	data_out=16'h81ad;
17'he0c8:	data_out=16'h80bc;
17'he0c9:	data_out=16'h8144;
17'he0ca:	data_out=16'h80c7;
17'he0cb:	data_out=16'h8071;
17'he0cc:	data_out=16'h8186;
17'he0cd:	data_out=16'h8140;
17'he0ce:	data_out=16'h80cd;
17'he0cf:	data_out=16'h8192;
17'he0d0:	data_out=16'h8182;
17'he0d1:	data_out=16'h37;
17'he0d2:	data_out=16'h8092;
17'he0d3:	data_out=16'h116;
17'he0d4:	data_out=16'h8029;
17'he0d5:	data_out=16'h85;
17'he0d6:	data_out=16'h8176;
17'he0d7:	data_out=16'h81b8;
17'he0d8:	data_out=16'h18;
17'he0d9:	data_out=16'h81cd;
17'he0da:	data_out=16'hee;
17'he0db:	data_out=16'hef;
17'he0dc:	data_out=16'ha8;
17'he0dd:	data_out=16'h811e;
17'he0de:	data_out=16'h802f;
17'he0df:	data_out=16'h8074;
17'he0e0:	data_out=16'h815d;
17'he0e1:	data_out=16'h800e;
17'he0e2:	data_out=16'he9;
17'he0e3:	data_out=16'h8019;
17'he0e4:	data_out=16'h809d;
17'he0e5:	data_out=16'h8093;
17'he0e6:	data_out=16'h800f;
17'he0e7:	data_out=16'h80cd;
17'he0e8:	data_out=16'h801f;
17'he0e9:	data_out=16'h8024;
17'he0ea:	data_out=16'h801e;
17'he0eb:	data_out=16'h806e;
17'he0ec:	data_out=16'h81ff;
17'he0ed:	data_out=16'h8020;
17'he0ee:	data_out=16'h801d;
17'he0ef:	data_out=16'h8022;
17'he0f0:	data_out=16'h8023;
17'he0f1:	data_out=16'h8086;
17'he0f2:	data_out=16'h80e8;
17'he0f3:	data_out=16'h805b;
17'he0f4:	data_out=16'h8034;
17'he0f5:	data_out=16'h10a;
17'he0f6:	data_out=16'h1f;
17'he0f7:	data_out=16'h81ea;
17'he0f8:	data_out=16'h4a;
17'he0f9:	data_out=16'h80dc;
17'he0fa:	data_out=16'h8020;
17'he0fb:	data_out=16'h801e;
17'he0fc:	data_out=16'h1d;
17'he0fd:	data_out=16'he7;
17'he0fe:	data_out=16'h8137;
17'he0ff:	data_out=16'h8199;
17'he100:	data_out=16'h8648;
17'he101:	data_out=16'h8001;
17'he102:	data_out=16'h828e;
17'he103:	data_out=16'h83ca;
17'he104:	data_out=16'h815c;
17'he105:	data_out=16'h424;
17'he106:	data_out=16'h1ca;
17'he107:	data_out=16'h840f;
17'he108:	data_out=16'h83da;
17'he109:	data_out=16'h8700;
17'he10a:	data_out=16'h82dc;
17'he10b:	data_out=16'h272;
17'he10c:	data_out=16'h80bd;
17'he10d:	data_out=16'h823e;
17'he10e:	data_out=16'h8148;
17'he10f:	data_out=16'h8248;
17'he110:	data_out=16'h8684;
17'he111:	data_out=16'hd6;
17'he112:	data_out=16'h81fb;
17'he113:	data_out=16'h845f;
17'he114:	data_out=16'h12a;
17'he115:	data_out=16'h82af;
17'he116:	data_out=16'h843d;
17'he117:	data_out=16'h17c;
17'he118:	data_out=16'h81e7;
17'he119:	data_out=16'h251;
17'he11a:	data_out=16'h80a8;
17'he11b:	data_out=16'h3c7;
17'he11c:	data_out=16'h37e;
17'he11d:	data_out=16'h1c4;
17'he11e:	data_out=16'h9b;
17'he11f:	data_out=16'h8123;
17'he120:	data_out=16'h3ff;
17'he121:	data_out=16'h812f;
17'he122:	data_out=16'h85dc;
17'he123:	data_out=16'h8406;
17'he124:	data_out=16'h8406;
17'he125:	data_out=16'h8658;
17'he126:	data_out=16'h889a;
17'he127:	data_out=16'h36e;
17'he128:	data_out=16'h80fc;
17'he129:	data_out=16'h84bb;
17'he12a:	data_out=16'h883c;
17'he12b:	data_out=16'h492;
17'he12c:	data_out=16'h83bd;
17'he12d:	data_out=16'h8a00;
17'he12e:	data_out=16'h847a;
17'he12f:	data_out=16'h173;
17'he130:	data_out=16'h8264;
17'he131:	data_out=16'h25d;
17'he132:	data_out=16'h826a;
17'he133:	data_out=16'h8d;
17'he134:	data_out=16'h2b;
17'he135:	data_out=16'h29d;
17'he136:	data_out=16'h8294;
17'he137:	data_out=16'h8206;
17'he138:	data_out=16'h441;
17'he139:	data_out=16'h1c0;
17'he13a:	data_out=16'h880d;
17'he13b:	data_out=16'h80d9;
17'he13c:	data_out=16'h8121;
17'he13d:	data_out=16'h83bb;
17'he13e:	data_out=16'h8106;
17'he13f:	data_out=16'h3dd;
17'he140:	data_out=16'h863d;
17'he141:	data_out=16'hfb;
17'he142:	data_out=16'h8993;
17'he143:	data_out=16'h210;
17'he144:	data_out=16'h21;
17'he145:	data_out=16'h82c7;
17'he146:	data_out=16'h81bf;
17'he147:	data_out=16'h885a;
17'he148:	data_out=16'h8180;
17'he149:	data_out=16'h8650;
17'he14a:	data_out=16'h83bf;
17'he14b:	data_out=16'h8425;
17'he14c:	data_out=16'h87a7;
17'he14d:	data_out=16'h85be;
17'he14e:	data_out=16'h8455;
17'he14f:	data_out=16'h877c;
17'he150:	data_out=16'h85f8;
17'he151:	data_out=16'h1f;
17'he152:	data_out=16'h85a7;
17'he153:	data_out=16'h670;
17'he154:	data_out=16'h30;
17'he155:	data_out=16'h80b5;
17'he156:	data_out=16'h87b5;
17'he157:	data_out=16'h87ef;
17'he158:	data_out=16'h811e;
17'he159:	data_out=16'h8711;
17'he15a:	data_out=16'h3b8;
17'he15b:	data_out=16'h4cd;
17'he15c:	data_out=16'h5a7;
17'he15d:	data_out=16'h853f;
17'he15e:	data_out=16'hd0;
17'he15f:	data_out=16'h81c6;
17'he160:	data_out=16'h898f;
17'he161:	data_out=16'h23f;
17'he162:	data_out=16'h332;
17'he163:	data_out=16'h118;
17'he164:	data_out=16'h6c;
17'he165:	data_out=16'h4f;
17'he166:	data_out=16'h2ef;
17'he167:	data_out=16'h8459;
17'he168:	data_out=16'h8126;
17'he169:	data_out=16'h84e5;
17'he16a:	data_out=16'h8151;
17'he16b:	data_out=16'h113;
17'he16c:	data_out=16'h89ff;
17'he16d:	data_out=16'he1;
17'he16e:	data_out=16'h8159;
17'he16f:	data_out=16'h8227;
17'he170:	data_out=16'h8148;
17'he171:	data_out=16'h8207;
17'he172:	data_out=16'h8385;
17'he173:	data_out=16'h80dc;
17'he174:	data_out=16'h826c;
17'he175:	data_out=16'h6b7;
17'he176:	data_out=16'h26e;
17'he177:	data_out=16'h890a;
17'he178:	data_out=16'h311;
17'he179:	data_out=16'h855f;
17'he17a:	data_out=16'h15c;
17'he17b:	data_out=16'h8101;
17'he17c:	data_out=16'h80f8;
17'he17d:	data_out=16'h429;
17'he17e:	data_out=16'h861b;
17'he17f:	data_out=16'h862c;
17'he180:	data_out=16'h84e0;
17'he181:	data_out=16'h8083;
17'he182:	data_out=16'h8838;
17'he183:	data_out=16'h8a00;
17'he184:	data_out=16'h83ac;
17'he185:	data_out=16'h9f0;
17'he186:	data_out=16'h2bf;
17'he187:	data_out=16'h8a00;
17'he188:	data_out=16'h886e;
17'he189:	data_out=16'h8a00;
17'he18a:	data_out=16'h89ff;
17'he18b:	data_out=16'h136;
17'he18c:	data_out=16'h8a00;
17'he18d:	data_out=16'h8601;
17'he18e:	data_out=16'h8108;
17'he18f:	data_out=16'h8a00;
17'he190:	data_out=16'h8606;
17'he191:	data_out=16'h817b;
17'he192:	data_out=16'h84ca;
17'he193:	data_out=16'h8949;
17'he194:	data_out=16'h9f8;
17'he195:	data_out=16'h860d;
17'he196:	data_out=16'h8a00;
17'he197:	data_out=16'h9ab;
17'he198:	data_out=16'h8056;
17'he199:	data_out=16'h626;
17'he19a:	data_out=16'h8671;
17'he19b:	data_out=16'h9f4;
17'he19c:	data_out=16'h9e7;
17'he19d:	data_out=16'h5ea;
17'he19e:	data_out=16'h9a5;
17'he19f:	data_out=16'h60;
17'he1a0:	data_out=16'ha00;
17'he1a1:	data_out=16'h80fc;
17'he1a2:	data_out=16'hbf;
17'he1a3:	data_out=16'h8a00;
17'he1a4:	data_out=16'h8a00;
17'he1a5:	data_out=16'h8a00;
17'he1a6:	data_out=16'h8a00;
17'he1a7:	data_out=16'ha00;
17'he1a8:	data_out=16'h80e3;
17'he1a9:	data_out=16'h8882;
17'he1aa:	data_out=16'h8a00;
17'he1ab:	data_out=16'ha00;
17'he1ac:	data_out=16'h8a00;
17'he1ad:	data_out=16'h89fe;
17'he1ae:	data_out=16'h89c1;
17'he1af:	data_out=16'h9fe;
17'he1b0:	data_out=16'h8a00;
17'he1b1:	data_out=16'h525;
17'he1b2:	data_out=16'h8a00;
17'he1b3:	data_out=16'ha00;
17'he1b4:	data_out=16'h8298;
17'he1b5:	data_out=16'h83ef;
17'he1b6:	data_out=16'h8543;
17'he1b7:	data_out=16'h874f;
17'he1b8:	data_out=16'ha00;
17'he1b9:	data_out=16'ha00;
17'he1ba:	data_out=16'h89fd;
17'he1bb:	data_out=16'h89fd;
17'he1bc:	data_out=16'h87a4;
17'he1bd:	data_out=16'h958;
17'he1be:	data_out=16'h80e5;
17'he1bf:	data_out=16'h9f1;
17'he1c0:	data_out=16'h8990;
17'he1c1:	data_out=16'h11;
17'he1c2:	data_out=16'h8a00;
17'he1c3:	data_out=16'h337;
17'he1c4:	data_out=16'h801d;
17'he1c5:	data_out=16'h86c6;
17'he1c6:	data_out=16'h88b2;
17'he1c7:	data_out=16'h89fb;
17'he1c8:	data_out=16'h3ec;
17'he1c9:	data_out=16'h8a00;
17'he1ca:	data_out=16'h87e1;
17'he1cb:	data_out=16'h8a00;
17'he1cc:	data_out=16'h8a00;
17'he1cd:	data_out=16'h3c5;
17'he1ce:	data_out=16'h89e3;
17'he1cf:	data_out=16'h8a00;
17'he1d0:	data_out=16'h880b;
17'he1d1:	data_out=16'h89ff;
17'he1d2:	data_out=16'h8a00;
17'he1d3:	data_out=16'ha00;
17'he1d4:	data_out=16'ha00;
17'he1d5:	data_out=16'h8a00;
17'he1d6:	data_out=16'h8a00;
17'he1d7:	data_out=16'h89fd;
17'he1d8:	data_out=16'h86d4;
17'he1d9:	data_out=16'h8956;
17'he1da:	data_out=16'h9f7;
17'he1db:	data_out=16'h842;
17'he1dc:	data_out=16'h9f2;
17'he1dd:	data_out=16'h89f9;
17'he1de:	data_out=16'h9fd;
17'he1df:	data_out=16'h2c6;
17'he1e0:	data_out=16'h8a00;
17'he1e1:	data_out=16'hb9;
17'he1e2:	data_out=16'h48d;
17'he1e3:	data_out=16'ha00;
17'he1e4:	data_out=16'ha00;
17'he1e5:	data_out=16'h8335;
17'he1e6:	data_out=16'h82c;
17'he1e7:	data_out=16'h89a7;
17'he1e8:	data_out=16'h80f2;
17'he1e9:	data_out=16'h89fb;
17'he1ea:	data_out=16'h810f;
17'he1eb:	data_out=16'h106;
17'he1ec:	data_out=16'h89f9;
17'he1ed:	data_out=16'ha00;
17'he1ee:	data_out=16'h8110;
17'he1ef:	data_out=16'h8a00;
17'he1f0:	data_out=16'h810b;
17'he1f1:	data_out=16'h892c;
17'he1f2:	data_out=16'h89f5;
17'he1f3:	data_out=16'h82cf;
17'he1f4:	data_out=16'h8a00;
17'he1f5:	data_out=16'hed;
17'he1f6:	data_out=16'h6c7;
17'he1f7:	data_out=16'h8a00;
17'he1f8:	data_out=16'h18;
17'he1f9:	data_out=16'h89fc;
17'he1fa:	data_out=16'h9fd;
17'he1fb:	data_out=16'h80e6;
17'he1fc:	data_out=16'h384;
17'he1fd:	data_out=16'h9e4;
17'he1fe:	data_out=16'h89ff;
17'he1ff:	data_out=16'h879f;
17'he200:	data_out=16'h395;
17'he201:	data_out=16'h661;
17'he202:	data_out=16'h8a00;
17'he203:	data_out=16'h84da;
17'he204:	data_out=16'h88bc;
17'he205:	data_out=16'h8a00;
17'he206:	data_out=16'h2f9;
17'he207:	data_out=16'h89f1;
17'he208:	data_out=16'h18b;
17'he209:	data_out=16'h56f;
17'he20a:	data_out=16'h89f8;
17'he20b:	data_out=16'h9ff;
17'he20c:	data_out=16'h89f0;
17'he20d:	data_out=16'h8a00;
17'he20e:	data_out=16'h871e;
17'he20f:	data_out=16'h89fc;
17'he210:	data_out=16'h9f0;
17'he211:	data_out=16'h66d;
17'he212:	data_out=16'h9f7;
17'he213:	data_out=16'h834d;
17'he214:	data_out=16'h9f8;
17'he215:	data_out=16'h8a00;
17'he216:	data_out=16'h8a00;
17'he217:	data_out=16'h9f5;
17'he218:	data_out=16'h80d9;
17'he219:	data_out=16'ha00;
17'he21a:	data_out=16'h8a00;
17'he21b:	data_out=16'h9f9;
17'he21c:	data_out=16'h9e5;
17'he21d:	data_out=16'h9fe;
17'he21e:	data_out=16'h9ee;
17'he21f:	data_out=16'h9ec;
17'he220:	data_out=16'ha00;
17'he221:	data_out=16'h8709;
17'he222:	data_out=16'h89d6;
17'he223:	data_out=16'h89f6;
17'he224:	data_out=16'h89ef;
17'he225:	data_out=16'h86a7;
17'he226:	data_out=16'h89ff;
17'he227:	data_out=16'ha00;
17'he228:	data_out=16'h869e;
17'he229:	data_out=16'h8a00;
17'he22a:	data_out=16'h89f8;
17'he22b:	data_out=16'ha00;
17'he22c:	data_out=16'h8a00;
17'he22d:	data_out=16'h89ed;
17'he22e:	data_out=16'h8356;
17'he22f:	data_out=16'h9fd;
17'he230:	data_out=16'h8a00;
17'he231:	data_out=16'h275;
17'he232:	data_out=16'h8a00;
17'he233:	data_out=16'ha00;
17'he234:	data_out=16'h564;
17'he235:	data_out=16'h12d;
17'he236:	data_out=16'ha00;
17'he237:	data_out=16'h85ff;
17'he238:	data_out=16'ha00;
17'he239:	data_out=16'ha00;
17'he23a:	data_out=16'h58b;
17'he23b:	data_out=16'h89f0;
17'he23c:	data_out=16'h470;
17'he23d:	data_out=16'h6db;
17'he23e:	data_out=16'h869d;
17'he23f:	data_out=16'h8a00;
17'he240:	data_out=16'h8a00;
17'he241:	data_out=16'h9ef;
17'he242:	data_out=16'h8a00;
17'he243:	data_out=16'h8672;
17'he244:	data_out=16'ha00;
17'he245:	data_out=16'h8a00;
17'he246:	data_out=16'h89b1;
17'he247:	data_out=16'h8586;
17'he248:	data_out=16'h6e1;
17'he249:	data_out=16'h8578;
17'he24a:	data_out=16'h8560;
17'he24b:	data_out=16'h89f3;
17'he24c:	data_out=16'h8a00;
17'he24d:	data_out=16'h8639;
17'he24e:	data_out=16'h86b9;
17'he24f:	data_out=16'h8a00;
17'he250:	data_out=16'h8a00;
17'he251:	data_out=16'h123;
17'he252:	data_out=16'h89fe;
17'he253:	data_out=16'ha00;
17'he254:	data_out=16'ha00;
17'he255:	data_out=16'h8016;
17'he256:	data_out=16'h89f5;
17'he257:	data_out=16'h89ff;
17'he258:	data_out=16'h832e;
17'he259:	data_out=16'h89ff;
17'he25a:	data_out=16'h9fd;
17'he25b:	data_out=16'ha00;
17'he25c:	data_out=16'h9e9;
17'he25d:	data_out=16'h89fc;
17'he25e:	data_out=16'h9e4;
17'he25f:	data_out=16'h303;
17'he260:	data_out=16'h8a00;
17'he261:	data_out=16'h8046;
17'he262:	data_out=16'h9ff;
17'he263:	data_out=16'ha00;
17'he264:	data_out=16'ha00;
17'he265:	data_out=16'h8e8;
17'he266:	data_out=16'ha00;
17'he267:	data_out=16'h89f0;
17'he268:	data_out=16'h86db;
17'he269:	data_out=16'h818e;
17'he26a:	data_out=16'h872d;
17'he26b:	data_out=16'h89c2;
17'he26c:	data_out=16'h89f4;
17'he26d:	data_out=16'ha00;
17'he26e:	data_out=16'h872e;
17'he26f:	data_out=16'h8a00;
17'he270:	data_out=16'h8727;
17'he271:	data_out=16'h81de;
17'he272:	data_out=16'h8a00;
17'he273:	data_out=16'h8a00;
17'he274:	data_out=16'h8a00;
17'he275:	data_out=16'h8a00;
17'he276:	data_out=16'h9ff;
17'he277:	data_out=16'h8a00;
17'he278:	data_out=16'h8a00;
17'he279:	data_out=16'h89d4;
17'he27a:	data_out=16'h9fd;
17'he27b:	data_out=16'h869f;
17'he27c:	data_out=16'h4f8;
17'he27d:	data_out=16'h1a0;
17'he27e:	data_out=16'h9fb;
17'he27f:	data_out=16'h89ff;
17'he280:	data_out=16'h89f5;
17'he281:	data_out=16'h8a00;
17'he282:	data_out=16'h8a00;
17'he283:	data_out=16'h89fd;
17'he284:	data_out=16'h891e;
17'he285:	data_out=16'h8a00;
17'he286:	data_out=16'h9fd;
17'he287:	data_out=16'h9ff;
17'he288:	data_out=16'h5ff;
17'he289:	data_out=16'ha00;
17'he28a:	data_out=16'h89fd;
17'he28b:	data_out=16'ha00;
17'he28c:	data_out=16'h9ff;
17'he28d:	data_out=16'h8a00;
17'he28e:	data_out=16'h8a00;
17'he28f:	data_out=16'h8a00;
17'he290:	data_out=16'h9a3;
17'he291:	data_out=16'h8779;
17'he292:	data_out=16'h8a2;
17'he293:	data_out=16'ha00;
17'he294:	data_out=16'h808a;
17'he295:	data_out=16'h8a00;
17'he296:	data_out=16'h8a00;
17'he297:	data_out=16'h6b6;
17'he298:	data_out=16'h8a00;
17'he299:	data_out=16'ha00;
17'he29a:	data_out=16'h8a00;
17'he29b:	data_out=16'h81c3;
17'he29c:	data_out=16'h8a00;
17'he29d:	data_out=16'h177;
17'he29e:	data_out=16'h89fc;
17'he29f:	data_out=16'h960;
17'he2a0:	data_out=16'h89fe;
17'he2a1:	data_out=16'h8a00;
17'he2a2:	data_out=16'h8967;
17'he2a3:	data_out=16'h9fe;
17'he2a4:	data_out=16'h9ff;
17'he2a5:	data_out=16'h56e;
17'he2a6:	data_out=16'h9ee;
17'he2a7:	data_out=16'h9fa;
17'he2a8:	data_out=16'h8a00;
17'he2a9:	data_out=16'h8a00;
17'he2aa:	data_out=16'h851e;
17'he2ab:	data_out=16'ha00;
17'he2ac:	data_out=16'h8a00;
17'he2ad:	data_out=16'ha00;
17'he2ae:	data_out=16'h13e;
17'he2af:	data_out=16'h89ff;
17'he2b0:	data_out=16'h8a00;
17'he2b1:	data_out=16'h89fb;
17'he2b2:	data_out=16'h8a00;
17'he2b3:	data_out=16'h495;
17'he2b4:	data_out=16'h89e8;
17'he2b5:	data_out=16'h88ae;
17'he2b6:	data_out=16'h8667;
17'he2b7:	data_out=16'h8a00;
17'he2b8:	data_out=16'h870e;
17'he2b9:	data_out=16'h85fe;
17'he2ba:	data_out=16'ha00;
17'he2bb:	data_out=16'h851f;
17'he2bc:	data_out=16'h8a00;
17'he2bd:	data_out=16'h89ff;
17'he2be:	data_out=16'h8a00;
17'he2bf:	data_out=16'h8a00;
17'he2c0:	data_out=16'h8a00;
17'he2c1:	data_out=16'h8a00;
17'he2c2:	data_out=16'h9fe;
17'he2c3:	data_out=16'h89fe;
17'he2c4:	data_out=16'h8908;
17'he2c5:	data_out=16'h8a00;
17'he2c6:	data_out=16'h8a00;
17'he2c7:	data_out=16'ha00;
17'he2c8:	data_out=16'ha00;
17'he2c9:	data_out=16'h369;
17'he2ca:	data_out=16'h9fe;
17'he2cb:	data_out=16'ha00;
17'he2cc:	data_out=16'h812b;
17'he2cd:	data_out=16'h88ab;
17'he2ce:	data_out=16'h5f;
17'he2cf:	data_out=16'h804;
17'he2d0:	data_out=16'h8a00;
17'he2d1:	data_out=16'h8a00;
17'he2d2:	data_out=16'h9fc;
17'he2d3:	data_out=16'h8f6;
17'he2d4:	data_out=16'h89f4;
17'he2d5:	data_out=16'h5cf;
17'he2d6:	data_out=16'h89fe;
17'he2d7:	data_out=16'h89fe;
17'he2d8:	data_out=16'h8a00;
17'he2d9:	data_out=16'h8a00;
17'he2da:	data_out=16'h9e1;
17'he2db:	data_out=16'h883f;
17'he2dc:	data_out=16'h8a00;
17'he2dd:	data_out=16'h8a00;
17'he2de:	data_out=16'h89ff;
17'he2df:	data_out=16'h89fd;
17'he2e0:	data_out=16'h9fe;
17'he2e1:	data_out=16'h8a00;
17'he2e2:	data_out=16'ha00;
17'he2e3:	data_out=16'h69b;
17'he2e4:	data_out=16'ha00;
17'he2e5:	data_out=16'h9fb;
17'he2e6:	data_out=16'ha00;
17'he2e7:	data_out=16'h89f5;
17'he2e8:	data_out=16'h8a00;
17'he2e9:	data_out=16'h9dc;
17'he2ea:	data_out=16'h8a00;
17'he2eb:	data_out=16'h8a00;
17'he2ec:	data_out=16'h8a00;
17'he2ed:	data_out=16'h5ce;
17'he2ee:	data_out=16'h8a00;
17'he2ef:	data_out=16'h8a00;
17'he2f0:	data_out=16'h8a00;
17'he2f1:	data_out=16'h89f7;
17'he2f2:	data_out=16'h8a00;
17'he2f3:	data_out=16'h8a00;
17'he2f4:	data_out=16'h8a00;
17'he2f5:	data_out=16'h8a00;
17'he2f6:	data_out=16'h9f0;
17'he2f7:	data_out=16'h89f0;
17'he2f8:	data_out=16'h8a00;
17'he2f9:	data_out=16'h8a00;
17'he2fa:	data_out=16'h801e;
17'he2fb:	data_out=16'h8a00;
17'he2fc:	data_out=16'h8a00;
17'he2fd:	data_out=16'h813b;
17'he2fe:	data_out=16'h9f8;
17'he2ff:	data_out=16'h8a00;
17'he300:	data_out=16'h89fc;
17'he301:	data_out=16'h8a00;
17'he302:	data_out=16'h8a00;
17'he303:	data_out=16'h89ff;
17'he304:	data_out=16'h88ea;
17'he305:	data_out=16'h8a00;
17'he306:	data_out=16'h9ff;
17'he307:	data_out=16'ha00;
17'he308:	data_out=16'h8a00;
17'he309:	data_out=16'ha00;
17'he30a:	data_out=16'h89f0;
17'he30b:	data_out=16'ha00;
17'he30c:	data_out=16'ha00;
17'he30d:	data_out=16'h8a00;
17'he30e:	data_out=16'h8a00;
17'he30f:	data_out=16'h89fa;
17'he310:	data_out=16'h961;
17'he311:	data_out=16'h89d3;
17'he312:	data_out=16'h50b;
17'he313:	data_out=16'h9f8;
17'he314:	data_out=16'h853d;
17'he315:	data_out=16'h8a00;
17'he316:	data_out=16'h8a00;
17'he317:	data_out=16'h862b;
17'he318:	data_out=16'h8a00;
17'he319:	data_out=16'h9c0;
17'he31a:	data_out=16'h8a00;
17'he31b:	data_out=16'h89ec;
17'he31c:	data_out=16'h8a00;
17'he31d:	data_out=16'h89e5;
17'he31e:	data_out=16'h89fd;
17'he31f:	data_out=16'h9c7;
17'he320:	data_out=16'h8a00;
17'he321:	data_out=16'h8a00;
17'he322:	data_out=16'h605;
17'he323:	data_out=16'ha00;
17'he324:	data_out=16'ha00;
17'he325:	data_out=16'h8f0;
17'he326:	data_out=16'h9e7;
17'he327:	data_out=16'h88b7;
17'he328:	data_out=16'h8a00;
17'he329:	data_out=16'h8a00;
17'he32a:	data_out=16'h86c6;
17'he32b:	data_out=16'ha00;
17'he32c:	data_out=16'h8a00;
17'he32d:	data_out=16'ha00;
17'he32e:	data_out=16'h472;
17'he32f:	data_out=16'h8a00;
17'he330:	data_out=16'h89f8;
17'he331:	data_out=16'h8a00;
17'he332:	data_out=16'h8a00;
17'he333:	data_out=16'h895d;
17'he334:	data_out=16'h89f8;
17'he335:	data_out=16'h88be;
17'he336:	data_out=16'h89fc;
17'he337:	data_out=16'h8a00;
17'he338:	data_out=16'h89fb;
17'he339:	data_out=16'h89fe;
17'he33a:	data_out=16'ha00;
17'he33b:	data_out=16'h433;
17'he33c:	data_out=16'h8a00;
17'he33d:	data_out=16'h8a00;
17'he33e:	data_out=16'h8a00;
17'he33f:	data_out=16'h8a00;
17'he340:	data_out=16'h8a00;
17'he341:	data_out=16'h8a00;
17'he342:	data_out=16'ha00;
17'he343:	data_out=16'h8a00;
17'he344:	data_out=16'h89d6;
17'he345:	data_out=16'h8a00;
17'he346:	data_out=16'h8a00;
17'he347:	data_out=16'ha00;
17'he348:	data_out=16'ha00;
17'he349:	data_out=16'h91b;
17'he34a:	data_out=16'h9eb;
17'he34b:	data_out=16'ha00;
17'he34c:	data_out=16'h936;
17'he34d:	data_out=16'h6e0;
17'he34e:	data_out=16'h86b5;
17'he34f:	data_out=16'ha00;
17'he350:	data_out=16'h8a00;
17'he351:	data_out=16'h8a00;
17'he352:	data_out=16'ha00;
17'he353:	data_out=16'h89fc;
17'he354:	data_out=16'h89fe;
17'he355:	data_out=16'h91a;
17'he356:	data_out=16'h876;
17'he357:	data_out=16'h8a00;
17'he358:	data_out=16'h8a00;
17'he359:	data_out=16'h89f7;
17'he35a:	data_out=16'h870b;
17'he35b:	data_out=16'h8981;
17'he35c:	data_out=16'h8a00;
17'he35d:	data_out=16'h8a00;
17'he35e:	data_out=16'h8a00;
17'he35f:	data_out=16'h89fc;
17'he360:	data_out=16'h9fd;
17'he361:	data_out=16'h8a00;
17'he362:	data_out=16'h9fb;
17'he363:	data_out=16'h89d7;
17'he364:	data_out=16'ha00;
17'he365:	data_out=16'h9fa;
17'he366:	data_out=16'h9ff;
17'he367:	data_out=16'h81a9;
17'he368:	data_out=16'h8a00;
17'he369:	data_out=16'h88b;
17'he36a:	data_out=16'h8a00;
17'he36b:	data_out=16'h8a00;
17'he36c:	data_out=16'h89fe;
17'he36d:	data_out=16'h89f7;
17'he36e:	data_out=16'h8a00;
17'he36f:	data_out=16'h8a00;
17'he370:	data_out=16'h8a00;
17'he371:	data_out=16'h89ee;
17'he372:	data_out=16'h8a00;
17'he373:	data_out=16'h8a00;
17'he374:	data_out=16'h8a00;
17'he375:	data_out=16'h8a00;
17'he376:	data_out=16'ha00;
17'he377:	data_out=16'h9cc;
17'he378:	data_out=16'h8a00;
17'he379:	data_out=16'h8a00;
17'he37a:	data_out=16'h89ff;
17'he37b:	data_out=16'h8a00;
17'he37c:	data_out=16'h8a00;
17'he37d:	data_out=16'h85d4;
17'he37e:	data_out=16'ha00;
17'he37f:	data_out=16'h8a00;
17'he380:	data_out=16'h8a00;
17'he381:	data_out=16'h8a00;
17'he382:	data_out=16'h89fe;
17'he383:	data_out=16'h89f2;
17'he384:	data_out=16'h89f9;
17'he385:	data_out=16'h8a00;
17'he386:	data_out=16'h9ef;
17'he387:	data_out=16'ha00;
17'he388:	data_out=16'h8a00;
17'he389:	data_out=16'ha00;
17'he38a:	data_out=16'h89d6;
17'he38b:	data_out=16'ha00;
17'he38c:	data_out=16'ha00;
17'he38d:	data_out=16'h8a00;
17'he38e:	data_out=16'h8a00;
17'he38f:	data_out=16'h8976;
17'he390:	data_out=16'h8d7;
17'he391:	data_out=16'h889d;
17'he392:	data_out=16'h84;
17'he393:	data_out=16'h97c;
17'he394:	data_out=16'h8557;
17'he395:	data_out=16'h8a00;
17'he396:	data_out=16'h8a00;
17'he397:	data_out=16'h8510;
17'he398:	data_out=16'h8a00;
17'he399:	data_out=16'ha00;
17'he39a:	data_out=16'h8a00;
17'he39b:	data_out=16'h897c;
17'he39c:	data_out=16'h8a00;
17'he39d:	data_out=16'h89d6;
17'he39e:	data_out=16'h89f6;
17'he39f:	data_out=16'h9d8;
17'he3a0:	data_out=16'h8a00;
17'he3a1:	data_out=16'h8a00;
17'he3a2:	data_out=16'h958;
17'he3a3:	data_out=16'ha00;
17'he3a4:	data_out=16'ha00;
17'he3a5:	data_out=16'h920;
17'he3a6:	data_out=16'h9f8;
17'he3a7:	data_out=16'h89dc;
17'he3a8:	data_out=16'h8a00;
17'he3a9:	data_out=16'h89f5;
17'he3aa:	data_out=16'h847a;
17'he3ab:	data_out=16'ha00;
17'he3ac:	data_out=16'h8a00;
17'he3ad:	data_out=16'ha00;
17'he3ae:	data_out=16'ha00;
17'he3af:	data_out=16'h89ff;
17'he3b0:	data_out=16'h89ae;
17'he3b1:	data_out=16'h8a00;
17'he3b2:	data_out=16'h8a00;
17'he3b3:	data_out=16'h89ed;
17'he3b4:	data_out=16'h89fb;
17'he3b5:	data_out=16'h89d9;
17'he3b6:	data_out=16'h89fd;
17'he3b7:	data_out=16'h89ce;
17'he3b8:	data_out=16'h8a00;
17'he3b9:	data_out=16'h89f3;
17'he3ba:	data_out=16'ha00;
17'he3bb:	data_out=16'h975;
17'he3bc:	data_out=16'h8a00;
17'he3bd:	data_out=16'h8a00;
17'he3be:	data_out=16'h8a00;
17'he3bf:	data_out=16'h8a00;
17'he3c0:	data_out=16'h89ff;
17'he3c1:	data_out=16'h8a00;
17'he3c2:	data_out=16'ha00;
17'he3c3:	data_out=16'h89fd;
17'he3c4:	data_out=16'h89fb;
17'he3c5:	data_out=16'h8a00;
17'he3c6:	data_out=16'h8a00;
17'he3c7:	data_out=16'ha00;
17'he3c8:	data_out=16'h9e5;
17'he3c9:	data_out=16'h912;
17'he3ca:	data_out=16'h573;
17'he3cb:	data_out=16'ha00;
17'he3cc:	data_out=16'h9c1;
17'he3cd:	data_out=16'h983;
17'he3ce:	data_out=16'h89ef;
17'he3cf:	data_out=16'ha00;
17'he3d0:	data_out=16'h89f9;
17'he3d1:	data_out=16'h8a00;
17'he3d2:	data_out=16'ha00;
17'he3d3:	data_out=16'h89f6;
17'he3d4:	data_out=16'h8a00;
17'he3d5:	data_out=16'h9cf;
17'he3d6:	data_out=16'h8013;
17'he3d7:	data_out=16'h89fe;
17'he3d8:	data_out=16'h8a00;
17'he3d9:	data_out=16'h89fd;
17'he3da:	data_out=16'h89af;
17'he3db:	data_out=16'h89cf;
17'he3dc:	data_out=16'h8a00;
17'he3dd:	data_out=16'h8a00;
17'he3de:	data_out=16'h89fd;
17'he3df:	data_out=16'h89f9;
17'he3e0:	data_out=16'h9fb;
17'he3e1:	data_out=16'h8a00;
17'he3e2:	data_out=16'ha00;
17'he3e3:	data_out=16'h89ee;
17'he3e4:	data_out=16'h446;
17'he3e5:	data_out=16'h9cb;
17'he3e6:	data_out=16'ha00;
17'he3e7:	data_out=16'ha00;
17'he3e8:	data_out=16'h8a00;
17'he3e9:	data_out=16'h89eb;
17'he3ea:	data_out=16'h8a00;
17'he3eb:	data_out=16'h8a00;
17'he3ec:	data_out=16'h8a00;
17'he3ed:	data_out=16'h89ee;
17'he3ee:	data_out=16'h8a00;
17'he3ef:	data_out=16'h89ff;
17'he3f0:	data_out=16'h8a00;
17'he3f1:	data_out=16'h8986;
17'he3f2:	data_out=16'h8a00;
17'he3f3:	data_out=16'h8a00;
17'he3f4:	data_out=16'h89e9;
17'he3f5:	data_out=16'h8a00;
17'he3f6:	data_out=16'ha00;
17'he3f7:	data_out=16'h9db;
17'he3f8:	data_out=16'h8a00;
17'he3f9:	data_out=16'h8a00;
17'he3fa:	data_out=16'h89d9;
17'he3fb:	data_out=16'h8a00;
17'he3fc:	data_out=16'h8a00;
17'he3fd:	data_out=16'h88ef;
17'he3fe:	data_out=16'ha00;
17'he3ff:	data_out=16'h8a00;
17'he400:	data_out=16'h8a00;
17'he401:	data_out=16'h89df;
17'he402:	data_out=16'h89c3;
17'he403:	data_out=16'h851b;
17'he404:	data_out=16'h89e5;
17'he405:	data_out=16'h8a00;
17'he406:	data_out=16'h9f9;
17'he407:	data_out=16'h9e1;
17'he408:	data_out=16'h89f7;
17'he409:	data_out=16'ha00;
17'he40a:	data_out=16'h86b9;
17'he40b:	data_out=16'ha00;
17'he40c:	data_out=16'h9e8;
17'he40d:	data_out=16'h89fc;
17'he40e:	data_out=16'h89af;
17'he40f:	data_out=16'h8372;
17'he410:	data_out=16'h9b8;
17'he411:	data_out=16'h8739;
17'he412:	data_out=16'h8603;
17'he413:	data_out=16'h9d5;
17'he414:	data_out=16'h849e;
17'he415:	data_out=16'h8a00;
17'he416:	data_out=16'h89f8;
17'he417:	data_out=16'h830c;
17'he418:	data_out=16'h8a00;
17'he419:	data_out=16'ha00;
17'he41a:	data_out=16'h8a00;
17'he41b:	data_out=16'h86a4;
17'he41c:	data_out=16'h89f7;
17'he41d:	data_out=16'h89b6;
17'he41e:	data_out=16'h88d8;
17'he41f:	data_out=16'h9eb;
17'he420:	data_out=16'h89f6;
17'he421:	data_out=16'h89a3;
17'he422:	data_out=16'h9f7;
17'he423:	data_out=16'h9f8;
17'he424:	data_out=16'h9f8;
17'he425:	data_out=16'h9e7;
17'he426:	data_out=16'h9fa;
17'he427:	data_out=16'h89d6;
17'he428:	data_out=16'h8991;
17'he429:	data_out=16'h9d5;
17'he42a:	data_out=16'h351;
17'he42b:	data_out=16'h9fd;
17'he42c:	data_out=16'h89fa;
17'he42d:	data_out=16'ha00;
17'he42e:	data_out=16'ha00;
17'he42f:	data_out=16'h89cc;
17'he430:	data_out=16'h8711;
17'he431:	data_out=16'h89ca;
17'he432:	data_out=16'h89d5;
17'he433:	data_out=16'h899f;
17'he434:	data_out=16'h89e0;
17'he435:	data_out=16'h8951;
17'he436:	data_out=16'h89d2;
17'he437:	data_out=16'h84f9;
17'he438:	data_out=16'h89f0;
17'he439:	data_out=16'h89c9;
17'he43a:	data_out=16'h9fb;
17'he43b:	data_out=16'ha00;
17'he43c:	data_out=16'h89cd;
17'he43d:	data_out=16'h89e8;
17'he43e:	data_out=16'h8992;
17'he43f:	data_out=16'h8a00;
17'he440:	data_out=16'h89fd;
17'he441:	data_out=16'h89f8;
17'he442:	data_out=16'h9fa;
17'he443:	data_out=16'h93;
17'he444:	data_out=16'h8870;
17'he445:	data_out=16'h8a00;
17'he446:	data_out=16'h8a00;
17'he447:	data_out=16'ha00;
17'he448:	data_out=16'h9f1;
17'he449:	data_out=16'h9f1;
17'he44a:	data_out=16'h89d8;
17'he44b:	data_out=16'ha00;
17'he44c:	data_out=16'h9fa;
17'he44d:	data_out=16'ha00;
17'he44e:	data_out=16'h894c;
17'he44f:	data_out=16'ha00;
17'he450:	data_out=16'h8941;
17'he451:	data_out=16'h89c9;
17'he452:	data_out=16'ha00;
17'he453:	data_out=16'h899e;
17'he454:	data_out=16'h89d2;
17'he455:	data_out=16'ha00;
17'he456:	data_out=16'h8889;
17'he457:	data_out=16'h6df;
17'he458:	data_out=16'h89fb;
17'he459:	data_out=16'h89ed;
17'he45a:	data_out=16'h896d;
17'he45b:	data_out=16'h89b0;
17'he45c:	data_out=16'h8a00;
17'he45d:	data_out=16'h89dd;
17'he45e:	data_out=16'h89bf;
17'he45f:	data_out=16'h89ed;
17'he460:	data_out=16'h9f4;
17'he461:	data_out=16'h89c5;
17'he462:	data_out=16'ha00;
17'he463:	data_out=16'h8977;
17'he464:	data_out=16'h89f8;
17'he465:	data_out=16'h813;
17'he466:	data_out=16'ha00;
17'he467:	data_out=16'ha00;
17'he468:	data_out=16'h8993;
17'he469:	data_out=16'h89e4;
17'he46a:	data_out=16'h89a9;
17'he46b:	data_out=16'h89ff;
17'he46c:	data_out=16'h8a00;
17'he46d:	data_out=16'h898b;
17'he46e:	data_out=16'h89a9;
17'he46f:	data_out=16'h89f7;
17'he470:	data_out=16'h89ae;
17'he471:	data_out=16'h87e1;
17'he472:	data_out=16'h89ff;
17'he473:	data_out=16'h89e8;
17'he474:	data_out=16'h87c3;
17'he475:	data_out=16'h8a00;
17'he476:	data_out=16'ha00;
17'he477:	data_out=16'h9fa;
17'he478:	data_out=16'h8a00;
17'he479:	data_out=16'h8a00;
17'he47a:	data_out=16'h881b;
17'he47b:	data_out=16'h8991;
17'he47c:	data_out=16'h8a00;
17'he47d:	data_out=16'h8497;
17'he47e:	data_out=16'ha00;
17'he47f:	data_out=16'h8a00;
17'he480:	data_out=16'h8a00;
17'he481:	data_out=16'h89bd;
17'he482:	data_out=16'h89d9;
17'he483:	data_out=16'h859f;
17'he484:	data_out=16'h89c7;
17'he485:	data_out=16'h890d;
17'he486:	data_out=16'ha00;
17'he487:	data_out=16'h9ef;
17'he488:	data_out=16'h89f4;
17'he489:	data_out=16'ha00;
17'he48a:	data_out=16'h83b3;
17'he48b:	data_out=16'ha00;
17'he48c:	data_out=16'h9f3;
17'he48d:	data_out=16'h89ff;
17'he48e:	data_out=16'h8952;
17'he48f:	data_out=16'h8871;
17'he490:	data_out=16'h9f5;
17'he491:	data_out=16'h1bf;
17'he492:	data_out=16'h89fe;
17'he493:	data_out=16'h88d8;
17'he494:	data_out=16'h881c;
17'he495:	data_out=16'h89f9;
17'he496:	data_out=16'h894d;
17'he497:	data_out=16'h86e4;
17'he498:	data_out=16'h8a00;
17'he499:	data_out=16'h9f6;
17'he49a:	data_out=16'h895a;
17'he49b:	data_out=16'h8941;
17'he49c:	data_out=16'h89db;
17'he49d:	data_out=16'h89b2;
17'he49e:	data_out=16'h88d9;
17'he49f:	data_out=16'h9e8;
17'he4a0:	data_out=16'h89e0;
17'he4a1:	data_out=16'h893e;
17'he4a2:	data_out=16'ha00;
17'he4a3:	data_out=16'h9f1;
17'he4a4:	data_out=16'h9f1;
17'he4a5:	data_out=16'h9ee;
17'he4a6:	data_out=16'h9c1;
17'he4a7:	data_out=16'h89b2;
17'he4a8:	data_out=16'h892c;
17'he4a9:	data_out=16'h9d5;
17'he4aa:	data_out=16'h8143;
17'he4ab:	data_out=16'h9fb;
17'he4ac:	data_out=16'h8963;
17'he4ad:	data_out=16'ha00;
17'he4ae:	data_out=16'h6a4;
17'he4af:	data_out=16'h899c;
17'he4b0:	data_out=16'h813a;
17'he4b1:	data_out=16'h89;
17'he4b2:	data_out=16'h81d2;
17'he4b3:	data_out=16'h89b4;
17'he4b4:	data_out=16'h89ef;
17'he4b5:	data_out=16'h86c7;
17'he4b6:	data_out=16'h89ca;
17'he4b7:	data_out=16'h8999;
17'he4b8:	data_out=16'h89f9;
17'he4b9:	data_out=16'h89df;
17'he4ba:	data_out=16'ha00;
17'he4bb:	data_out=16'ha00;
17'he4bc:	data_out=16'h89c7;
17'he4bd:	data_out=16'h89d4;
17'he4be:	data_out=16'h892d;
17'he4bf:	data_out=16'h891b;
17'he4c0:	data_out=16'h894f;
17'he4c1:	data_out=16'h89d2;
17'he4c2:	data_out=16'ha00;
17'he4c3:	data_out=16'h9f3;
17'he4c4:	data_out=16'h3ca;
17'he4c5:	data_out=16'h89f8;
17'he4c6:	data_out=16'h8a00;
17'he4c7:	data_out=16'h9c8;
17'he4c8:	data_out=16'h9fb;
17'he4c9:	data_out=16'h9f1;
17'he4ca:	data_out=16'h89aa;
17'he4cb:	data_out=16'ha00;
17'he4cc:	data_out=16'h9f4;
17'he4cd:	data_out=16'ha00;
17'he4ce:	data_out=16'h8a00;
17'he4cf:	data_out=16'ha00;
17'he4d0:	data_out=16'h80ba;
17'he4d1:	data_out=16'h89ec;
17'he4d2:	data_out=16'h9fe;
17'he4d3:	data_out=16'h8975;
17'he4d4:	data_out=16'h89ce;
17'he4d5:	data_out=16'h9fa;
17'he4d6:	data_out=16'h89f8;
17'he4d7:	data_out=16'h8ab;
17'he4d8:	data_out=16'h89fc;
17'he4d9:	data_out=16'h839b;
17'he4da:	data_out=16'h89de;
17'he4db:	data_out=16'h893d;
17'he4dc:	data_out=16'h89c6;
17'he4dd:	data_out=16'h89a0;
17'he4de:	data_out=16'h88f7;
17'he4df:	data_out=16'h89f4;
17'he4e0:	data_out=16'h9e8;
17'he4e1:	data_out=16'h836b;
17'he4e2:	data_out=16'h4fa;
17'he4e3:	data_out=16'h89ab;
17'he4e4:	data_out=16'h8a00;
17'he4e5:	data_out=16'h9ed;
17'he4e6:	data_out=16'ha00;
17'he4e7:	data_out=16'ha00;
17'he4e8:	data_out=16'h8919;
17'he4e9:	data_out=16'h89fd;
17'he4ea:	data_out=16'h8944;
17'he4eb:	data_out=16'h897a;
17'he4ec:	data_out=16'h8a00;
17'he4ed:	data_out=16'h89b0;
17'he4ee:	data_out=16'h8944;
17'he4ef:	data_out=16'h81a1;
17'he4f0:	data_out=16'h894e;
17'he4f1:	data_out=16'h89b9;
17'he4f2:	data_out=16'h8592;
17'he4f3:	data_out=16'h846c;
17'he4f4:	data_out=16'h81cd;
17'he4f5:	data_out=16'h898a;
17'he4f6:	data_out=16'ha00;
17'he4f7:	data_out=16'h9fd;
17'he4f8:	data_out=16'h475;
17'he4f9:	data_out=16'h8a00;
17'he4fa:	data_out=16'h8929;
17'he4fb:	data_out=16'h892d;
17'he4fc:	data_out=16'h8a00;
17'he4fd:	data_out=16'h8552;
17'he4fe:	data_out=16'ha00;
17'he4ff:	data_out=16'h8a00;
17'he500:	data_out=16'h8a00;
17'he501:	data_out=16'h8a00;
17'he502:	data_out=16'h8a00;
17'he503:	data_out=16'h87c5;
17'he504:	data_out=16'h8994;
17'he505:	data_out=16'h88b5;
17'he506:	data_out=16'ha00;
17'he507:	data_out=16'h9ee;
17'he508:	data_out=16'h8a00;
17'he509:	data_out=16'ha00;
17'he50a:	data_out=16'h8801;
17'he50b:	data_out=16'h951;
17'he50c:	data_out=16'h9fb;
17'he50d:	data_out=16'h8a00;
17'he50e:	data_out=16'h89f8;
17'he50f:	data_out=16'h89d3;
17'he510:	data_out=16'ha00;
17'he511:	data_out=16'h8b5;
17'he512:	data_out=16'h8a00;
17'he513:	data_out=16'h89fe;
17'he514:	data_out=16'h89c8;
17'he515:	data_out=16'h89fd;
17'he516:	data_out=16'h8945;
17'he517:	data_out=16'h898f;
17'he518:	data_out=16'h8a00;
17'he519:	data_out=16'h9f3;
17'he51a:	data_out=16'h894d;
17'he51b:	data_out=16'h89eb;
17'he51c:	data_out=16'h8a00;
17'he51d:	data_out=16'h89d0;
17'he51e:	data_out=16'h89e2;
17'he51f:	data_out=16'h896a;
17'he520:	data_out=16'h89fa;
17'he521:	data_out=16'h89f7;
17'he522:	data_out=16'ha00;
17'he523:	data_out=16'ha00;
17'he524:	data_out=16'ha00;
17'he525:	data_out=16'ha00;
17'he526:	data_out=16'h87f0;
17'he527:	data_out=16'h89e6;
17'he528:	data_out=16'h89f6;
17'he529:	data_out=16'h9c6;
17'he52a:	data_out=16'h8908;
17'he52b:	data_out=16'h8726;
17'he52c:	data_out=16'h8930;
17'he52d:	data_out=16'ha00;
17'he52e:	data_out=16'h87e0;
17'he52f:	data_out=16'h89da;
17'he530:	data_out=16'h822a;
17'he531:	data_out=16'h18d;
17'he532:	data_out=16'h833d;
17'he533:	data_out=16'h89fd;
17'he534:	data_out=16'h8a00;
17'he535:	data_out=16'h892b;
17'he536:	data_out=16'h8a00;
17'he537:	data_out=16'h89fc;
17'he538:	data_out=16'h8a00;
17'he539:	data_out=16'h89fe;
17'he53a:	data_out=16'ha00;
17'he53b:	data_out=16'ha00;
17'he53c:	data_out=16'h8a00;
17'he53d:	data_out=16'h89ee;
17'he53e:	data_out=16'h89f6;
17'he53f:	data_out=16'h88c9;
17'he540:	data_out=16'h8783;
17'he541:	data_out=16'h8a00;
17'he542:	data_out=16'ha00;
17'he543:	data_out=16'ha00;
17'he544:	data_out=16'h77;
17'he545:	data_out=16'h89fd;
17'he546:	data_out=16'h8a00;
17'he547:	data_out=16'h82f6;
17'he548:	data_out=16'h8983;
17'he549:	data_out=16'ha00;
17'he54a:	data_out=16'h89cd;
17'he54b:	data_out=16'ha00;
17'he54c:	data_out=16'h9f9;
17'he54d:	data_out=16'ha00;
17'he54e:	data_out=16'h8a00;
17'he54f:	data_out=16'ha00;
17'he550:	data_out=16'h169;
17'he551:	data_out=16'h89ff;
17'he552:	data_out=16'ha00;
17'he553:	data_out=16'h89d2;
17'he554:	data_out=16'h89fd;
17'he555:	data_out=16'h89b6;
17'he556:	data_out=16'h8a00;
17'he557:	data_out=16'h89f9;
17'he558:	data_out=16'h8a00;
17'he559:	data_out=16'h9b;
17'he55a:	data_out=16'h8a00;
17'he55b:	data_out=16'h89b4;
17'he55c:	data_out=16'h8a00;
17'he55d:	data_out=16'h898d;
17'he55e:	data_out=16'h88d2;
17'he55f:	data_out=16'h89fe;
17'he560:	data_out=16'h9f2;
17'he561:	data_out=16'h849d;
17'he562:	data_out=16'h8803;
17'he563:	data_out=16'h89fd;
17'he564:	data_out=16'h8a00;
17'he565:	data_out=16'ha00;
17'he566:	data_out=16'ha00;
17'he567:	data_out=16'ha00;
17'he568:	data_out=16'h89f6;
17'he569:	data_out=16'h8a00;
17'he56a:	data_out=16'h89f9;
17'he56b:	data_out=16'h88ac;
17'he56c:	data_out=16'h8a00;
17'he56d:	data_out=16'h89ff;
17'he56e:	data_out=16'h89f9;
17'he56f:	data_out=16'h8613;
17'he570:	data_out=16'h89f8;
17'he571:	data_out=16'h89ff;
17'he572:	data_out=16'h8203;
17'he573:	data_out=16'h87e1;
17'he574:	data_out=16'h834a;
17'he575:	data_out=16'h899e;
17'he576:	data_out=16'ha00;
17'he577:	data_out=16'h80c9;
17'he578:	data_out=16'h9f2;
17'he579:	data_out=16'h8a00;
17'he57a:	data_out=16'h89e3;
17'he57b:	data_out=16'h89f6;
17'he57c:	data_out=16'h8a00;
17'he57d:	data_out=16'h8968;
17'he57e:	data_out=16'ha00;
17'he57f:	data_out=16'h89fb;
17'he580:	data_out=16'h8a00;
17'he581:	data_out=16'h8a00;
17'he582:	data_out=16'h8a00;
17'he583:	data_out=16'h8911;
17'he584:	data_out=16'h813a;
17'he585:	data_out=16'h9d1;
17'he586:	data_out=16'ha00;
17'he587:	data_out=16'h898f;
17'he588:	data_out=16'h8a00;
17'he589:	data_out=16'ha00;
17'he58a:	data_out=16'h8a00;
17'he58b:	data_out=16'h8900;
17'he58c:	data_out=16'h898b;
17'he58d:	data_out=16'h8a00;
17'he58e:	data_out=16'h9f5;
17'he58f:	data_out=16'h8a00;
17'he590:	data_out=16'ha00;
17'he591:	data_out=16'h9d8;
17'he592:	data_out=16'h8a00;
17'he593:	data_out=16'h89ff;
17'he594:	data_out=16'h8a00;
17'he595:	data_out=16'h89fc;
17'he596:	data_out=16'h89e8;
17'he597:	data_out=16'h8a00;
17'he598:	data_out=16'h8a00;
17'he599:	data_out=16'h9b5;
17'he59a:	data_out=16'h9d7;
17'he59b:	data_out=16'h8a00;
17'he59c:	data_out=16'h8a00;
17'he59d:	data_out=16'h8a00;
17'he59e:	data_out=16'h89ff;
17'he59f:	data_out=16'h88d7;
17'he5a0:	data_out=16'h89f4;
17'he5a1:	data_out=16'h9f9;
17'he5a2:	data_out=16'ha00;
17'he5a3:	data_out=16'ha00;
17'he5a4:	data_out=16'ha00;
17'he5a5:	data_out=16'ha00;
17'he5a6:	data_out=16'h8a00;
17'he5a7:	data_out=16'h89fe;
17'he5a8:	data_out=16'h9fb;
17'he5a9:	data_out=16'h61d;
17'he5aa:	data_out=16'h89f1;
17'he5ab:	data_out=16'h89fe;
17'he5ac:	data_out=16'h891c;
17'he5ad:	data_out=16'h9d3;
17'he5ae:	data_out=16'h89aa;
17'he5af:	data_out=16'h8a00;
17'he5b0:	data_out=16'h8299;
17'he5b1:	data_out=16'h85a0;
17'he5b2:	data_out=16'h119;
17'he5b3:	data_out=16'h8a00;
17'he5b4:	data_out=16'h8a00;
17'he5b5:	data_out=16'h89fe;
17'he5b6:	data_out=16'h8a00;
17'he5b7:	data_out=16'h8a00;
17'he5b8:	data_out=16'h89ff;
17'he5b9:	data_out=16'h8a00;
17'he5ba:	data_out=16'h6f7;
17'he5bb:	data_out=16'hd2;
17'he5bc:	data_out=16'h8a00;
17'he5bd:	data_out=16'h89b5;
17'he5be:	data_out=16'h9fb;
17'he5bf:	data_out=16'h9d0;
17'he5c0:	data_out=16'h305;
17'he5c1:	data_out=16'h8a00;
17'he5c2:	data_out=16'ha00;
17'he5c3:	data_out=16'ha00;
17'he5c4:	data_out=16'h88aa;
17'he5c5:	data_out=16'h89fc;
17'he5c6:	data_out=16'h8a00;
17'he5c7:	data_out=16'h89e3;
17'he5c8:	data_out=16'h8973;
17'he5c9:	data_out=16'ha00;
17'he5ca:	data_out=16'h89f3;
17'he5cb:	data_out=16'ha00;
17'he5cc:	data_out=16'ha00;
17'he5cd:	data_out=16'ha00;
17'he5ce:	data_out=16'h8a00;
17'he5cf:	data_out=16'ha00;
17'he5d0:	data_out=16'ha00;
17'he5d1:	data_out=16'h8a00;
17'he5d2:	data_out=16'ha00;
17'he5d3:	data_out=16'h8a00;
17'he5d4:	data_out=16'h89fc;
17'he5d5:	data_out=16'h89f5;
17'he5d6:	data_out=16'h8a00;
17'he5d7:	data_out=16'h919;
17'he5d8:	data_out=16'h8a00;
17'he5d9:	data_out=16'h9ee;
17'he5da:	data_out=16'h8a00;
17'he5db:	data_out=16'h89f9;
17'he5dc:	data_out=16'h8a00;
17'he5dd:	data_out=16'h86f9;
17'he5de:	data_out=16'h878a;
17'he5df:	data_out=16'h89fd;
17'he5e0:	data_out=16'h893c;
17'he5e1:	data_out=16'h9d1;
17'he5e2:	data_out=16'h89d9;
17'he5e3:	data_out=16'h8a00;
17'he5e4:	data_out=16'h8a00;
17'he5e5:	data_out=16'ha00;
17'he5e6:	data_out=16'h88b2;
17'he5e7:	data_out=16'ha00;
17'he5e8:	data_out=16'h9fc;
17'he5e9:	data_out=16'h8a00;
17'he5ea:	data_out=16'h9f2;
17'he5eb:	data_out=16'h405;
17'he5ec:	data_out=16'h8a00;
17'he5ed:	data_out=16'h8a00;
17'he5ee:	data_out=16'h9f2;
17'he5ef:	data_out=16'h31;
17'he5f0:	data_out=16'h9f4;
17'he5f1:	data_out=16'h8a00;
17'he5f2:	data_out=16'h9c5;
17'he5f3:	data_out=16'h994;
17'he5f4:	data_out=16'h8459;
17'he5f5:	data_out=16'h85c6;
17'he5f6:	data_out=16'h86ca;
17'he5f7:	data_out=16'h81e0;
17'he5f8:	data_out=16'h9fd;
17'he5f9:	data_out=16'h8a00;
17'he5fa:	data_out=16'h8a00;
17'he5fb:	data_out=16'h9fb;
17'he5fc:	data_out=16'h8a00;
17'he5fd:	data_out=16'h85c7;
17'he5fe:	data_out=16'ha00;
17'he5ff:	data_out=16'h9f6;
17'he600:	data_out=16'h8a00;
17'he601:	data_out=16'h8a00;
17'he602:	data_out=16'h8a00;
17'he603:	data_out=16'h899d;
17'he604:	data_out=16'h8025;
17'he605:	data_out=16'h9e5;
17'he606:	data_out=16'ha00;
17'he607:	data_out=16'h8a00;
17'he608:	data_out=16'h8a00;
17'he609:	data_out=16'h8716;
17'he60a:	data_out=16'h89fe;
17'he60b:	data_out=16'h89f8;
17'he60c:	data_out=16'h8a00;
17'he60d:	data_out=16'h8a00;
17'he60e:	data_out=16'ha00;
17'he60f:	data_out=16'h89ff;
17'he610:	data_out=16'ha00;
17'he611:	data_out=16'h9fd;
17'he612:	data_out=16'h8a00;
17'he613:	data_out=16'h8a00;
17'he614:	data_out=16'h89f5;
17'he615:	data_out=16'h88dc;
17'he616:	data_out=16'h89fd;
17'he617:	data_out=16'h89fc;
17'he618:	data_out=16'h8a00;
17'he619:	data_out=16'h89a9;
17'he61a:	data_out=16'h9ec;
17'he61b:	data_out=16'h8a00;
17'he61c:	data_out=16'h86b2;
17'he61d:	data_out=16'h8a00;
17'he61e:	data_out=16'h89e1;
17'he61f:	data_out=16'h84e9;
17'he620:	data_out=16'h2b7;
17'he621:	data_out=16'ha00;
17'he622:	data_out=16'ha00;
17'he623:	data_out=16'h89ff;
17'he624:	data_out=16'h89ff;
17'he625:	data_out=16'ha00;
17'he626:	data_out=16'h8a00;
17'he627:	data_out=16'h89ff;
17'he628:	data_out=16'ha00;
17'he629:	data_out=16'h95c;
17'he62a:	data_out=16'h89c2;
17'he62b:	data_out=16'h8a00;
17'he62c:	data_out=16'h87b6;
17'he62d:	data_out=16'h9e0;
17'he62e:	data_out=16'h161;
17'he62f:	data_out=16'h8717;
17'he630:	data_out=16'h8a00;
17'he631:	data_out=16'h8941;
17'he632:	data_out=16'h322;
17'he633:	data_out=16'h89f6;
17'he634:	data_out=16'h8a00;
17'he635:	data_out=16'h89ff;
17'he636:	data_out=16'h8a00;
17'he637:	data_out=16'h8a00;
17'he638:	data_out=16'h9f5;
17'he639:	data_out=16'h89fb;
17'he63a:	data_out=16'h8889;
17'he63b:	data_out=16'h8a00;
17'he63c:	data_out=16'h8a00;
17'he63d:	data_out=16'h9f9;
17'he63e:	data_out=16'ha00;
17'he63f:	data_out=16'h9e5;
17'he640:	data_out=16'h9e0;
17'he641:	data_out=16'h8a00;
17'he642:	data_out=16'h8770;
17'he643:	data_out=16'ha00;
17'he644:	data_out=16'h89fc;
17'he645:	data_out=16'h88e0;
17'he646:	data_out=16'h8a00;
17'he647:	data_out=16'h89f8;
17'he648:	data_out=16'h675;
17'he649:	data_out=16'h9fe;
17'he64a:	data_out=16'h8a00;
17'he64b:	data_out=16'h57f;
17'he64c:	data_out=16'ha00;
17'he64d:	data_out=16'ha00;
17'he64e:	data_out=16'h8a00;
17'he64f:	data_out=16'ha00;
17'he650:	data_out=16'ha00;
17'he651:	data_out=16'h8a00;
17'he652:	data_out=16'h89f9;
17'he653:	data_out=16'h8a00;
17'he654:	data_out=16'h86aa;
17'he655:	data_out=16'h89f2;
17'he656:	data_out=16'h8a00;
17'he657:	data_out=16'h9d3;
17'he658:	data_out=16'h8a00;
17'he659:	data_out=16'ha00;
17'he65a:	data_out=16'h8a00;
17'he65b:	data_out=16'h89b0;
17'he65c:	data_out=16'h8a00;
17'he65d:	data_out=16'h9cd;
17'he65e:	data_out=16'he0;
17'he65f:	data_out=16'h876f;
17'he660:	data_out=16'h8a00;
17'he661:	data_out=16'h9f0;
17'he662:	data_out=16'h89d2;
17'he663:	data_out=16'h8a00;
17'he664:	data_out=16'h8a00;
17'he665:	data_out=16'h86d2;
17'he666:	data_out=16'h8a00;
17'he667:	data_out=16'ha00;
17'he668:	data_out=16'ha00;
17'he669:	data_out=16'h8a00;
17'he66a:	data_out=16'ha00;
17'he66b:	data_out=16'h9ff;
17'he66c:	data_out=16'h8a00;
17'he66d:	data_out=16'h8a00;
17'he66e:	data_out=16'ha00;
17'he66f:	data_out=16'h250;
17'he670:	data_out=16'ha00;
17'he671:	data_out=16'h8a00;
17'he672:	data_out=16'ha00;
17'he673:	data_out=16'h9e2;
17'he674:	data_out=16'h8a00;
17'he675:	data_out=16'h9c5;
17'he676:	data_out=16'h89c5;
17'he677:	data_out=16'h879b;
17'he678:	data_out=16'ha00;
17'he679:	data_out=16'h8a00;
17'he67a:	data_out=16'h8a00;
17'he67b:	data_out=16'ha00;
17'he67c:	data_out=16'h8a00;
17'he67d:	data_out=16'h9ff;
17'he67e:	data_out=16'ha00;
17'he67f:	data_out=16'ha00;
17'he680:	data_out=16'h8a00;
17'he681:	data_out=16'h89ff;
17'he682:	data_out=16'h8a00;
17'he683:	data_out=16'h939;
17'he684:	data_out=16'h87a1;
17'he685:	data_out=16'ha00;
17'he686:	data_out=16'ha00;
17'he687:	data_out=16'h8a00;
17'he688:	data_out=16'h8a00;
17'he689:	data_out=16'h89da;
17'he68a:	data_out=16'h8832;
17'he68b:	data_out=16'h8a00;
17'he68c:	data_out=16'h8a00;
17'he68d:	data_out=16'h8a00;
17'he68e:	data_out=16'ha00;
17'he68f:	data_out=16'h8a00;
17'he690:	data_out=16'h968;
17'he691:	data_out=16'ha00;
17'he692:	data_out=16'h8a00;
17'he693:	data_out=16'h14d;
17'he694:	data_out=16'h954;
17'he695:	data_out=16'h83a8;
17'he696:	data_out=16'h8294;
17'he697:	data_out=16'h21f;
17'he698:	data_out=16'h8a00;
17'he699:	data_out=16'h8a00;
17'he69a:	data_out=16'ha00;
17'he69b:	data_out=16'h8a00;
17'he69c:	data_out=16'h854;
17'he69d:	data_out=16'h8a00;
17'he69e:	data_out=16'h9a5;
17'he69f:	data_out=16'h9fe;
17'he6a0:	data_out=16'h9f1;
17'he6a1:	data_out=16'ha00;
17'he6a2:	data_out=16'ha00;
17'he6a3:	data_out=16'h8a00;
17'he6a4:	data_out=16'h8a00;
17'he6a5:	data_out=16'h9bb;
17'he6a6:	data_out=16'h8a00;
17'he6a7:	data_out=16'h8a00;
17'he6a8:	data_out=16'ha00;
17'he6a9:	data_out=16'h9bd;
17'he6aa:	data_out=16'h856b;
17'he6ab:	data_out=16'h8a00;
17'he6ac:	data_out=16'h58d;
17'he6ad:	data_out=16'h9bb;
17'he6ae:	data_out=16'h9f6;
17'he6af:	data_out=16'h956;
17'he6b0:	data_out=16'h8a00;
17'he6b1:	data_out=16'h89fd;
17'he6b2:	data_out=16'h7e;
17'he6b3:	data_out=16'h9b5;
17'he6b4:	data_out=16'h8a00;
17'he6b5:	data_out=16'h8a00;
17'he6b6:	data_out=16'h8a00;
17'he6b7:	data_out=16'h8a00;
17'he6b8:	data_out=16'ha00;
17'he6b9:	data_out=16'h9bb;
17'he6ba:	data_out=16'h8a00;
17'he6bb:	data_out=16'h8a00;
17'he6bc:	data_out=16'h8244;
17'he6bd:	data_out=16'ha00;
17'he6be:	data_out=16'ha00;
17'he6bf:	data_out=16'ha00;
17'he6c0:	data_out=16'h9cc;
17'he6c1:	data_out=16'h8a00;
17'he6c2:	data_out=16'h8a00;
17'he6c3:	data_out=16'ha00;
17'he6c4:	data_out=16'h89ff;
17'he6c5:	data_out=16'h837e;
17'he6c6:	data_out=16'h8a00;
17'he6c7:	data_out=16'h8a00;
17'he6c8:	data_out=16'h97b;
17'he6c9:	data_out=16'h958;
17'he6ca:	data_out=16'h8a00;
17'he6cb:	data_out=16'h8a00;
17'he6cc:	data_out=16'h9fb;
17'he6cd:	data_out=16'ha00;
17'he6ce:	data_out=16'h812d;
17'he6cf:	data_out=16'h893c;
17'he6d0:	data_out=16'h9fa;
17'he6d1:	data_out=16'h89ee;
17'he6d2:	data_out=16'h8a00;
17'he6d3:	data_out=16'h82e5;
17'he6d4:	data_out=16'h9ad;
17'he6d5:	data_out=16'h89ef;
17'he6d6:	data_out=16'h8a00;
17'he6d7:	data_out=16'h99a;
17'he6d8:	data_out=16'h8a00;
17'he6d9:	data_out=16'ha00;
17'he6da:	data_out=16'h8a00;
17'he6db:	data_out=16'h89fa;
17'he6dc:	data_out=16'h86a;
17'he6dd:	data_out=16'ha00;
17'he6de:	data_out=16'ha00;
17'he6df:	data_out=16'h9f9;
17'he6e0:	data_out=16'h8a00;
17'he6e1:	data_out=16'h9f7;
17'he6e2:	data_out=16'h133;
17'he6e3:	data_out=16'h982;
17'he6e4:	data_out=16'h8a00;
17'he6e5:	data_out=16'h8a00;
17'he6e6:	data_out=16'h8a00;
17'he6e7:	data_out=16'ha00;
17'he6e8:	data_out=16'ha00;
17'he6e9:	data_out=16'h8a00;
17'he6ea:	data_out=16'ha00;
17'he6eb:	data_out=16'ha00;
17'he6ec:	data_out=16'h89fe;
17'he6ed:	data_out=16'h98f;
17'he6ee:	data_out=16'ha00;
17'he6ef:	data_out=16'h96b;
17'he6f0:	data_out=16'ha00;
17'he6f1:	data_out=16'h8a00;
17'he6f2:	data_out=16'ha00;
17'he6f3:	data_out=16'ha00;
17'he6f4:	data_out=16'h8a00;
17'he6f5:	data_out=16'h9db;
17'he6f6:	data_out=16'h8a00;
17'he6f7:	data_out=16'h8555;
17'he6f8:	data_out=16'ha00;
17'he6f9:	data_out=16'h83a6;
17'he6fa:	data_out=16'h960;
17'he6fb:	data_out=16'ha00;
17'he6fc:	data_out=16'h8a00;
17'he6fd:	data_out=16'ha00;
17'he6fe:	data_out=16'ha00;
17'he6ff:	data_out=16'ha00;
17'he700:	data_out=16'h8a00;
17'he701:	data_out=16'h8a00;
17'he702:	data_out=16'h8a00;
17'he703:	data_out=16'h9ba;
17'he704:	data_out=16'h89f9;
17'he705:	data_out=16'h9dd;
17'he706:	data_out=16'ha00;
17'he707:	data_out=16'h8a00;
17'he708:	data_out=16'h8a00;
17'he709:	data_out=16'h816;
17'he70a:	data_out=16'h8a00;
17'he70b:	data_out=16'h8a00;
17'he70c:	data_out=16'h8a00;
17'he70d:	data_out=16'h1ce;
17'he70e:	data_out=16'ha00;
17'he70f:	data_out=16'h8927;
17'he710:	data_out=16'h91a;
17'he711:	data_out=16'h8198;
17'he712:	data_out=16'h7d0;
17'he713:	data_out=16'h9e5;
17'he714:	data_out=16'h9ca;
17'he715:	data_out=16'h9cf;
17'he716:	data_out=16'h98f;
17'he717:	data_out=16'h9b3;
17'he718:	data_out=16'h8a00;
17'he719:	data_out=16'h8a00;
17'he71a:	data_out=16'h9f2;
17'he71b:	data_out=16'h8a00;
17'he71c:	data_out=16'h8f7;
17'he71d:	data_out=16'h8a00;
17'he71e:	data_out=16'h9ef;
17'he71f:	data_out=16'ha00;
17'he720:	data_out=16'h9d6;
17'he721:	data_out=16'ha00;
17'he722:	data_out=16'ha00;
17'he723:	data_out=16'h8a00;
17'he724:	data_out=16'h8a00;
17'he725:	data_out=16'h942;
17'he726:	data_out=16'h8a00;
17'he727:	data_out=16'h8a00;
17'he728:	data_out=16'ha00;
17'he729:	data_out=16'h844;
17'he72a:	data_out=16'h83c0;
17'he72b:	data_out=16'h8a00;
17'he72c:	data_out=16'h9d4;
17'he72d:	data_out=16'h8a00;
17'he72e:	data_out=16'h9df;
17'he72f:	data_out=16'h98d;
17'he730:	data_out=16'h8a00;
17'he731:	data_out=16'h8a00;
17'he732:	data_out=16'h89f8;
17'he733:	data_out=16'h9fe;
17'he734:	data_out=16'h8a00;
17'he735:	data_out=16'h8a00;
17'he736:	data_out=16'h8a00;
17'he737:	data_out=16'h8a00;
17'he738:	data_out=16'ha00;
17'he739:	data_out=16'ha00;
17'he73a:	data_out=16'h43d;
17'he73b:	data_out=16'h8a00;
17'he73c:	data_out=16'h89fe;
17'he73d:	data_out=16'h9de;
17'he73e:	data_out=16'ha00;
17'he73f:	data_out=16'h9df;
17'he740:	data_out=16'h959;
17'he741:	data_out=16'h8a00;
17'he742:	data_out=16'h8a00;
17'he743:	data_out=16'ha00;
17'he744:	data_out=16'h8a00;
17'he745:	data_out=16'h9d1;
17'he746:	data_out=16'h8a00;
17'he747:	data_out=16'h8a00;
17'he748:	data_out=16'h9ca;
17'he749:	data_out=16'h8570;
17'he74a:	data_out=16'h8a00;
17'he74b:	data_out=16'h8a00;
17'he74c:	data_out=16'h9ad;
17'he74d:	data_out=16'ha00;
17'he74e:	data_out=16'h4f3;
17'he74f:	data_out=16'h89f4;
17'he750:	data_out=16'ha00;
17'he751:	data_out=16'h68e;
17'he752:	data_out=16'h8a00;
17'he753:	data_out=16'h8a00;
17'he754:	data_out=16'h941;
17'he755:	data_out=16'h8f4;
17'he756:	data_out=16'h8a00;
17'he757:	data_out=16'h7fb;
17'he758:	data_out=16'h89fe;
17'he759:	data_out=16'h9fb;
17'he75a:	data_out=16'h89fe;
17'he75b:	data_out=16'h8a00;
17'he75c:	data_out=16'h62a;
17'he75d:	data_out=16'h9fd;
17'he75e:	data_out=16'ha00;
17'he75f:	data_out=16'h9f9;
17'he760:	data_out=16'h8a00;
17'he761:	data_out=16'h82df;
17'he762:	data_out=16'h942;
17'he763:	data_out=16'h9dc;
17'he764:	data_out=16'h8a00;
17'he765:	data_out=16'h8a00;
17'he766:	data_out=16'h8a00;
17'he767:	data_out=16'ha00;
17'he768:	data_out=16'ha00;
17'he769:	data_out=16'h8a00;
17'he76a:	data_out=16'ha00;
17'he76b:	data_out=16'h9fb;
17'he76c:	data_out=16'h8a00;
17'he76d:	data_out=16'h9e2;
17'he76e:	data_out=16'ha00;
17'he76f:	data_out=16'h980;
17'he770:	data_out=16'ha00;
17'he771:	data_out=16'h8321;
17'he772:	data_out=16'h9ff;
17'he773:	data_out=16'h9fe;
17'he774:	data_out=16'h8a00;
17'he775:	data_out=16'h8954;
17'he776:	data_out=16'h8a00;
17'he777:	data_out=16'h880;
17'he778:	data_out=16'ha00;
17'he779:	data_out=16'h6a9;
17'he77a:	data_out=16'h9ca;
17'he77b:	data_out=16'ha00;
17'he77c:	data_out=16'h8a00;
17'he77d:	data_out=16'ha00;
17'he77e:	data_out=16'h9fe;
17'he77f:	data_out=16'ha00;
17'he780:	data_out=16'h8a00;
17'he781:	data_out=16'h8a00;
17'he782:	data_out=16'h8a00;
17'he783:	data_out=16'h980;
17'he784:	data_out=16'h8a00;
17'he785:	data_out=16'h8a00;
17'he786:	data_out=16'ha00;
17'he787:	data_out=16'h8a00;
17'he788:	data_out=16'h8a00;
17'he789:	data_out=16'h95d;
17'he78a:	data_out=16'h8a00;
17'he78b:	data_out=16'h8a00;
17'he78c:	data_out=16'h8a00;
17'he78d:	data_out=16'h8029;
17'he78e:	data_out=16'h9ff;
17'he78f:	data_out=16'h976;
17'he790:	data_out=16'h9b5;
17'he791:	data_out=16'h8775;
17'he792:	data_out=16'h9d0;
17'he793:	data_out=16'h9f3;
17'he794:	data_out=16'h9b7;
17'he795:	data_out=16'h89b3;
17'he796:	data_out=16'h8818;
17'he797:	data_out=16'h99e;
17'he798:	data_out=16'h823d;
17'he799:	data_out=16'h8a00;
17'he79a:	data_out=16'h89f7;
17'he79b:	data_out=16'h8a00;
17'he79c:	data_out=16'h78e;
17'he79d:	data_out=16'h8a00;
17'he79e:	data_out=16'h9ca;
17'he79f:	data_out=16'h9d0;
17'he7a0:	data_out=16'h954;
17'he7a1:	data_out=16'ha00;
17'he7a2:	data_out=16'h9e6;
17'he7a3:	data_out=16'h8a00;
17'he7a4:	data_out=16'h8a00;
17'he7a5:	data_out=16'h95c;
17'he7a6:	data_out=16'h8a00;
17'he7a7:	data_out=16'h8a00;
17'he7a8:	data_out=16'ha00;
17'he7a9:	data_out=16'h89fa;
17'he7aa:	data_out=16'h433;
17'he7ab:	data_out=16'h8a00;
17'he7ac:	data_out=16'h8601;
17'he7ad:	data_out=16'h8751;
17'he7ae:	data_out=16'h9bb;
17'he7af:	data_out=16'h957;
17'he7b0:	data_out=16'h8a00;
17'he7b1:	data_out=16'h8a00;
17'he7b2:	data_out=16'h8a00;
17'he7b3:	data_out=16'ha00;
17'he7b4:	data_out=16'h8a00;
17'he7b5:	data_out=16'h8a00;
17'he7b6:	data_out=16'h8a00;
17'he7b7:	data_out=16'h89ff;
17'he7b8:	data_out=16'ha00;
17'he7b9:	data_out=16'ha00;
17'he7ba:	data_out=16'h8cc;
17'he7bb:	data_out=16'h8a00;
17'he7bc:	data_out=16'h8a00;
17'he7bd:	data_out=16'h993;
17'he7be:	data_out=16'ha00;
17'he7bf:	data_out=16'h8a00;
17'he7c0:	data_out=16'h8a00;
17'he7c1:	data_out=16'h8a00;
17'he7c2:	data_out=16'h8a00;
17'he7c3:	data_out=16'h9c4;
17'he7c4:	data_out=16'h8a00;
17'he7c5:	data_out=16'h8998;
17'he7c6:	data_out=16'h8a00;
17'he7c7:	data_out=16'h9a7;
17'he7c8:	data_out=16'h9f0;
17'he7c9:	data_out=16'h879d;
17'he7ca:	data_out=16'h8a00;
17'he7cb:	data_out=16'h8a00;
17'he7cc:	data_out=16'h9e5;
17'he7cd:	data_out=16'ha00;
17'he7ce:	data_out=16'h9c7;
17'he7cf:	data_out=16'h89e1;
17'he7d0:	data_out=16'h9d1;
17'he7d1:	data_out=16'h8473;
17'he7d2:	data_out=16'h8a00;
17'he7d3:	data_out=16'h8a00;
17'he7d4:	data_out=16'h8e3;
17'he7d5:	data_out=16'h81af;
17'he7d6:	data_out=16'h8a00;
17'he7d7:	data_out=16'h92c;
17'he7d8:	data_out=16'h89fb;
17'he7d9:	data_out=16'h9a1;
17'he7da:	data_out=16'h89f8;
17'he7db:	data_out=16'h8a00;
17'he7dc:	data_out=16'h8a00;
17'he7dd:	data_out=16'h9f5;
17'he7de:	data_out=16'ha00;
17'he7df:	data_out=16'h9fb;
17'he7e0:	data_out=16'h8a00;
17'he7e1:	data_out=16'h8a00;
17'he7e2:	data_out=16'h3aa;
17'he7e3:	data_out=16'h9f2;
17'he7e4:	data_out=16'h8a00;
17'he7e5:	data_out=16'h8a00;
17'he7e6:	data_out=16'h8a00;
17'he7e7:	data_out=16'h967;
17'he7e8:	data_out=16'ha00;
17'he7e9:	data_out=16'h8a00;
17'he7ea:	data_out=16'h9fd;
17'he7eb:	data_out=16'h9bc;
17'he7ec:	data_out=16'h8a00;
17'he7ed:	data_out=16'h9f7;
17'he7ee:	data_out=16'h9fd;
17'he7ef:	data_out=16'h8a00;
17'he7f0:	data_out=16'h9fe;
17'he7f1:	data_out=16'h8a7;
17'he7f2:	data_out=16'h9d1;
17'he7f3:	data_out=16'h962;
17'he7f4:	data_out=16'h8a00;
17'he7f5:	data_out=16'h8a00;
17'he7f6:	data_out=16'h8a00;
17'he7f7:	data_out=16'h94a;
17'he7f8:	data_out=16'h180;
17'he7f9:	data_out=16'h537;
17'he7fa:	data_out=16'h9cc;
17'he7fb:	data_out=16'ha00;
17'he7fc:	data_out=16'h935;
17'he7fd:	data_out=16'h9fe;
17'he7fe:	data_out=16'ha00;
17'he7ff:	data_out=16'ha00;
17'he800:	data_out=16'h89e3;
17'he801:	data_out=16'h8a00;
17'he802:	data_out=16'h89e8;
17'he803:	data_out=16'h8180;
17'he804:	data_out=16'h8a00;
17'he805:	data_out=16'h8a00;
17'he806:	data_out=16'h9f6;
17'he807:	data_out=16'h8a00;
17'he808:	data_out=16'h8a00;
17'he809:	data_out=16'h9b1;
17'he80a:	data_out=16'h8a00;
17'he80b:	data_out=16'h9f1;
17'he80c:	data_out=16'h8a00;
17'he80d:	data_out=16'h89e7;
17'he80e:	data_out=16'h9fb;
17'he80f:	data_out=16'h9ae;
17'he810:	data_out=16'h9cf;
17'he811:	data_out=16'h8427;
17'he812:	data_out=16'h9d9;
17'he813:	data_out=16'ha00;
17'he814:	data_out=16'h9cd;
17'he815:	data_out=16'h8a00;
17'he816:	data_out=16'h8a00;
17'he817:	data_out=16'h9bc;
17'he818:	data_out=16'h9cd;
17'he819:	data_out=16'h89b6;
17'he81a:	data_out=16'h8a00;
17'he81b:	data_out=16'h89fc;
17'he81c:	data_out=16'ha6;
17'he81d:	data_out=16'h8a00;
17'he81e:	data_out=16'h9eb;
17'he81f:	data_out=16'h9ae;
17'he820:	data_out=16'h848e;
17'he821:	data_out=16'h9fc;
17'he822:	data_out=16'h9c7;
17'he823:	data_out=16'h8a00;
17'he824:	data_out=16'h8a00;
17'he825:	data_out=16'h9af;
17'he826:	data_out=16'h8a00;
17'he827:	data_out=16'h8a00;
17'he828:	data_out=16'h9fb;
17'he829:	data_out=16'h89ff;
17'he82a:	data_out=16'h55a;
17'he82b:	data_out=16'h89fd;
17'he82c:	data_out=16'h89fb;
17'he82d:	data_out=16'h935;
17'he82e:	data_out=16'h953;
17'he82f:	data_out=16'h888e;
17'he830:	data_out=16'h89da;
17'he831:	data_out=16'h8a00;
17'he832:	data_out=16'h8a00;
17'he833:	data_out=16'ha00;
17'he834:	data_out=16'h8a00;
17'he835:	data_out=16'h8a00;
17'he836:	data_out=16'h8a00;
17'he837:	data_out=16'h89f8;
17'he838:	data_out=16'ha00;
17'he839:	data_out=16'ha00;
17'he83a:	data_out=16'h9bf;
17'he83b:	data_out=16'h8a00;
17'he83c:	data_out=16'h8a00;
17'he83d:	data_out=16'h9db;
17'he83e:	data_out=16'h9fb;
17'he83f:	data_out=16'h8a00;
17'he840:	data_out=16'h8a00;
17'he841:	data_out=16'h89fe;
17'he842:	data_out=16'h89eb;
17'he843:	data_out=16'h904;
17'he844:	data_out=16'h8a00;
17'he845:	data_out=16'h8a00;
17'he846:	data_out=16'h8a00;
17'he847:	data_out=16'h9f0;
17'he848:	data_out=16'h9db;
17'he849:	data_out=16'h993;
17'he84a:	data_out=16'h8a00;
17'he84b:	data_out=16'h89c9;
17'he84c:	data_out=16'h9ce;
17'he84d:	data_out=16'h9ea;
17'he84e:	data_out=16'h9bd;
17'he84f:	data_out=16'h9cd;
17'he850:	data_out=16'h82ed;
17'he851:	data_out=16'h88d8;
17'he852:	data_out=16'h8a00;
17'he853:	data_out=16'h89fd;
17'he854:	data_out=16'h8020;
17'he855:	data_out=16'h85d9;
17'he856:	data_out=16'h8a00;
17'he857:	data_out=16'h998;
17'he858:	data_out=16'h89d4;
17'he859:	data_out=16'h88d7;
17'he85a:	data_out=16'h8111;
17'he85b:	data_out=16'h8a00;
17'he85c:	data_out=16'h8a00;
17'he85d:	data_out=16'h881e;
17'he85e:	data_out=16'h805d;
17'he85f:	data_out=16'h9fa;
17'he860:	data_out=16'h8a00;
17'he861:	data_out=16'h8a00;
17'he862:	data_out=16'h81aa;
17'he863:	data_out=16'h9f9;
17'he864:	data_out=16'h8a00;
17'he865:	data_out=16'h8a00;
17'he866:	data_out=16'h9e6;
17'he867:	data_out=16'h8a00;
17'he868:	data_out=16'h9fc;
17'he869:	data_out=16'h81e9;
17'he86a:	data_out=16'h9fb;
17'he86b:	data_out=16'h87b1;
17'he86c:	data_out=16'h89dc;
17'he86d:	data_out=16'h9ff;
17'he86e:	data_out=16'h9fb;
17'he86f:	data_out=16'h8a00;
17'he870:	data_out=16'h9fb;
17'he871:	data_out=16'h7a4;
17'he872:	data_out=16'h9f1;
17'he873:	data_out=16'h8961;
17'he874:	data_out=16'h89f8;
17'he875:	data_out=16'h8a00;
17'he876:	data_out=16'h8a00;
17'he877:	data_out=16'h9b9;
17'he878:	data_out=16'h89f5;
17'he879:	data_out=16'h73f;
17'he87a:	data_out=16'h9e0;
17'he87b:	data_out=16'h9fb;
17'he87c:	data_out=16'h9b6;
17'he87d:	data_out=16'h9db;
17'he87e:	data_out=16'ha00;
17'he87f:	data_out=16'h9ee;
17'he880:	data_out=16'h89c7;
17'he881:	data_out=16'h89f3;
17'he882:	data_out=16'h9fc;
17'he883:	data_out=16'h887a;
17'he884:	data_out=16'h89f2;
17'he885:	data_out=16'h8a00;
17'he886:	data_out=16'h9f4;
17'he887:	data_out=16'h975;
17'he888:	data_out=16'h9f9;
17'he889:	data_out=16'ha00;
17'he88a:	data_out=16'h89d5;
17'he88b:	data_out=16'ha00;
17'he88c:	data_out=16'h979;
17'he88d:	data_out=16'h89db;
17'he88e:	data_out=16'ha00;
17'he88f:	data_out=16'h9ff;
17'he890:	data_out=16'h9ee;
17'he891:	data_out=16'h17d;
17'he892:	data_out=16'h9fb;
17'he893:	data_out=16'h9fd;
17'he894:	data_out=16'h9fb;
17'he895:	data_out=16'h89ea;
17'he896:	data_out=16'h89e8;
17'he897:	data_out=16'h3fe;
17'he898:	data_out=16'h9fd;
17'he899:	data_out=16'ha00;
17'he89a:	data_out=16'h8a00;
17'he89b:	data_out=16'h9ff;
17'he89c:	data_out=16'h89ae;
17'he89d:	data_out=16'h89b0;
17'he89e:	data_out=16'ha00;
17'he89f:	data_out=16'h9dc;
17'he8a0:	data_out=16'h877f;
17'he8a1:	data_out=16'ha00;
17'he8a2:	data_out=16'h9e8;
17'he8a3:	data_out=16'h683;
17'he8a4:	data_out=16'h670;
17'he8a5:	data_out=16'h9f9;
17'he8a6:	data_out=16'h9fc;
17'he8a7:	data_out=16'h8600;
17'he8a8:	data_out=16'ha00;
17'he8a9:	data_out=16'h89e9;
17'he8aa:	data_out=16'h9fe;
17'he8ab:	data_out=16'h9ee;
17'he8ac:	data_out=16'h89f3;
17'he8ad:	data_out=16'ha00;
17'he8ae:	data_out=16'h9e4;
17'he8af:	data_out=16'h8928;
17'he8b0:	data_out=16'h8117;
17'he8b1:	data_out=16'h89ff;
17'he8b2:	data_out=16'h89ff;
17'he8b3:	data_out=16'ha00;
17'he8b4:	data_out=16'h89f4;
17'he8b5:	data_out=16'h8904;
17'he8b6:	data_out=16'ha00;
17'he8b7:	data_out=16'h9f6;
17'he8b8:	data_out=16'h5de;
17'he8b9:	data_out=16'ha00;
17'he8ba:	data_out=16'ha00;
17'he8bb:	data_out=16'h89f9;
17'he8bc:	data_out=16'h8a00;
17'he8bd:	data_out=16'h833c;
17'he8be:	data_out=16'ha00;
17'he8bf:	data_out=16'h8a00;
17'he8c0:	data_out=16'h89fd;
17'he8c1:	data_out=16'h89d5;
17'he8c2:	data_out=16'h80c3;
17'he8c3:	data_out=16'h86f5;
17'he8c4:	data_out=16'h89ef;
17'he8c5:	data_out=16'h89ec;
17'he8c6:	data_out=16'h8536;
17'he8c7:	data_out=16'ha00;
17'he8c8:	data_out=16'h9f2;
17'he8c9:	data_out=16'h9e8;
17'he8ca:	data_out=16'h9cc;
17'he8cb:	data_out=16'h880a;
17'he8cc:	data_out=16'h9fd;
17'he8cd:	data_out=16'h9f9;
17'he8ce:	data_out=16'h9fd;
17'he8cf:	data_out=16'ha00;
17'he8d0:	data_out=16'h89a3;
17'he8d1:	data_out=16'h899a;
17'he8d2:	data_out=16'h86ec;
17'he8d3:	data_out=16'h102;
17'he8d4:	data_out=16'h9fa;
17'he8d5:	data_out=16'h633;
17'he8d6:	data_out=16'h9f9;
17'he8d7:	data_out=16'ha00;
17'he8d8:	data_out=16'h899c;
17'he8d9:	data_out=16'h8961;
17'he8da:	data_out=16'h9eb;
17'he8db:	data_out=16'h89b4;
17'he8dc:	data_out=16'h8a00;
17'he8dd:	data_out=16'h892c;
17'he8de:	data_out=16'h885c;
17'he8df:	data_out=16'ha00;
17'he8e0:	data_out=16'h9d9;
17'he8e1:	data_out=16'h8a00;
17'he8e2:	data_out=16'h9eb;
17'he8e3:	data_out=16'ha00;
17'he8e4:	data_out=16'h89f9;
17'he8e5:	data_out=16'h8981;
17'he8e6:	data_out=16'ha00;
17'he8e7:	data_out=16'h89c8;
17'he8e8:	data_out=16'ha00;
17'he8e9:	data_out=16'h9ff;
17'he8ea:	data_out=16'ha00;
17'he8eb:	data_out=16'h896a;
17'he8ec:	data_out=16'h89a0;
17'he8ed:	data_out=16'ha00;
17'he8ee:	data_out=16'ha00;
17'he8ef:	data_out=16'h8a00;
17'he8f0:	data_out=16'ha00;
17'he8f1:	data_out=16'h9ee;
17'he8f2:	data_out=16'h8943;
17'he8f3:	data_out=16'h89f1;
17'he8f4:	data_out=16'h8344;
17'he8f5:	data_out=16'h8a00;
17'he8f6:	data_out=16'h9e8;
17'he8f7:	data_out=16'ha00;
17'he8f8:	data_out=16'h8a00;
17'he8f9:	data_out=16'h9fd;
17'he8fa:	data_out=16'h9fd;
17'he8fb:	data_out=16'ha00;
17'he8fc:	data_out=16'h9fb;
17'he8fd:	data_out=16'h9d2;
17'he8fe:	data_out=16'ha00;
17'he8ff:	data_out=16'h8a00;
17'he900:	data_out=16'h89ef;
17'he901:	data_out=16'h8a00;
17'he902:	data_out=16'h9fa;
17'he903:	data_out=16'h89a9;
17'he904:	data_out=16'h89e7;
17'he905:	data_out=16'h8a00;
17'he906:	data_out=16'h833e;
17'he907:	data_out=16'ha00;
17'he908:	data_out=16'ha00;
17'he909:	data_out=16'ha00;
17'he90a:	data_out=16'h8a00;
17'he90b:	data_out=16'ha00;
17'he90c:	data_out=16'h9e9;
17'he90d:	data_out=16'h89d8;
17'he90e:	data_out=16'h9fe;
17'he90f:	data_out=16'ha00;
17'he910:	data_out=16'h957;
17'he911:	data_out=16'h882a;
17'he912:	data_out=16'h9f7;
17'he913:	data_out=16'h866d;
17'he914:	data_out=16'h9fa;
17'he915:	data_out=16'h89ff;
17'he916:	data_out=16'h89fa;
17'he917:	data_out=16'h895d;
17'he918:	data_out=16'h9ff;
17'he919:	data_out=16'ha00;
17'he91a:	data_out=16'h8a00;
17'he91b:	data_out=16'ha00;
17'he91c:	data_out=16'h8a00;
17'he91d:	data_out=16'h89f2;
17'he91e:	data_out=16'h9fc;
17'he91f:	data_out=16'h9f1;
17'he920:	data_out=16'h89b5;
17'he921:	data_out=16'h9fd;
17'he922:	data_out=16'h8795;
17'he923:	data_out=16'ha00;
17'he924:	data_out=16'ha00;
17'he925:	data_out=16'h7ba;
17'he926:	data_out=16'h9f6;
17'he927:	data_out=16'h5fa;
17'he928:	data_out=16'h9fd;
17'he929:	data_out=16'h89d0;
17'he92a:	data_out=16'h9fe;
17'he92b:	data_out=16'ha00;
17'he92c:	data_out=16'h8a00;
17'he92d:	data_out=16'h438;
17'he92e:	data_out=16'h9e3;
17'he92f:	data_out=16'h89eb;
17'he930:	data_out=16'h821a;
17'he931:	data_out=16'h89fe;
17'he932:	data_out=16'h89fe;
17'he933:	data_out=16'h9ff;
17'he934:	data_out=16'h89fd;
17'he935:	data_out=16'h8934;
17'he936:	data_out=16'ha00;
17'he937:	data_out=16'h9fd;
17'he938:	data_out=16'h8a00;
17'he939:	data_out=16'h9ff;
17'he93a:	data_out=16'ha00;
17'he93b:	data_out=16'h838e;
17'he93c:	data_out=16'h8a00;
17'he93d:	data_out=16'h8969;
17'he93e:	data_out=16'h9fd;
17'he93f:	data_out=16'h8a00;
17'he940:	data_out=16'h89fe;
17'he941:	data_out=16'h51f;
17'he942:	data_out=16'h873e;
17'he943:	data_out=16'h89c5;
17'he944:	data_out=16'h89dd;
17'he945:	data_out=16'h8a00;
17'he946:	data_out=16'h87de;
17'he947:	data_out=16'ha00;
17'he948:	data_out=16'h89e;
17'he949:	data_out=16'h80dd;
17'he94a:	data_out=16'ha00;
17'he94b:	data_out=16'h33d;
17'he94c:	data_out=16'h9f0;
17'he94d:	data_out=16'h84de;
17'he94e:	data_out=16'h9ff;
17'he94f:	data_out=16'h9ff;
17'he950:	data_out=16'h8a00;
17'he951:	data_out=16'h89b6;
17'he952:	data_out=16'h297;
17'he953:	data_out=16'h9a5;
17'he954:	data_out=16'h848e;
17'he955:	data_out=16'h9fc;
17'he956:	data_out=16'h8540;
17'he957:	data_out=16'h82f9;
17'he958:	data_out=16'h894b;
17'he959:	data_out=16'h89e9;
17'he95a:	data_out=16'h9ef;
17'he95b:	data_out=16'h89a4;
17'he95c:	data_out=16'h8a00;
17'he95d:	data_out=16'h89e9;
17'he95e:	data_out=16'h89f7;
17'he95f:	data_out=16'h9fe;
17'he960:	data_out=16'h84b8;
17'he961:	data_out=16'h8a00;
17'he962:	data_out=16'h9fd;
17'he963:	data_out=16'h9ff;
17'he964:	data_out=16'h89ff;
17'he965:	data_out=16'h899d;
17'he966:	data_out=16'ha00;
17'he967:	data_out=16'h93c;
17'he968:	data_out=16'h9fd;
17'he969:	data_out=16'ha00;
17'he96a:	data_out=16'h9fe;
17'he96b:	data_out=16'h89fe;
17'he96c:	data_out=16'h89ed;
17'he96d:	data_out=16'h9ff;
17'he96e:	data_out=16'h9fe;
17'he96f:	data_out=16'h89ff;
17'he970:	data_out=16'h9fe;
17'he971:	data_out=16'h9f8;
17'he972:	data_out=16'h8a00;
17'he973:	data_out=16'h8a00;
17'he974:	data_out=16'h827c;
17'he975:	data_out=16'h8a00;
17'he976:	data_out=16'ha00;
17'he977:	data_out=16'ha00;
17'he978:	data_out=16'h8a00;
17'he979:	data_out=16'h9fc;
17'he97a:	data_out=16'h9fe;
17'he97b:	data_out=16'h9fd;
17'he97c:	data_out=16'h9fe;
17'he97d:	data_out=16'h816f;
17'he97e:	data_out=16'h8af;
17'he97f:	data_out=16'h8a00;
17'he980:	data_out=16'h8a00;
17'he981:	data_out=16'h8a00;
17'he982:	data_out=16'h1c5;
17'he983:	data_out=16'h89cc;
17'he984:	data_out=16'h89db;
17'he985:	data_out=16'h8a00;
17'he986:	data_out=16'h8959;
17'he987:	data_out=16'ha00;
17'he988:	data_out=16'h9ea;
17'he989:	data_out=16'ha00;
17'he98a:	data_out=16'h8a00;
17'he98b:	data_out=16'ha00;
17'he98c:	data_out=16'ha00;
17'he98d:	data_out=16'h8a00;
17'he98e:	data_out=16'h896f;
17'he98f:	data_out=16'h9fb;
17'he990:	data_out=16'h93d;
17'he991:	data_out=16'h89f3;
17'he992:	data_out=16'h973;
17'he993:	data_out=16'h89d2;
17'he994:	data_out=16'h898b;
17'he995:	data_out=16'h8a00;
17'he996:	data_out=16'h89fb;
17'he997:	data_out=16'h89da;
17'he998:	data_out=16'h9f2;
17'he999:	data_out=16'ha00;
17'he99a:	data_out=16'h89fc;
17'he99b:	data_out=16'h9f8;
17'he99c:	data_out=16'h8a00;
17'he99d:	data_out=16'h89eb;
17'he99e:	data_out=16'h89d1;
17'he99f:	data_out=16'h40;
17'he9a0:	data_out=16'h89f2;
17'he9a1:	data_out=16'h8711;
17'he9a2:	data_out=16'h89c5;
17'he9a3:	data_out=16'ha00;
17'he9a4:	data_out=16'ha00;
17'he9a5:	data_out=16'h88df;
17'he9a6:	data_out=16'h8856;
17'he9a7:	data_out=16'h99a;
17'he9a8:	data_out=16'h8391;
17'he9a9:	data_out=16'h89d9;
17'he9aa:	data_out=16'ha00;
17'he9ab:	data_out=16'ha00;
17'he9ac:	data_out=16'h8a00;
17'he9ad:	data_out=16'h899c;
17'he9ae:	data_out=16'h9e4;
17'he9af:	data_out=16'h85e7;
17'he9b0:	data_out=16'h8672;
17'he9b1:	data_out=16'h89fd;
17'he9b2:	data_out=16'h87c2;
17'he9b3:	data_out=16'h8924;
17'he9b4:	data_out=16'h8a00;
17'he9b5:	data_out=16'h884e;
17'he9b6:	data_out=16'ha00;
17'he9b7:	data_out=16'h417;
17'he9b8:	data_out=16'h8a00;
17'he9b9:	data_out=16'h89ef;
17'he9ba:	data_out=16'ha00;
17'he9bb:	data_out=16'ha00;
17'he9bc:	data_out=16'h8a00;
17'he9bd:	data_out=16'h89fb;
17'he9be:	data_out=16'h8383;
17'he9bf:	data_out=16'h8a00;
17'he9c0:	data_out=16'h8994;
17'he9c1:	data_out=16'h92d;
17'he9c2:	data_out=16'h8322;
17'he9c3:	data_out=16'h8e7;
17'he9c4:	data_out=16'h89dd;
17'he9c5:	data_out=16'h8a00;
17'he9c6:	data_out=16'h89f7;
17'he9c7:	data_out=16'ha00;
17'he9c8:	data_out=16'h522;
17'he9c9:	data_out=16'h86fc;
17'he9ca:	data_out=16'ha00;
17'he9cb:	data_out=16'h98d;
17'he9cc:	data_out=16'h845e;
17'he9cd:	data_out=16'h898e;
17'he9ce:	data_out=16'ha00;
17'he9cf:	data_out=16'h775;
17'he9d0:	data_out=16'h89da;
17'he9d1:	data_out=16'h89ff;
17'he9d2:	data_out=16'hce;
17'he9d3:	data_out=16'h99a;
17'he9d4:	data_out=16'h835b;
17'he9d5:	data_out=16'h8555;
17'he9d6:	data_out=16'h89aa;
17'he9d7:	data_out=16'h89c4;
17'he9d8:	data_out=16'h89fa;
17'he9d9:	data_out=16'h89d6;
17'he9da:	data_out=16'h83c9;
17'he9db:	data_out=16'h89e5;
17'he9dc:	data_out=16'h8a00;
17'he9dd:	data_out=16'h89f0;
17'he9de:	data_out=16'h86a7;
17'he9df:	data_out=16'h9e1;
17'he9e0:	data_out=16'h89b2;
17'he9e1:	data_out=16'h8a00;
17'he9e2:	data_out=16'h8283;
17'he9e3:	data_out=16'h8416;
17'he9e4:	data_out=16'h89ec;
17'he9e5:	data_out=16'h1bc;
17'he9e6:	data_out=16'ha00;
17'he9e7:	data_out=16'ha00;
17'he9e8:	data_out=16'h8592;
17'he9e9:	data_out=16'h9ec;
17'he9ea:	data_out=16'h89e9;
17'he9eb:	data_out=16'h89f8;
17'he9ec:	data_out=16'h8a00;
17'he9ed:	data_out=16'h856c;
17'he9ee:	data_out=16'h89e9;
17'he9ef:	data_out=16'h89f5;
17'he9f0:	data_out=16'h89e4;
17'he9f1:	data_out=16'h9f8;
17'he9f2:	data_out=16'h8a00;
17'he9f3:	data_out=16'h8a00;
17'he9f4:	data_out=16'h8699;
17'he9f5:	data_out=16'h8a00;
17'he9f6:	data_out=16'ha00;
17'he9f7:	data_out=16'h9fa;
17'he9f8:	data_out=16'h8a00;
17'he9f9:	data_out=16'h9d3;
17'he9fa:	data_out=16'h88d9;
17'he9fb:	data_out=16'h837b;
17'he9fc:	data_out=16'h9f4;
17'he9fd:	data_out=16'h8384;
17'he9fe:	data_out=16'h89e8;
17'he9ff:	data_out=16'h8a00;
17'hea00:	data_out=16'h8a00;
17'hea01:	data_out=16'h8a00;
17'hea02:	data_out=16'h87a0;
17'hea03:	data_out=16'h89fe;
17'hea04:	data_out=16'h8465;
17'hea05:	data_out=16'h8a00;
17'hea06:	data_out=16'h8991;
17'hea07:	data_out=16'ha00;
17'hea08:	data_out=16'h9b1;
17'hea09:	data_out=16'h9f9;
17'hea0a:	data_out=16'h8a00;
17'hea0b:	data_out=16'ha00;
17'hea0c:	data_out=16'ha00;
17'hea0d:	data_out=16'h89fc;
17'hea0e:	data_out=16'h89fc;
17'hea0f:	data_out=16'h9f4;
17'hea10:	data_out=16'hc8;
17'hea11:	data_out=16'h89ff;
17'hea12:	data_out=16'h8687;
17'hea13:	data_out=16'h89f7;
17'hea14:	data_out=16'h89f0;
17'hea15:	data_out=16'h89ff;
17'hea16:	data_out=16'h89fd;
17'hea17:	data_out=16'h89f1;
17'hea18:	data_out=16'h9ca;
17'hea19:	data_out=16'ha00;
17'hea1a:	data_out=16'h89fb;
17'hea1b:	data_out=16'h278;
17'hea1c:	data_out=16'h8a00;
17'hea1d:	data_out=16'h8a00;
17'hea1e:	data_out=16'h89f7;
17'hea1f:	data_out=16'h8964;
17'hea20:	data_out=16'h89fa;
17'hea21:	data_out=16'h89fb;
17'hea22:	data_out=16'h89d7;
17'hea23:	data_out=16'ha00;
17'hea24:	data_out=16'ha00;
17'hea25:	data_out=16'h8936;
17'hea26:	data_out=16'h89de;
17'hea27:	data_out=16'h988;
17'hea28:	data_out=16'h89fb;
17'hea29:	data_out=16'h8a00;
17'hea2a:	data_out=16'h9fb;
17'hea2b:	data_out=16'ha00;
17'hea2c:	data_out=16'h89fe;
17'hea2d:	data_out=16'h89fe;
17'hea2e:	data_out=16'h4ab;
17'hea2f:	data_out=16'h85b1;
17'hea30:	data_out=16'h89c0;
17'hea31:	data_out=16'h8a00;
17'hea32:	data_out=16'h84cb;
17'hea33:	data_out=16'h89f9;
17'hea34:	data_out=16'h8a00;
17'hea35:	data_out=16'hab;
17'hea36:	data_out=16'h9e9;
17'hea37:	data_out=16'h8672;
17'hea38:	data_out=16'h8a00;
17'hea39:	data_out=16'h89fb;
17'hea3a:	data_out=16'h9f6;
17'hea3b:	data_out=16'ha00;
17'hea3c:	data_out=16'h8a00;
17'hea3d:	data_out=16'h89fc;
17'hea3e:	data_out=16'h89fb;
17'hea3f:	data_out=16'h8a00;
17'hea40:	data_out=16'h85b9;
17'hea41:	data_out=16'h965;
17'hea42:	data_out=16'h79a;
17'hea43:	data_out=16'h9ee;
17'hea44:	data_out=16'h88bc;
17'hea45:	data_out=16'h89ff;
17'hea46:	data_out=16'h8a00;
17'hea47:	data_out=16'h9fd;
17'hea48:	data_out=16'h306;
17'hea49:	data_out=16'h87b2;
17'hea4a:	data_out=16'ha00;
17'hea4b:	data_out=16'h9f3;
17'hea4c:	data_out=16'h84a6;
17'hea4d:	data_out=16'h89e4;
17'hea4e:	data_out=16'ha00;
17'hea4f:	data_out=16'h9e7;
17'hea50:	data_out=16'h89e8;
17'hea51:	data_out=16'h89fc;
17'hea52:	data_out=16'h96;
17'hea53:	data_out=16'h992;
17'hea54:	data_out=16'h8663;
17'hea55:	data_out=16'h87b0;
17'hea56:	data_out=16'h8916;
17'hea57:	data_out=16'h89f7;
17'hea58:	data_out=16'h8a00;
17'hea59:	data_out=16'h89d6;
17'hea5a:	data_out=16'h89d7;
17'hea5b:	data_out=16'h89b4;
17'hea5c:	data_out=16'h8a00;
17'hea5d:	data_out=16'h867a;
17'hea5e:	data_out=16'h859c;
17'hea5f:	data_out=16'h6c4;
17'hea60:	data_out=16'h89fd;
17'hea61:	data_out=16'h8a00;
17'hea62:	data_out=16'h823c;
17'hea63:	data_out=16'h89f1;
17'hea64:	data_out=16'h8a00;
17'hea65:	data_out=16'h60;
17'hea66:	data_out=16'ha00;
17'hea67:	data_out=16'ha00;
17'hea68:	data_out=16'h89fa;
17'hea69:	data_out=16'h9c2;
17'hea6a:	data_out=16'h89fd;
17'hea6b:	data_out=16'h89f1;
17'hea6c:	data_out=16'h8a00;
17'hea6d:	data_out=16'h89f3;
17'hea6e:	data_out=16'h89fd;
17'hea6f:	data_out=16'h85de;
17'hea70:	data_out=16'h89fc;
17'hea71:	data_out=16'h9f6;
17'hea72:	data_out=16'h8a00;
17'hea73:	data_out=16'h8a00;
17'hea74:	data_out=16'h89f8;
17'hea75:	data_out=16'h8a00;
17'hea76:	data_out=16'ha00;
17'hea77:	data_out=16'h9ed;
17'hea78:	data_out=16'h89ff;
17'hea79:	data_out=16'h9b3;
17'hea7a:	data_out=16'h89ee;
17'hea7b:	data_out=16'h89fb;
17'hea7c:	data_out=16'h9d8;
17'hea7d:	data_out=16'h8904;
17'hea7e:	data_out=16'h8a00;
17'hea7f:	data_out=16'h8a00;
17'hea80:	data_out=16'h88cc;
17'hea81:	data_out=16'h8a00;
17'hea82:	data_out=16'h8565;
17'hea83:	data_out=16'h89f7;
17'hea84:	data_out=16'ha00;
17'hea85:	data_out=16'h89ed;
17'hea86:	data_out=16'h89e5;
17'hea87:	data_out=16'ha00;
17'hea88:	data_out=16'h9be;
17'hea89:	data_out=16'h9fd;
17'hea8a:	data_out=16'h89f9;
17'hea8b:	data_out=16'ha00;
17'hea8c:	data_out=16'ha00;
17'hea8d:	data_out=16'h89f9;
17'hea8e:	data_out=16'h89fb;
17'hea8f:	data_out=16'ha00;
17'hea90:	data_out=16'h298;
17'hea91:	data_out=16'h2e5;
17'hea92:	data_out=16'h80be;
17'hea93:	data_out=16'h89a8;
17'hea94:	data_out=16'h89e5;
17'hea95:	data_out=16'h89b6;
17'hea96:	data_out=16'h8661;
17'hea97:	data_out=16'h89cb;
17'hea98:	data_out=16'h8691;
17'hea99:	data_out=16'ha00;
17'hea9a:	data_out=16'h164;
17'hea9b:	data_out=16'h8709;
17'hea9c:	data_out=16'h8a00;
17'hea9d:	data_out=16'h8859;
17'hea9e:	data_out=16'h8738;
17'hea9f:	data_out=16'h8348;
17'heaa0:	data_out=16'h816e;
17'heaa1:	data_out=16'h89fa;
17'heaa2:	data_out=16'h89e3;
17'heaa3:	data_out=16'h851c;
17'heaa4:	data_out=16'h84e4;
17'heaa5:	data_out=16'h881c;
17'heaa6:	data_out=16'h875b;
17'heaa7:	data_out=16'h9ea;
17'heaa8:	data_out=16'h89fb;
17'heaa9:	data_out=16'h8a00;
17'heaaa:	data_out=16'ha00;
17'heaab:	data_out=16'ha00;
17'heaac:	data_out=16'h879e;
17'heaad:	data_out=16'h89ff;
17'heaae:	data_out=16'ha00;
17'heaaf:	data_out=16'h9aa;
17'heab0:	data_out=16'h89e7;
17'heab1:	data_out=16'h89fa;
17'heab2:	data_out=16'h85ae;
17'heab3:	data_out=16'h89f5;
17'heab4:	data_out=16'h8a00;
17'heab5:	data_out=16'h9dc;
17'heab6:	data_out=16'h9e8;
17'heab7:	data_out=16'h832d;
17'heab8:	data_out=16'h8a00;
17'heab9:	data_out=16'h89fb;
17'heaba:	data_out=16'h9ef;
17'heabb:	data_out=16'ha00;
17'heabc:	data_out=16'h8a00;
17'heabd:	data_out=16'h8876;
17'heabe:	data_out=16'h89fb;
17'heabf:	data_out=16'h89ee;
17'heac0:	data_out=16'h883;
17'heac1:	data_out=16'h992;
17'heac2:	data_out=16'h9f1;
17'heac3:	data_out=16'h9fb;
17'heac4:	data_out=16'ha00;
17'heac5:	data_out=16'h89ab;
17'heac6:	data_out=16'h8a00;
17'heac7:	data_out=16'ha00;
17'heac8:	data_out=16'h9c5;
17'heac9:	data_out=16'h8815;
17'heaca:	data_out=16'ha00;
17'heacb:	data_out=16'h9ee;
17'heacc:	data_out=16'h9e8;
17'heacd:	data_out=16'h89ee;
17'heace:	data_out=16'ha00;
17'heacf:	data_out=16'h9ee;
17'head0:	data_out=16'h86fe;
17'head1:	data_out=16'h89fd;
17'head2:	data_out=16'h84d9;
17'head3:	data_out=16'h9f0;
17'head4:	data_out=16'h7b3;
17'head5:	data_out=16'h859a;
17'head6:	data_out=16'h8744;
17'head7:	data_out=16'h89ed;
17'head8:	data_out=16'h8a00;
17'head9:	data_out=16'h8800;
17'heada:	data_out=16'h89eb;
17'headb:	data_out=16'h6ea;
17'headc:	data_out=16'h8a00;
17'headd:	data_out=16'h9ba;
17'heade:	data_out=16'h9b8;
17'headf:	data_out=16'h594;
17'heae0:	data_out=16'h892a;
17'heae1:	data_out=16'h89e9;
17'heae2:	data_out=16'h8eb;
17'heae3:	data_out=16'h89ec;
17'heae4:	data_out=16'h89fb;
17'heae5:	data_out=16'h9d2;
17'heae6:	data_out=16'ha00;
17'heae7:	data_out=16'ha00;
17'heae8:	data_out=16'h89fa;
17'heae9:	data_out=16'h9d7;
17'heaea:	data_out=16'h89fb;
17'heaeb:	data_out=16'h865a;
17'heaec:	data_out=16'h863d;
17'heaed:	data_out=16'h89ee;
17'heaee:	data_out=16'h89fb;
17'heaef:	data_out=16'h1a;
17'heaf0:	data_out=16'h89fb;
17'heaf1:	data_out=16'ha00;
17'heaf2:	data_out=16'h89fd;
17'heaf3:	data_out=16'h89ea;
17'heaf4:	data_out=16'h89fb;
17'heaf5:	data_out=16'h8a00;
17'heaf6:	data_out=16'ha00;
17'heaf7:	data_out=16'h9fb;
17'heaf8:	data_out=16'h83c6;
17'heaf9:	data_out=16'h9af;
17'heafa:	data_out=16'h8972;
17'heafb:	data_out=16'h89fb;
17'heafc:	data_out=16'h480;
17'heafd:	data_out=16'h4b8;
17'heafe:	data_out=16'h8a00;
17'heaff:	data_out=16'h8a00;
17'heb00:	data_out=16'h89fb;
17'heb01:	data_out=16'h847b;
17'heb02:	data_out=16'h897c;
17'heb03:	data_out=16'h89f7;
17'heb04:	data_out=16'ha00;
17'heb05:	data_out=16'h89d7;
17'heb06:	data_out=16'h89f1;
17'heb07:	data_out=16'ha00;
17'heb08:	data_out=16'h9ec;
17'heb09:	data_out=16'h9d7;
17'heb0a:	data_out=16'h89e8;
17'heb0b:	data_out=16'ha00;
17'heb0c:	data_out=16'h9f4;
17'heb0d:	data_out=16'h89fd;
17'heb0e:	data_out=16'h89fa;
17'heb0f:	data_out=16'h8f0;
17'heb10:	data_out=16'h89bb;
17'heb11:	data_out=16'h9af;
17'heb12:	data_out=16'h14e;
17'heb13:	data_out=16'h89fa;
17'heb14:	data_out=16'h89e0;
17'heb15:	data_out=16'h89fe;
17'heb16:	data_out=16'h88ff;
17'heb17:	data_out=16'h87d9;
17'heb18:	data_out=16'h89ff;
17'heb19:	data_out=16'ha00;
17'heb1a:	data_out=16'h9fd;
17'heb1b:	data_out=16'h885d;
17'heb1c:	data_out=16'h8a00;
17'heb1d:	data_out=16'h85e;
17'heb1e:	data_out=16'h89e6;
17'heb1f:	data_out=16'h2f;
17'heb20:	data_out=16'h89ec;
17'heb21:	data_out=16'h89f9;
17'heb22:	data_out=16'hb8;
17'heb23:	data_out=16'h824;
17'heb24:	data_out=16'h84c;
17'heb25:	data_out=16'h81cd;
17'heb26:	data_out=16'h71a;
17'heb27:	data_out=16'h9ef;
17'heb28:	data_out=16'h89f9;
17'heb29:	data_out=16'h8a00;
17'heb2a:	data_out=16'ha00;
17'heb2b:	data_out=16'ha00;
17'heb2c:	data_out=16'h897e;
17'heb2d:	data_out=16'h89ed;
17'heb2e:	data_out=16'ha00;
17'heb2f:	data_out=16'h8147;
17'heb30:	data_out=16'h89e6;
17'heb31:	data_out=16'h89f4;
17'heb32:	data_out=16'h88b7;
17'heb33:	data_out=16'h89f5;
17'heb34:	data_out=16'h8a00;
17'heb35:	data_out=16'h9f3;
17'heb36:	data_out=16'h3bb;
17'heb37:	data_out=16'h8628;
17'heb38:	data_out=16'h8a00;
17'heb39:	data_out=16'h89fd;
17'heb3a:	data_out=16'h9a3;
17'heb3b:	data_out=16'h9ff;
17'heb3c:	data_out=16'h89f9;
17'heb3d:	data_out=16'h89f9;
17'heb3e:	data_out=16'h89f8;
17'heb3f:	data_out=16'h89d9;
17'heb40:	data_out=16'ha00;
17'heb41:	data_out=16'h115;
17'heb42:	data_out=16'h9f6;
17'heb43:	data_out=16'h9f1;
17'heb44:	data_out=16'ha00;
17'heb45:	data_out=16'h89fe;
17'heb46:	data_out=16'h8a00;
17'heb47:	data_out=16'h9ec;
17'heb48:	data_out=16'h9aa;
17'heb49:	data_out=16'h85d7;
17'heb4a:	data_out=16'ha00;
17'heb4b:	data_out=16'h9f5;
17'heb4c:	data_out=16'h835;
17'heb4d:	data_out=16'h8322;
17'heb4e:	data_out=16'ha00;
17'heb4f:	data_out=16'h9cd;
17'heb50:	data_out=16'h89bf;
17'heb51:	data_out=16'h89ff;
17'heb52:	data_out=16'h83f9;
17'heb53:	data_out=16'ha00;
17'heb54:	data_out=16'h85a0;
17'heb55:	data_out=16'h87c3;
17'heb56:	data_out=16'h88ac;
17'heb57:	data_out=16'h89fe;
17'heb58:	data_out=16'h8a00;
17'heb59:	data_out=16'h89c4;
17'heb5a:	data_out=16'h89f1;
17'heb5b:	data_out=16'ha00;
17'heb5c:	data_out=16'h89f4;
17'heb5d:	data_out=16'h8242;
17'heb5e:	data_out=16'h211;
17'heb5f:	data_out=16'h87e9;
17'heb60:	data_out=16'h8774;
17'heb61:	data_out=16'h8594;
17'heb62:	data_out=16'h9f8;
17'heb63:	data_out=16'h8948;
17'heb64:	data_out=16'h850e;
17'heb65:	data_out=16'h9de;
17'heb66:	data_out=16'ha00;
17'heb67:	data_out=16'ha00;
17'heb68:	data_out=16'h89f8;
17'heb69:	data_out=16'h9dd;
17'heb6a:	data_out=16'h89fa;
17'heb6b:	data_out=16'h89de;
17'heb6c:	data_out=16'h89f8;
17'heb6d:	data_out=16'h89f1;
17'heb6e:	data_out=16'h89fa;
17'heb6f:	data_out=16'h9fe;
17'heb70:	data_out=16'h89fa;
17'heb71:	data_out=16'h9fe;
17'heb72:	data_out=16'h89f5;
17'heb73:	data_out=16'h89dd;
17'heb74:	data_out=16'h89f0;
17'heb75:	data_out=16'h89f7;
17'heb76:	data_out=16'ha00;
17'heb77:	data_out=16'h5c1;
17'heb78:	data_out=16'h89d5;
17'heb79:	data_out=16'h9c8;
17'heb7a:	data_out=16'h8937;
17'heb7b:	data_out=16'h89f8;
17'heb7c:	data_out=16'h89fe;
17'heb7d:	data_out=16'h3e8;
17'heb7e:	data_out=16'h8a00;
17'heb7f:	data_out=16'h8a00;
17'heb80:	data_out=16'h89f3;
17'heb81:	data_out=16'h9de;
17'heb82:	data_out=16'h89cf;
17'heb83:	data_out=16'h89f0;
17'heb84:	data_out=16'ha00;
17'heb85:	data_out=16'h89cf;
17'heb86:	data_out=16'h89fb;
17'heb87:	data_out=16'ha00;
17'heb88:	data_out=16'h43b;
17'heb89:	data_out=16'h7c8;
17'heb8a:	data_out=16'h9e9;
17'heb8b:	data_out=16'ha00;
17'heb8c:	data_out=16'h9f5;
17'heb8d:	data_out=16'h89fd;
17'heb8e:	data_out=16'h89b8;
17'heb8f:	data_out=16'h867f;
17'heb90:	data_out=16'h8a00;
17'heb91:	data_out=16'h9f1;
17'heb92:	data_out=16'h89f7;
17'heb93:	data_out=16'h89ef;
17'heb94:	data_out=16'h89ee;
17'heb95:	data_out=16'h89fb;
17'heb96:	data_out=16'h89ec;
17'heb97:	data_out=16'h89e4;
17'heb98:	data_out=16'h89fe;
17'heb99:	data_out=16'ha00;
17'heb9a:	data_out=16'h9fd;
17'heb9b:	data_out=16'h89ea;
17'heb9c:	data_out=16'h89fb;
17'heb9d:	data_out=16'h9dc;
17'heb9e:	data_out=16'h89f3;
17'heb9f:	data_out=16'h831c;
17'heba0:	data_out=16'h89fc;
17'heba1:	data_out=16'h89f5;
17'heba2:	data_out=16'h481;
17'heba3:	data_out=16'h975;
17'heba4:	data_out=16'h989;
17'heba5:	data_out=16'h8526;
17'heba6:	data_out=16'h596;
17'heba7:	data_out=16'h9fd;
17'heba8:	data_out=16'h89f6;
17'heba9:	data_out=16'h89e4;
17'hebaa:	data_out=16'h220;
17'hebab:	data_out=16'ha00;
17'hebac:	data_out=16'h89f1;
17'hebad:	data_out=16'h8255;
17'hebae:	data_out=16'h9e;
17'hebaf:	data_out=16'h88e3;
17'hebb0:	data_out=16'h86b8;
17'hebb1:	data_out=16'h9c3;
17'hebb2:	data_out=16'h81e3;
17'hebb3:	data_out=16'h8a00;
17'hebb4:	data_out=16'h8c9;
17'hebb5:	data_out=16'h9ff;
17'hebb6:	data_out=16'h8983;
17'hebb7:	data_out=16'h89cf;
17'hebb8:	data_out=16'h82e3;
17'hebb9:	data_out=16'h8a00;
17'hebba:	data_out=16'h804;
17'hebbb:	data_out=16'h9ff;
17'hebbc:	data_out=16'h89dd;
17'hebbd:	data_out=16'h89fd;
17'hebbe:	data_out=16'h89f6;
17'hebbf:	data_out=16'h89d0;
17'hebc0:	data_out=16'h662;
17'hebc1:	data_out=16'h89b2;
17'hebc2:	data_out=16'h9fd;
17'hebc3:	data_out=16'h850d;
17'hebc4:	data_out=16'ha00;
17'hebc5:	data_out=16'h89fb;
17'hebc6:	data_out=16'h8a00;
17'hebc7:	data_out=16'h9e5;
17'hebc8:	data_out=16'h80f;
17'hebc9:	data_out=16'h89f7;
17'hebca:	data_out=16'h9f6;
17'hebcb:	data_out=16'ha00;
17'hebcc:	data_out=16'h8b0;
17'hebcd:	data_out=16'h142;
17'hebce:	data_out=16'h9ff;
17'hebcf:	data_out=16'h8e9;
17'hebd0:	data_out=16'h89f5;
17'hebd1:	data_out=16'h89e5;
17'hebd2:	data_out=16'h9ed;
17'hebd3:	data_out=16'h9fe;
17'hebd4:	data_out=16'h89ee;
17'hebd5:	data_out=16'h89d6;
17'hebd6:	data_out=16'h89e6;
17'hebd7:	data_out=16'h89f2;
17'hebd8:	data_out=16'h89f2;
17'hebd9:	data_out=16'h89c5;
17'hebda:	data_out=16'h89ef;
17'hebdb:	data_out=16'ha00;
17'hebdc:	data_out=16'h800d;
17'hebdd:	data_out=16'h8917;
17'hebde:	data_out=16'h86a9;
17'hebdf:	data_out=16'h8979;
17'hebe0:	data_out=16'h57b;
17'hebe1:	data_out=16'h9fc;
17'hebe2:	data_out=16'h8180;
17'hebe3:	data_out=16'h89fa;
17'hebe4:	data_out=16'h9cf;
17'hebe5:	data_out=16'h9d0;
17'hebe6:	data_out=16'ha00;
17'hebe7:	data_out=16'h9ff;
17'hebe8:	data_out=16'h89f5;
17'hebe9:	data_out=16'h96f;
17'hebea:	data_out=16'h89ae;
17'hebeb:	data_out=16'h81f5;
17'hebec:	data_out=16'h89e3;
17'hebed:	data_out=16'h89fc;
17'hebee:	data_out=16'h89ae;
17'hebef:	data_out=16'h8091;
17'hebf0:	data_out=16'h89b5;
17'hebf1:	data_out=16'h825a;
17'hebf2:	data_out=16'h89e7;
17'hebf3:	data_out=16'h883f;
17'hebf4:	data_out=16'h89f8;
17'hebf5:	data_out=16'h89ce;
17'hebf6:	data_out=16'ha00;
17'hebf7:	data_out=16'h8707;
17'hebf8:	data_out=16'h89df;
17'hebf9:	data_out=16'h81c3;
17'hebfa:	data_out=16'h89f0;
17'hebfb:	data_out=16'h89f6;
17'hebfc:	data_out=16'h89fc;
17'hebfd:	data_out=16'h173;
17'hebfe:	data_out=16'h8a00;
17'hebff:	data_out=16'h8a00;
17'hec00:	data_out=16'h9e5;
17'hec01:	data_out=16'h9f4;
17'hec02:	data_out=16'h89f0;
17'hec03:	data_out=16'h89f2;
17'hec04:	data_out=16'ha00;
17'hec05:	data_out=16'h902;
17'hec06:	data_out=16'h89f0;
17'hec07:	data_out=16'h4ae;
17'hec08:	data_out=16'h89f4;
17'hec09:	data_out=16'h970;
17'hec0a:	data_out=16'h9ff;
17'hec0b:	data_out=16'h9fa;
17'hec0c:	data_out=16'h830d;
17'hec0d:	data_out=16'h8a00;
17'hec0e:	data_out=16'h84ea;
17'hec0f:	data_out=16'h89e8;
17'hec10:	data_out=16'h80c;
17'hec11:	data_out=16'h9f1;
17'hec12:	data_out=16'h89f9;
17'hec13:	data_out=16'h89f3;
17'hec14:	data_out=16'h89f4;
17'hec15:	data_out=16'h516;
17'hec16:	data_out=16'h89f6;
17'hec17:	data_out=16'h89e8;
17'hec18:	data_out=16'h8a00;
17'hec19:	data_out=16'ha00;
17'hec1a:	data_out=16'ha00;
17'hec1b:	data_out=16'h89f8;
17'hec1c:	data_out=16'h8504;
17'hec1d:	data_out=16'h9f2;
17'hec1e:	data_out=16'h89f9;
17'hec1f:	data_out=16'h87bc;
17'hec20:	data_out=16'h9ee;
17'hec21:	data_out=16'h84bc;
17'hec22:	data_out=16'h962;
17'hec23:	data_out=16'h81c3;
17'hec24:	data_out=16'h81b1;
17'hec25:	data_out=16'h8ce;
17'hec26:	data_out=16'h89f6;
17'hec27:	data_out=16'h9f3;
17'hec28:	data_out=16'h8470;
17'hec29:	data_out=16'h89f8;
17'hec2a:	data_out=16'h89c0;
17'hec2b:	data_out=16'ha00;
17'hec2c:	data_out=16'h8545;
17'hec2d:	data_out=16'h83f4;
17'hec2e:	data_out=16'h89e0;
17'hec2f:	data_out=16'h7f8;
17'hec30:	data_out=16'h8245;
17'hec31:	data_out=16'h9eb;
17'hec32:	data_out=16'h4ae;
17'hec33:	data_out=16'h89fb;
17'hec34:	data_out=16'h9de;
17'hec35:	data_out=16'h9f3;
17'hec36:	data_out=16'h89f2;
17'hec37:	data_out=16'h89ec;
17'hec38:	data_out=16'h9e1;
17'hec39:	data_out=16'h8a00;
17'hec3a:	data_out=16'h939;
17'hec3b:	data_out=16'h9f7;
17'hec3c:	data_out=16'h89e1;
17'hec3d:	data_out=16'h9dc;
17'hec3e:	data_out=16'h8475;
17'hec3f:	data_out=16'h8f3;
17'hec40:	data_out=16'ha00;
17'hec41:	data_out=16'h89fe;
17'hec42:	data_out=16'h9fc;
17'hec43:	data_out=16'h894a;
17'hec44:	data_out=16'h9f5;
17'hec45:	data_out=16'h4de;
17'hec46:	data_out=16'h8a00;
17'hec47:	data_out=16'h9e9;
17'hec48:	data_out=16'hc4;
17'hec49:	data_out=16'h8ff;
17'hec4a:	data_out=16'h9f4;
17'hec4b:	data_out=16'h9fe;
17'hec4c:	data_out=16'h996;
17'hec4d:	data_out=16'h957;
17'hec4e:	data_out=16'h80d5;
17'hec4f:	data_out=16'h9b1;
17'hec50:	data_out=16'h85b3;
17'hec51:	data_out=16'h89f4;
17'hec52:	data_out=16'h79b;
17'hec53:	data_out=16'h9fa;
17'hec54:	data_out=16'h9f1;
17'hec55:	data_out=16'h89ef;
17'hec56:	data_out=16'h89ff;
17'hec57:	data_out=16'h89fe;
17'hec58:	data_out=16'h89f9;
17'hec59:	data_out=16'h9fe;
17'hec5a:	data_out=16'h89ef;
17'hec5b:	data_out=16'ha00;
17'hec5c:	data_out=16'h467;
17'hec5d:	data_out=16'h8257;
17'hec5e:	data_out=16'h825;
17'hec5f:	data_out=16'h81ae;
17'hec60:	data_out=16'h89fd;
17'hec61:	data_out=16'ha00;
17'hec62:	data_out=16'h89e6;
17'hec63:	data_out=16'h89f4;
17'hec64:	data_out=16'h9eb;
17'hec65:	data_out=16'h9f4;
17'hec66:	data_out=16'h9fe;
17'hec67:	data_out=16'h87d;
17'hec68:	data_out=16'h8466;
17'hec69:	data_out=16'h898e;
17'hec6a:	data_out=16'h8518;
17'hec6b:	data_out=16'h9f8;
17'hec6c:	data_out=16'h320;
17'hec6d:	data_out=16'h89f5;
17'hec6e:	data_out=16'h851a;
17'hec6f:	data_out=16'h85da;
17'hec70:	data_out=16'h84d9;
17'hec71:	data_out=16'h89e6;
17'hec72:	data_out=16'ha00;
17'hec73:	data_out=16'ha00;
17'hec74:	data_out=16'h85cc;
17'hec75:	data_out=16'h89dc;
17'hec76:	data_out=16'ha00;
17'hec77:	data_out=16'h88cd;
17'hec78:	data_out=16'h89e1;
17'hec79:	data_out=16'h875c;
17'hec7a:	data_out=16'h89f2;
17'hec7b:	data_out=16'h8478;
17'hec7c:	data_out=16'h872e;
17'hec7d:	data_out=16'h391;
17'hec7e:	data_out=16'h248;
17'hec7f:	data_out=16'h4ff;
17'hec80:	data_out=16'ha00;
17'hec81:	data_out=16'ha00;
17'hec82:	data_out=16'h8a00;
17'hec83:	data_out=16'h640;
17'hec84:	data_out=16'ha00;
17'hec85:	data_out=16'ha00;
17'hec86:	data_out=16'ha00;
17'hec87:	data_out=16'h89a9;
17'hec88:	data_out=16'h8a00;
17'hec89:	data_out=16'ha00;
17'hec8a:	data_out=16'ha00;
17'hec8b:	data_out=16'h860b;
17'hec8c:	data_out=16'h8a00;
17'hec8d:	data_out=16'h8a00;
17'hec8e:	data_out=16'h830c;
17'hec8f:	data_out=16'h89ff;
17'hec90:	data_out=16'ha00;
17'hec91:	data_out=16'ha00;
17'hec92:	data_out=16'h8a00;
17'hec93:	data_out=16'h80cc;
17'hec94:	data_out=16'h84b6;
17'hec95:	data_out=16'ha00;
17'hec96:	data_out=16'h828f;
17'hec97:	data_out=16'h89f9;
17'hec98:	data_out=16'h85bc;
17'hec99:	data_out=16'ha00;
17'hec9a:	data_out=16'ha00;
17'hec9b:	data_out=16'h8a00;
17'hec9c:	data_out=16'h90f;
17'hec9d:	data_out=16'ha00;
17'hec9e:	data_out=16'h8229;
17'hec9f:	data_out=16'ha00;
17'heca0:	data_out=16'ha00;
17'heca1:	data_out=16'h8331;
17'heca2:	data_out=16'ha00;
17'heca3:	data_out=16'h8a00;
17'heca4:	data_out=16'h8a00;
17'heca5:	data_out=16'ha00;
17'heca6:	data_out=16'h8a00;
17'heca7:	data_out=16'ha00;
17'heca8:	data_out=16'h8360;
17'heca9:	data_out=16'h8a00;
17'hecaa:	data_out=16'h89f9;
17'hecab:	data_out=16'ha00;
17'hecac:	data_out=16'h7f8;
17'hecad:	data_out=16'h53;
17'hecae:	data_out=16'h89f9;
17'hecaf:	data_out=16'ha00;
17'hecb0:	data_out=16'h8a00;
17'hecb1:	data_out=16'ha00;
17'hecb2:	data_out=16'h8492;
17'hecb3:	data_out=16'ha00;
17'hecb4:	data_out=16'ha00;
17'hecb5:	data_out=16'ha00;
17'hecb6:	data_out=16'h89c6;
17'hecb7:	data_out=16'h8a00;
17'hecb8:	data_out=16'ha00;
17'hecb9:	data_out=16'ha00;
17'hecba:	data_out=16'ha00;
17'hecbb:	data_out=16'h1f7;
17'hecbc:	data_out=16'h89f2;
17'hecbd:	data_out=16'ha00;
17'hecbe:	data_out=16'h8364;
17'hecbf:	data_out=16'ha00;
17'hecc0:	data_out=16'ha00;
17'hecc1:	data_out=16'h8a00;
17'hecc2:	data_out=16'h8426;
17'hecc3:	data_out=16'ha00;
17'hecc4:	data_out=16'ha00;
17'hecc5:	data_out=16'ha00;
17'hecc6:	data_out=16'h8a00;
17'hecc7:	data_out=16'ha00;
17'hecc8:	data_out=16'h4e1;
17'hecc9:	data_out=16'ha00;
17'hecca:	data_out=16'h83bb;
17'heccb:	data_out=16'h8943;
17'heccc:	data_out=16'h49b;
17'heccd:	data_out=16'ha00;
17'hecce:	data_out=16'h8877;
17'heccf:	data_out=16'h9e7;
17'hecd0:	data_out=16'ha00;
17'hecd1:	data_out=16'h8a00;
17'hecd2:	data_out=16'h8718;
17'hecd3:	data_out=16'ha00;
17'hecd4:	data_out=16'ha00;
17'hecd5:	data_out=16'h89fe;
17'hecd6:	data_out=16'h9bf;
17'hecd7:	data_out=16'ha00;
17'hecd8:	data_out=16'h8a00;
17'hecd9:	data_out=16'ha00;
17'hecda:	data_out=16'h8a00;
17'hecdb:	data_out=16'ha00;
17'hecdc:	data_out=16'h77f;
17'hecdd:	data_out=16'h667;
17'hecde:	data_out=16'ha00;
17'hecdf:	data_out=16'h71d;
17'hece0:	data_out=16'h8a00;
17'hece1:	data_out=16'ha00;
17'hece2:	data_out=16'h89f5;
17'hece3:	data_out=16'h994;
17'hece4:	data_out=16'ha00;
17'hece5:	data_out=16'ha00;
17'hece6:	data_out=16'ha00;
17'hece7:	data_out=16'ha00;
17'hece8:	data_out=16'h833a;
17'hece9:	data_out=16'h8a00;
17'hecea:	data_out=16'h82e4;
17'heceb:	data_out=16'ha00;
17'hecec:	data_out=16'h2bc;
17'heced:	data_out=16'ha00;
17'hecee:	data_out=16'h82e6;
17'hecef:	data_out=16'h8de;
17'hecf0:	data_out=16'h8306;
17'hecf1:	data_out=16'h8a00;
17'hecf2:	data_out=16'ha00;
17'hecf3:	data_out=16'ha00;
17'hecf4:	data_out=16'h8a00;
17'hecf5:	data_out=16'h89fe;
17'hecf6:	data_out=16'ha00;
17'hecf7:	data_out=16'ha00;
17'hecf8:	data_out=16'h7ab;
17'hecf9:	data_out=16'h8934;
17'hecfa:	data_out=16'h80ce;
17'hecfb:	data_out=16'h8368;
17'hecfc:	data_out=16'h80c8;
17'hecfd:	data_out=16'ha00;
17'hecfe:	data_out=16'ha00;
17'hecff:	data_out=16'ha00;
17'hed00:	data_out=16'ha00;
17'hed01:	data_out=16'ha00;
17'hed02:	data_out=16'h8a00;
17'hed03:	data_out=16'h68f;
17'hed04:	data_out=16'ha00;
17'hed05:	data_out=16'h998;
17'hed06:	data_out=16'h13e;
17'hed07:	data_out=16'h81f8;
17'hed08:	data_out=16'h89ff;
17'hed09:	data_out=16'ha00;
17'hed0a:	data_out=16'ha00;
17'hed0b:	data_out=16'h8864;
17'hed0c:	data_out=16'h8a00;
17'hed0d:	data_out=16'h8a00;
17'hed0e:	data_out=16'h823c;
17'hed0f:	data_out=16'h8a00;
17'hed10:	data_out=16'ha00;
17'hed11:	data_out=16'ha00;
17'hed12:	data_out=16'h89b1;
17'hed13:	data_out=16'h840d;
17'hed14:	data_out=16'h457;
17'hed15:	data_out=16'h7d9;
17'hed16:	data_out=16'h840e;
17'hed17:	data_out=16'h8610;
17'hed18:	data_out=16'h811f;
17'hed19:	data_out=16'ha00;
17'hed1a:	data_out=16'ha00;
17'hed1b:	data_out=16'h87f7;
17'hed1c:	data_out=16'h97b;
17'hed1d:	data_out=16'ha00;
17'hed1e:	data_out=16'h294;
17'hed1f:	data_out=16'h9b8;
17'hed20:	data_out=16'ha00;
17'hed21:	data_out=16'h8253;
17'hed22:	data_out=16'ha00;
17'hed23:	data_out=16'h8a00;
17'hed24:	data_out=16'h8a00;
17'hed25:	data_out=16'h218;
17'hed26:	data_out=16'h8a00;
17'hed27:	data_out=16'ha00;
17'hed28:	data_out=16'h8270;
17'hed29:	data_out=16'h8090;
17'hed2a:	data_out=16'h8a00;
17'hed2b:	data_out=16'ha00;
17'hed2c:	data_out=16'h88;
17'hed2d:	data_out=16'h852d;
17'hed2e:	data_out=16'h8a00;
17'hed2f:	data_out=16'ha00;
17'hed30:	data_out=16'h8a00;
17'hed31:	data_out=16'ha00;
17'hed32:	data_out=16'h8a00;
17'hed33:	data_out=16'ha00;
17'hed34:	data_out=16'ha00;
17'hed35:	data_out=16'h82a5;
17'hed36:	data_out=16'h8825;
17'hed37:	data_out=16'h8a00;
17'hed38:	data_out=16'ha00;
17'hed39:	data_out=16'ha00;
17'hed3a:	data_out=16'ha00;
17'hed3b:	data_out=16'h394;
17'hed3c:	data_out=16'h8a00;
17'hed3d:	data_out=16'ha00;
17'hed3e:	data_out=16'h8272;
17'hed3f:	data_out=16'h99f;
17'hed40:	data_out=16'ha00;
17'hed41:	data_out=16'h8a00;
17'hed42:	data_out=16'h8a00;
17'hed43:	data_out=16'h66;
17'hed44:	data_out=16'ha00;
17'hed45:	data_out=16'h79d;
17'hed46:	data_out=16'h8a00;
17'hed47:	data_out=16'h4b4;
17'hed48:	data_out=16'h80db;
17'hed49:	data_out=16'h360;
17'hed4a:	data_out=16'h87fb;
17'hed4b:	data_out=16'h8a00;
17'hed4c:	data_out=16'h85e1;
17'hed4d:	data_out=16'ha00;
17'hed4e:	data_out=16'h8a00;
17'hed4f:	data_out=16'h8216;
17'hed50:	data_out=16'h7f0;
17'hed51:	data_out=16'h8a00;
17'hed52:	data_out=16'h876a;
17'hed53:	data_out=16'ha00;
17'hed54:	data_out=16'ha00;
17'hed55:	data_out=16'h8a00;
17'hed56:	data_out=16'h856;
17'hed57:	data_out=16'ha00;
17'hed58:	data_out=16'h8a00;
17'hed59:	data_out=16'ha00;
17'hed5a:	data_out=16'h8a00;
17'hed5b:	data_out=16'ha00;
17'hed5c:	data_out=16'h8f2;
17'hed5d:	data_out=16'h82d0;
17'hed5e:	data_out=16'ha00;
17'hed5f:	data_out=16'h318;
17'hed60:	data_out=16'h8a00;
17'hed61:	data_out=16'ha00;
17'hed62:	data_out=16'h8a00;
17'hed63:	data_out=16'ha00;
17'hed64:	data_out=16'ha00;
17'hed65:	data_out=16'ha00;
17'hed66:	data_out=16'ha00;
17'hed67:	data_out=16'h3a9;
17'hed68:	data_out=16'h825b;
17'hed69:	data_out=16'h8a00;
17'hed6a:	data_out=16'h822d;
17'hed6b:	data_out=16'ha00;
17'hed6c:	data_out=16'h1c;
17'hed6d:	data_out=16'ha00;
17'hed6e:	data_out=16'h822e;
17'hed6f:	data_out=16'h810e;
17'hed70:	data_out=16'h8239;
17'hed71:	data_out=16'h8a00;
17'hed72:	data_out=16'ha00;
17'hed73:	data_out=16'ha00;
17'hed74:	data_out=16'h8a00;
17'hed75:	data_out=16'h8a00;
17'hed76:	data_out=16'ha00;
17'hed77:	data_out=16'h649;
17'hed78:	data_out=16'h808d;
17'hed79:	data_out=16'h8a00;
17'hed7a:	data_out=16'h616;
17'hed7b:	data_out=16'h8274;
17'hed7c:	data_out=16'he3;
17'hed7d:	data_out=16'h3f1;
17'hed7e:	data_out=16'ha00;
17'hed7f:	data_out=16'ha00;
17'hed80:	data_out=16'h4e6;
17'hed81:	data_out=16'h254;
17'hed82:	data_out=16'h8339;
17'hed83:	data_out=16'h19;
17'hed84:	data_out=16'h1d;
17'hed85:	data_out=16'h99;
17'hed86:	data_out=16'h8133;
17'hed87:	data_out=16'h80b4;
17'hed88:	data_out=16'h8141;
17'hed89:	data_out=16'h23a;
17'hed8a:	data_out=16'h12e;
17'hed8b:	data_out=16'h81bd;
17'hed8c:	data_out=16'h851b;
17'hed8d:	data_out=16'h8116;
17'hed8e:	data_out=16'h8055;
17'hed8f:	data_out=16'h81ed;
17'hed90:	data_out=16'hc3;
17'hed91:	data_out=16'h1fc;
17'hed92:	data_out=16'h828f;
17'hed93:	data_out=16'h801c;
17'hed94:	data_out=16'h8073;
17'hed95:	data_out=16'h1a4;
17'hed96:	data_out=16'h4f;
17'hed97:	data_out=16'h81a3;
17'hed98:	data_out=16'h805d;
17'hed99:	data_out=16'h1ff;
17'hed9a:	data_out=16'h8079;
17'hed9b:	data_out=16'h13;
17'hed9c:	data_out=16'h430;
17'hed9d:	data_out=16'h1f3;
17'hed9e:	data_out=16'hbe;
17'hed9f:	data_out=16'h80c2;
17'heda0:	data_out=16'h4f5;
17'heda1:	data_out=16'h8058;
17'heda2:	data_out=16'h198;
17'heda3:	data_out=16'h8271;
17'heda4:	data_out=16'h826f;
17'heda5:	data_out=16'h80ba;
17'heda6:	data_out=16'h807e;
17'heda7:	data_out=16'h20f;
17'heda8:	data_out=16'h806e;
17'heda9:	data_out=16'h6c;
17'hedaa:	data_out=16'h82ca;
17'hedab:	data_out=16'h6c2;
17'hedac:	data_out=16'h8024;
17'hedad:	data_out=16'h80d7;
17'hedae:	data_out=16'h8308;
17'hedaf:	data_out=16'h212;
17'hedb0:	data_out=16'h81f0;
17'hedb1:	data_out=16'h4ed;
17'hedb2:	data_out=16'h81b8;
17'hedb3:	data_out=16'hb8;
17'hedb4:	data_out=16'h4d1;
17'hedb5:	data_out=16'h8164;
17'hedb6:	data_out=16'h81c6;
17'hedb7:	data_out=16'h833a;
17'hedb8:	data_out=16'h6db;
17'hedb9:	data_out=16'h1ff;
17'hedba:	data_out=16'h11;
17'hedbb:	data_out=16'h1f8;
17'hedbc:	data_out=16'h82fc;
17'hedbd:	data_out=16'h6c3;
17'hedbe:	data_out=16'h8061;
17'hedbf:	data_out=16'hac;
17'hedc0:	data_out=16'h804b;
17'hedc1:	data_out=16'h82c9;
17'hedc2:	data_out=16'h8374;
17'hedc3:	data_out=16'h811e;
17'hedc4:	data_out=16'h1a7;
17'hedc5:	data_out=16'h19d;
17'hedc6:	data_out=16'h8119;
17'hedc7:	data_out=16'h8160;
17'hedc8:	data_out=16'h81d4;
17'hedc9:	data_out=16'h8064;
17'hedca:	data_out=16'h8285;
17'hedcb:	data_out=16'h84fa;
17'hedcc:	data_out=16'h8296;
17'hedcd:	data_out=16'h2bd;
17'hedce:	data_out=16'h81a2;
17'hedcf:	data_out=16'h81ba;
17'hedd0:	data_out=16'h8078;
17'hedd1:	data_out=16'h80fc;
17'hedd2:	data_out=16'h81d6;
17'hedd3:	data_out=16'h18d;
17'hedd4:	data_out=16'h2ad;
17'hedd5:	data_out=16'h8328;
17'hedd6:	data_out=16'h8092;
17'hedd7:	data_out=16'h8031;
17'hedd8:	data_out=16'h837e;
17'hedd9:	data_out=16'h8044;
17'hedda:	data_out=16'h825b;
17'heddb:	data_out=16'h199;
17'heddc:	data_out=16'hde;
17'heddd:	data_out=16'h808b;
17'hedde:	data_out=16'h119;
17'heddf:	data_out=16'h54;
17'hede0:	data_out=16'h80f1;
17'hede1:	data_out=16'h2ca;
17'hede2:	data_out=16'h833b;
17'hede3:	data_out=16'h50;
17'hede4:	data_out=16'h58d;
17'hede5:	data_out=16'he8;
17'hede6:	data_out=16'h174;
17'hede7:	data_out=16'h80c6;
17'hede8:	data_out=16'h8064;
17'hede9:	data_out=16'h8355;
17'hedea:	data_out=16'h8054;
17'hedeb:	data_out=16'h2ce;
17'hedec:	data_out=16'h806d;
17'heded:	data_out=16'hca;
17'hedee:	data_out=16'h8064;
17'hedef:	data_out=16'h806a;
17'hedf0:	data_out=16'h805e;
17'hedf1:	data_out=16'h833a;
17'hedf2:	data_out=16'h1a5;
17'hedf3:	data_out=16'h2de;
17'hedf4:	data_out=16'h8206;
17'hedf5:	data_out=16'h8207;
17'hedf6:	data_out=16'h354;
17'hedf7:	data_out=16'h80f9;
17'hedf8:	data_out=16'h9e;
17'hedf9:	data_out=16'h83df;
17'hedfa:	data_out=16'h8044;
17'hedfb:	data_out=16'h8061;
17'hedfc:	data_out=16'h80de;
17'hedfd:	data_out=16'h80e9;
17'hedfe:	data_out=16'h24f;
17'hedff:	data_out=16'h8033;
17'hee00:	data_out=16'h4;
17'hee01:	data_out=16'h8008;
17'hee02:	data_out=16'h3;
17'hee03:	data_out=16'h8;
17'hee04:	data_out=16'h5;
17'hee05:	data_out=16'h2;
17'hee06:	data_out=16'h8000;
17'hee07:	data_out=16'h8007;
17'hee08:	data_out=16'h4;
17'hee09:	data_out=16'h8003;
17'hee0a:	data_out=16'h1;
17'hee0b:	data_out=16'h8001;
17'hee0c:	data_out=16'h8000;
17'hee0d:	data_out=16'h1;
17'hee0e:	data_out=16'h5;
17'hee0f:	data_out=16'h5;
17'hee10:	data_out=16'h8005;
17'hee11:	data_out=16'h8009;
17'hee12:	data_out=16'h9;
17'hee13:	data_out=16'h0;
17'hee14:	data_out=16'h5;
17'hee15:	data_out=16'h8006;
17'hee16:	data_out=16'h8002;
17'hee17:	data_out=16'h8002;
17'hee18:	data_out=16'h2;
17'hee19:	data_out=16'h8004;
17'hee1a:	data_out=16'h8007;
17'hee1b:	data_out=16'h8008;
17'hee1c:	data_out=16'h8008;
17'hee1d:	data_out=16'h8003;
17'hee1e:	data_out=16'h3;
17'hee1f:	data_out=16'h5;
17'hee20:	data_out=16'h8002;
17'hee21:	data_out=16'h8003;
17'hee22:	data_out=16'h4;
17'hee23:	data_out=16'h8006;
17'hee24:	data_out=16'h8;
17'hee25:	data_out=16'h8006;
17'hee26:	data_out=16'h8004;
17'hee27:	data_out=16'h3;
17'hee28:	data_out=16'h1;
17'hee29:	data_out=16'h6;
17'hee2a:	data_out=16'h8008;
17'hee2b:	data_out=16'h8009;
17'hee2c:	data_out=16'h8002;
17'hee2d:	data_out=16'h6;
17'hee2e:	data_out=16'h5;
17'hee2f:	data_out=16'h3;
17'hee30:	data_out=16'h6;
17'hee31:	data_out=16'h5;
17'hee32:	data_out=16'h8006;
17'hee33:	data_out=16'h3;
17'hee34:	data_out=16'h8;
17'hee35:	data_out=16'h1;
17'hee36:	data_out=16'h8009;
17'hee37:	data_out=16'h1;
17'hee38:	data_out=16'h6;
17'hee39:	data_out=16'h8007;
17'hee3a:	data_out=16'h2;
17'hee3b:	data_out=16'h6;
17'hee3c:	data_out=16'h8001;
17'hee3d:	data_out=16'h8004;
17'hee3e:	data_out=16'h2;
17'hee3f:	data_out=16'h6;
17'hee40:	data_out=16'h2;
17'hee41:	data_out=16'h8003;
17'hee42:	data_out=16'h9;
17'hee43:	data_out=16'h0;
17'hee44:	data_out=16'h0;
17'hee45:	data_out=16'h8004;
17'hee46:	data_out=16'h8006;
17'hee47:	data_out=16'h8008;
17'hee48:	data_out=16'h8007;
17'hee49:	data_out=16'h8005;
17'hee4a:	data_out=16'h8008;
17'hee4b:	data_out=16'h1;
17'hee4c:	data_out=16'h8008;
17'hee4d:	data_out=16'h6;
17'hee4e:	data_out=16'h8005;
17'hee4f:	data_out=16'h7;
17'hee50:	data_out=16'h1;
17'hee51:	data_out=16'h8002;
17'hee52:	data_out=16'h1;
17'hee53:	data_out=16'h0;
17'hee54:	data_out=16'h8;
17'hee55:	data_out=16'h1;
17'hee56:	data_out=16'h8008;
17'hee57:	data_out=16'h4;
17'hee58:	data_out=16'h4;
17'hee59:	data_out=16'h3;
17'hee5a:	data_out=16'h1;
17'hee5b:	data_out=16'h8006;
17'hee5c:	data_out=16'h8;
17'hee5d:	data_out=16'h8006;
17'hee5e:	data_out=16'h9;
17'hee5f:	data_out=16'h1;
17'hee60:	data_out=16'h1;
17'hee61:	data_out=16'h9;
17'hee62:	data_out=16'h8008;
17'hee63:	data_out=16'h8008;
17'hee64:	data_out=16'h8004;
17'hee65:	data_out=16'h8005;
17'hee66:	data_out=16'h8007;
17'hee67:	data_out=16'h8001;
17'hee68:	data_out=16'h8001;
17'hee69:	data_out=16'h8006;
17'hee6a:	data_out=16'h9;
17'hee6b:	data_out=16'h8000;
17'hee6c:	data_out=16'h8009;
17'hee6d:	data_out=16'h8006;
17'hee6e:	data_out=16'h8002;
17'hee6f:	data_out=16'h2;
17'hee70:	data_out=16'h1;
17'hee71:	data_out=16'h9;
17'hee72:	data_out=16'h8007;
17'hee73:	data_out=16'h8000;
17'hee74:	data_out=16'h1;
17'hee75:	data_out=16'h8006;
17'hee76:	data_out=16'h8005;
17'hee77:	data_out=16'h8005;
17'hee78:	data_out=16'h6;
17'hee79:	data_out=16'h5;
17'hee7a:	data_out=16'h8002;
17'hee7b:	data_out=16'h5;
17'hee7c:	data_out=16'h9;
17'hee7d:	data_out=16'h8002;
17'hee7e:	data_out=16'h8003;
17'hee7f:	data_out=16'h0;
17'hee80:	data_out=16'h8054;
17'hee81:	data_out=16'h37;
17'hee82:	data_out=16'h2;
17'hee83:	data_out=16'h800b;
17'hee84:	data_out=16'h803b;
17'hee85:	data_out=16'h87;
17'hee86:	data_out=16'h5d;
17'hee87:	data_out=16'h8017;
17'hee88:	data_out=16'h56;
17'hee89:	data_out=16'h8065;
17'hee8a:	data_out=16'h8019;
17'hee8b:	data_out=16'had;
17'hee8c:	data_out=16'h5e;
17'hee8d:	data_out=16'h2;
17'hee8e:	data_out=16'h8005;
17'hee8f:	data_out=16'h25;
17'hee90:	data_out=16'h806d;
17'hee91:	data_out=16'h3;
17'hee92:	data_out=16'h15;
17'hee93:	data_out=16'h8037;
17'hee94:	data_out=16'h55;
17'hee95:	data_out=16'h804c;
17'hee96:	data_out=16'h803c;
17'hee97:	data_out=16'h72;
17'hee98:	data_out=16'h8029;
17'hee99:	data_out=16'h8014;
17'hee9a:	data_out=16'h802e;
17'hee9b:	data_out=16'h9d;
17'hee9c:	data_out=16'ha9;
17'hee9d:	data_out=16'h50;
17'hee9e:	data_out=16'h7d;
17'hee9f:	data_out=16'h3f;
17'heea0:	data_out=16'h82;
17'heea1:	data_out=16'h8006;
17'heea2:	data_out=16'h803f;
17'heea3:	data_out=16'h805e;
17'heea4:	data_out=16'h806a;
17'heea5:	data_out=16'h804a;
17'heea6:	data_out=16'h8016;
17'heea7:	data_out=16'h88;
17'heea8:	data_out=16'h2;
17'heea9:	data_out=16'h801a;
17'heeaa:	data_out=16'h8032;
17'heeab:	data_out=16'h42;
17'heeac:	data_out=16'h8004;
17'heead:	data_out=16'h80b0;
17'heeae:	data_out=16'h8013;
17'heeaf:	data_out=16'h5f;
17'heeb0:	data_out=16'h23;
17'heeb1:	data_out=16'h2c;
17'heeb2:	data_out=16'h18;
17'heeb3:	data_out=16'h46;
17'heeb4:	data_out=16'h8005;
17'heeb5:	data_out=16'h7b;
17'heeb6:	data_out=16'h6d;
17'heeb7:	data_out=16'h17;
17'heeb8:	data_out=16'h58;
17'heeb9:	data_out=16'h42;
17'heeba:	data_out=16'h80a5;
17'heebb:	data_out=16'h37;
17'heebc:	data_out=16'h50;
17'heebd:	data_out=16'h805e;
17'heebe:	data_out=16'h4;
17'heebf:	data_out=16'h3e;
17'heec0:	data_out=16'h8096;
17'heec1:	data_out=16'hb9;
17'heec2:	data_out=16'h8048;
17'heec3:	data_out=16'h6a;
17'heec4:	data_out=16'h800f;
17'heec5:	data_out=16'h8051;
17'heec6:	data_out=16'h55;
17'heec7:	data_out=16'h809e;
17'heec8:	data_out=16'h800f;
17'heec9:	data_out=16'h8051;
17'heeca:	data_out=16'h8025;
17'heecb:	data_out=16'h1f;
17'heecc:	data_out=16'h8066;
17'heecd:	data_out=16'h803b;
17'heece:	data_out=16'h8018;
17'heecf:	data_out=16'h8077;
17'heed0:	data_out=16'h8091;
17'heed1:	data_out=16'h46;
17'heed2:	data_out=16'h8073;
17'heed3:	data_out=16'hde;
17'heed4:	data_out=16'h6d;
17'heed5:	data_out=16'h8b;
17'heed6:	data_out=16'h8062;
17'heed7:	data_out=16'h80ae;
17'heed8:	data_out=16'h3b;
17'heed9:	data_out=16'h80ab;
17'heeda:	data_out=16'h9b;
17'heedb:	data_out=16'hc1;
17'heedc:	data_out=16'h8c;
17'heedd:	data_out=16'h8046;
17'heede:	data_out=16'h5e;
17'heedf:	data_out=16'h8013;
17'heee0:	data_out=16'h8059;
17'heee1:	data_out=16'h35;
17'heee2:	data_out=16'hf6;
17'heee3:	data_out=16'h3f;
17'heee4:	data_out=16'h8019;
17'heee5:	data_out=16'h800e;
17'heee6:	data_out=16'h8003;
17'heee7:	data_out=16'h8027;
17'heee8:	data_out=16'h8005;
17'heee9:	data_out=16'h3c;
17'heeea:	data_out=16'h800b;
17'heeeb:	data_out=16'h3;
17'heeec:	data_out=16'h80cb;
17'heeed:	data_out=16'h49;
17'heeee:	data_out=16'h8008;
17'heeef:	data_out=16'h1d;
17'heef0:	data_out=16'h800c;
17'heef1:	data_out=16'h3;
17'heef2:	data_out=16'h8055;
17'heef3:	data_out=16'h4;
17'heef4:	data_out=16'h22;
17'heef5:	data_out=16'hd6;
17'heef6:	data_out=16'h41;
17'heef7:	data_out=16'h80ad;
17'heef8:	data_out=16'h4f;
17'heef9:	data_out=16'h8002;
17'heefa:	data_out=16'h4c;
17'heefb:	data_out=16'h8;
17'heefc:	data_out=16'h2d;
17'heefd:	data_out=16'hc2;
17'heefe:	data_out=16'h8046;
17'heeff:	data_out=16'h80a1;
17'hef00:	data_out=16'h8896;
17'hef01:	data_out=16'h82e1;
17'hef02:	data_out=16'h8367;
17'hef03:	data_out=16'h8564;
17'hef04:	data_out=16'h80aa;
17'hef05:	data_out=16'h3fd;
17'hef06:	data_out=16'h36f;
17'hef07:	data_out=16'h8388;
17'hef08:	data_out=16'h877a;
17'hef09:	data_out=16'h8604;
17'hef0a:	data_out=16'h861a;
17'hef0b:	data_out=16'h2b8;
17'hef0c:	data_out=16'h826b;
17'hef0d:	data_out=16'h832d;
17'hef0e:	data_out=16'h8159;
17'hef0f:	data_out=16'h8327;
17'hef10:	data_out=16'h86bb;
17'hef11:	data_out=16'hfa;
17'hef12:	data_out=16'h819b;
17'hef13:	data_out=16'h85d8;
17'hef14:	data_out=16'h1e1;
17'hef15:	data_out=16'h8363;
17'hef16:	data_out=16'h86bc;
17'hef17:	data_out=16'h191;
17'hef18:	data_out=16'h81a8;
17'hef19:	data_out=16'h3a2;
17'hef1a:	data_out=16'h8092;
17'hef1b:	data_out=16'h430;
17'hef1c:	data_out=16'h309;
17'hef1d:	data_out=16'h95;
17'hef1e:	data_out=16'h8;
17'hef1f:	data_out=16'he9;
17'hef20:	data_out=16'h515;
17'hef21:	data_out=16'h814b;
17'hef22:	data_out=16'h8560;
17'hef23:	data_out=16'h8477;
17'hef24:	data_out=16'h8478;
17'hef25:	data_out=16'h868d;
17'hef26:	data_out=16'h8a00;
17'hef27:	data_out=16'h2f9;
17'hef28:	data_out=16'h812f;
17'hef29:	data_out=16'h861c;
17'hef2a:	data_out=16'h890e;
17'hef2b:	data_out=16'h66c;
17'hef2c:	data_out=16'h85f1;
17'hef2d:	data_out=16'h8a00;
17'hef2e:	data_out=16'h84e9;
17'hef2f:	data_out=16'hf9;
17'hef30:	data_out=16'h8567;
17'hef31:	data_out=16'h147;
17'hef32:	data_out=16'h8539;
17'hef33:	data_out=16'h195;
17'hef34:	data_out=16'h1b9;
17'hef35:	data_out=16'h19a;
17'hef36:	data_out=16'h847d;
17'hef37:	data_out=16'h828b;
17'hef38:	data_out=16'h579;
17'hef39:	data_out=16'h1db;
17'hef3a:	data_out=16'h86d1;
17'hef3b:	data_out=16'h8332;
17'hef3c:	data_out=16'h84b6;
17'hef3d:	data_out=16'h8307;
17'hef3e:	data_out=16'h812f;
17'hef3f:	data_out=16'h3ce;
17'hef40:	data_out=16'h8539;
17'hef41:	data_out=16'h804b;
17'hef42:	data_out=16'h8a00;
17'hef43:	data_out=16'h34a;
17'hef44:	data_out=16'h80b8;
17'hef45:	data_out=16'h838a;
17'hef46:	data_out=16'h8460;
17'hef47:	data_out=16'h87cb;
17'hef48:	data_out=16'h57;
17'hef49:	data_out=16'h866e;
17'hef4a:	data_out=16'h83d0;
17'hef4b:	data_out=16'h8758;
17'hef4c:	data_out=16'h87cf;
17'hef4d:	data_out=16'h8525;
17'hef4e:	data_out=16'h8528;
17'hef4f:	data_out=16'h873f;
17'hef50:	data_out=16'h853c;
17'hef51:	data_out=16'h8236;
17'hef52:	data_out=16'h8672;
17'hef53:	data_out=16'h63f;
17'hef54:	data_out=16'h8049;
17'hef55:	data_out=16'h83d3;
17'hef56:	data_out=16'h8778;
17'hef57:	data_out=16'h874a;
17'hef58:	data_out=16'h8468;
17'hef59:	data_out=16'h8683;
17'hef5a:	data_out=16'h22b;
17'hef5b:	data_out=16'h3d1;
17'hef5c:	data_out=16'h51c;
17'hef5d:	data_out=16'h8717;
17'hef5e:	data_out=16'h3b;
17'hef5f:	data_out=16'h81c0;
17'hef60:	data_out=16'h8a00;
17'hef61:	data_out=16'h13d;
17'hef62:	data_out=16'h30e;
17'hef63:	data_out=16'h229;
17'hef64:	data_out=16'h301;
17'hef65:	data_out=16'h8008;
17'hef66:	data_out=16'h44a;
17'hef67:	data_out=16'h82d8;
17'hef68:	data_out=16'h8141;
17'hef69:	data_out=16'h8963;
17'hef6a:	data_out=16'h8162;
17'hef6b:	data_out=16'h16e;
17'hef6c:	data_out=16'h8a00;
17'hef6d:	data_out=16'h1ec;
17'hef6e:	data_out=16'h8162;
17'hef6f:	data_out=16'h846c;
17'hef70:	data_out=16'h815d;
17'hef71:	data_out=16'h80c8;
17'hef72:	data_out=16'h8525;
17'hef73:	data_out=16'h8122;
17'hef74:	data_out=16'h8585;
17'hef75:	data_out=16'h31b;
17'hef76:	data_out=16'h39d;
17'hef77:	data_out=16'h8823;
17'hef78:	data_out=16'h3b9;
17'hef79:	data_out=16'h85fb;
17'hef7a:	data_out=16'h241;
17'hef7b:	data_out=16'h812f;
17'hef7c:	data_out=16'h809b;
17'hef7d:	data_out=16'h67e;
17'hef7e:	data_out=16'h8590;
17'hef7f:	data_out=16'h85b0;
17'hef80:	data_out=16'h89ef;
17'hef81:	data_out=16'h804b;
17'hef82:	data_out=16'h8860;
17'hef83:	data_out=16'h8a00;
17'hef84:	data_out=16'h2d7;
17'hef85:	data_out=16'h9f9;
17'hef86:	data_out=16'h981;
17'hef87:	data_out=16'h8a00;
17'hef88:	data_out=16'h8764;
17'hef89:	data_out=16'h8a00;
17'hef8a:	data_out=16'h89fd;
17'hef8b:	data_out=16'h9be;
17'hef8c:	data_out=16'h8a00;
17'hef8d:	data_out=16'h8262;
17'hef8e:	data_out=16'h8105;
17'hef8f:	data_out=16'h89ff;
17'hef90:	data_out=16'h89e8;
17'hef91:	data_out=16'h840;
17'hef92:	data_out=16'h82a7;
17'hef93:	data_out=16'h897c;
17'hef94:	data_out=16'h9fc;
17'hef95:	data_out=16'h84fa;
17'hef96:	data_out=16'h8a00;
17'hef97:	data_out=16'h9f1;
17'hef98:	data_out=16'h81a3;
17'hef99:	data_out=16'ha00;
17'hef9a:	data_out=16'h336;
17'hef9b:	data_out=16'h9f9;
17'hef9c:	data_out=16'h9f9;
17'hef9d:	data_out=16'h9ff;
17'hef9e:	data_out=16'h8f7;
17'hef9f:	data_out=16'h70b;
17'hefa0:	data_out=16'ha00;
17'hefa1:	data_out=16'h80d0;
17'hefa2:	data_out=16'h89fd;
17'hefa3:	data_out=16'h8a00;
17'hefa4:	data_out=16'h8a00;
17'hefa5:	data_out=16'h8a00;
17'hefa6:	data_out=16'h8a00;
17'hefa7:	data_out=16'ha00;
17'hefa8:	data_out=16'h8062;
17'hefa9:	data_out=16'h8a00;
17'hefaa:	data_out=16'h8a00;
17'hefab:	data_out=16'ha00;
17'hefac:	data_out=16'h8a00;
17'hefad:	data_out=16'h8a00;
17'hefae:	data_out=16'h89f9;
17'hefaf:	data_out=16'ha00;
17'hefb0:	data_out=16'h8a00;
17'hefb1:	data_out=16'h90d;
17'hefb2:	data_out=16'h89fb;
17'hefb3:	data_out=16'ha00;
17'hefb4:	data_out=16'h1b3;
17'hefb5:	data_out=16'h6c9;
17'hefb6:	data_out=16'h849e;
17'hefb7:	data_out=16'h8776;
17'hefb8:	data_out=16'ha00;
17'hefb9:	data_out=16'ha00;
17'hefba:	data_out=16'h8a00;
17'hefbb:	data_out=16'h89d8;
17'hefbc:	data_out=16'h839d;
17'hefbd:	data_out=16'h9fd;
17'hefbe:	data_out=16'h8061;
17'hefbf:	data_out=16'h9f9;
17'hefc0:	data_out=16'h8936;
17'hefc1:	data_out=16'h96d;
17'hefc2:	data_out=16'h8a00;
17'hefc3:	data_out=16'h9f5;
17'hefc4:	data_out=16'ha00;
17'hefc5:	data_out=16'h85db;
17'hefc6:	data_out=16'h8977;
17'hefc7:	data_out=16'h8a00;
17'hefc8:	data_out=16'h424;
17'hefc9:	data_out=16'h8a00;
17'hefca:	data_out=16'h846d;
17'hefcb:	data_out=16'h8a00;
17'hefcc:	data_out=16'h8a00;
17'hefcd:	data_out=16'h87d5;
17'hefce:	data_out=16'h89a8;
17'hefcf:	data_out=16'h8a00;
17'hefd0:	data_out=16'h876b;
17'hefd1:	data_out=16'h8121;
17'hefd2:	data_out=16'h8a00;
17'hefd3:	data_out=16'ha00;
17'hefd4:	data_out=16'ha00;
17'hefd5:	data_out=16'h888d;
17'hefd6:	data_out=16'h89ff;
17'hefd7:	data_out=16'h89f6;
17'hefd8:	data_out=16'h83c2;
17'hefd9:	data_out=16'h89df;
17'hefda:	data_out=16'h9fa;
17'hefdb:	data_out=16'ha00;
17'hefdc:	data_out=16'h9f8;
17'hefdd:	data_out=16'h89f8;
17'hefde:	data_out=16'ha00;
17'hefdf:	data_out=16'h49;
17'hefe0:	data_out=16'h8a00;
17'hefe1:	data_out=16'h9f7;
17'hefe2:	data_out=16'h47e;
17'hefe3:	data_out=16'ha00;
17'hefe4:	data_out=16'ha00;
17'hefe5:	data_out=16'h41c;
17'hefe6:	data_out=16'ha00;
17'hefe7:	data_out=16'h89ea;
17'hefe8:	data_out=16'h80a8;
17'hefe9:	data_out=16'h89fc;
17'hefea:	data_out=16'h8127;
17'hefeb:	data_out=16'h9fc;
17'hefec:	data_out=16'h89f9;
17'hefed:	data_out=16'ha00;
17'hefee:	data_out=16'h8127;
17'hefef:	data_out=16'h89fb;
17'heff0:	data_out=16'h8113;
17'heff1:	data_out=16'h87b2;
17'heff2:	data_out=16'h89ec;
17'heff3:	data_out=16'h88a;
17'heff4:	data_out=16'h8a00;
17'heff5:	data_out=16'h9ef;
17'heff6:	data_out=16'h9ff;
17'heff7:	data_out=16'h8a00;
17'heff8:	data_out=16'h9fd;
17'heff9:	data_out=16'h89f6;
17'heffa:	data_out=16'h9ff;
17'heffb:	data_out=16'h8062;
17'heffc:	data_out=16'h41c;
17'heffd:	data_out=16'ha00;
17'heffe:	data_out=16'h89fd;
17'hefff:	data_out=16'h8786;
17'hf000:	data_out=16'ha00;
17'hf001:	data_out=16'h9fe;
17'hf002:	data_out=16'h8648;
17'hf003:	data_out=16'h8a00;
17'hf004:	data_out=16'ha00;
17'hf005:	data_out=16'h4b2;
17'hf006:	data_out=16'h22c;
17'hf007:	data_out=16'h89f2;
17'hf008:	data_out=16'h7c4;
17'hf009:	data_out=16'h89f8;
17'hf00a:	data_out=16'h390;
17'hf00b:	data_out=16'h9ff;
17'hf00c:	data_out=16'h89f7;
17'hf00d:	data_out=16'h8a00;
17'hf00e:	data_out=16'h852b;
17'hf00f:	data_out=16'h89f9;
17'hf010:	data_out=16'h405;
17'hf011:	data_out=16'ha00;
17'hf012:	data_out=16'h9f4;
17'hf013:	data_out=16'h83a5;
17'hf014:	data_out=16'h9f5;
17'hf015:	data_out=16'h816a;
17'hf016:	data_out=16'h8a00;
17'hf017:	data_out=16'h9dc;
17'hf018:	data_out=16'h66c;
17'hf019:	data_out=16'ha00;
17'hf01a:	data_out=16'h876e;
17'hf01b:	data_out=16'h9ec;
17'hf01c:	data_out=16'h94c;
17'hf01d:	data_out=16'h9ff;
17'hf01e:	data_out=16'h9f1;
17'hf01f:	data_out=16'h9fe;
17'hf020:	data_out=16'ha00;
17'hf021:	data_out=16'h8540;
17'hf022:	data_out=16'h89fe;
17'hf023:	data_out=16'h88ac;
17'hf024:	data_out=16'h888b;
17'hf025:	data_out=16'h8a00;
17'hf026:	data_out=16'h8a00;
17'hf027:	data_out=16'ha00;
17'hf028:	data_out=16'h84f4;
17'hf029:	data_out=16'h8a00;
17'hf02a:	data_out=16'h89f8;
17'hf02b:	data_out=16'ha00;
17'hf02c:	data_out=16'h8a00;
17'hf02d:	data_out=16'h89fa;
17'hf02e:	data_out=16'h80cc;
17'hf02f:	data_out=16'ha00;
17'hf030:	data_out=16'h8a00;
17'hf031:	data_out=16'h9fe;
17'hf032:	data_out=16'h8a00;
17'hf033:	data_out=16'ha00;
17'hf034:	data_out=16'h931;
17'hf035:	data_out=16'h9ff;
17'hf036:	data_out=16'h9fe;
17'hf037:	data_out=16'h8466;
17'hf038:	data_out=16'ha00;
17'hf039:	data_out=16'h9ff;
17'hf03a:	data_out=16'h854c;
17'hf03b:	data_out=16'h5ec;
17'hf03c:	data_out=16'hec;
17'hf03d:	data_out=16'h9fd;
17'hf03e:	data_out=16'h84f4;
17'hf03f:	data_out=16'h48f;
17'hf040:	data_out=16'h896a;
17'hf041:	data_out=16'h9e5;
17'hf042:	data_out=16'h8a00;
17'hf043:	data_out=16'h8a00;
17'hf044:	data_out=16'ha00;
17'hf045:	data_out=16'h82c5;
17'hf046:	data_out=16'h8991;
17'hf047:	data_out=16'h89ed;
17'hf048:	data_out=16'ha00;
17'hf049:	data_out=16'h8a00;
17'hf04a:	data_out=16'h3f3;
17'hf04b:	data_out=16'h89ff;
17'hf04c:	data_out=16'h8a00;
17'hf04d:	data_out=16'h89fc;
17'hf04e:	data_out=16'h8d;
17'hf04f:	data_out=16'h8a00;
17'hf050:	data_out=16'h89fd;
17'hf051:	data_out=16'h829b;
17'hf052:	data_out=16'h89fc;
17'hf053:	data_out=16'ha00;
17'hf054:	data_out=16'ha00;
17'hf055:	data_out=16'h89fe;
17'hf056:	data_out=16'h87cf;
17'hf057:	data_out=16'h89c7;
17'hf058:	data_out=16'h83df;
17'hf059:	data_out=16'h89ca;
17'hf05a:	data_out=16'h9f3;
17'hf05b:	data_out=16'ha00;
17'hf05c:	data_out=16'h9e4;
17'hf05d:	data_out=16'h89e8;
17'hf05e:	data_out=16'ha00;
17'hf05f:	data_out=16'ha00;
17'hf060:	data_out=16'h8a00;
17'hf061:	data_out=16'h68e;
17'hf062:	data_out=16'h3d7;
17'hf063:	data_out=16'ha00;
17'hf064:	data_out=16'ha00;
17'hf065:	data_out=16'h9ff;
17'hf066:	data_out=16'ha00;
17'hf067:	data_out=16'h89d4;
17'hf068:	data_out=16'h852a;
17'hf069:	data_out=16'h8290;
17'hf06a:	data_out=16'h8522;
17'hf06b:	data_out=16'h9fd;
17'hf06c:	data_out=16'h89f0;
17'hf06d:	data_out=16'ha00;
17'hf06e:	data_out=16'h8524;
17'hf06f:	data_out=16'h8a00;
17'hf070:	data_out=16'h8527;
17'hf071:	data_out=16'h9c0;
17'hf072:	data_out=16'h89e8;
17'hf073:	data_out=16'h803a;
17'hf074:	data_out=16'h8a00;
17'hf075:	data_out=16'h84fb;
17'hf076:	data_out=16'h9fe;
17'hf077:	data_out=16'h89fe;
17'hf078:	data_out=16'h8a00;
17'hf079:	data_out=16'h8350;
17'hf07a:	data_out=16'h9fb;
17'hf07b:	data_out=16'h84f7;
17'hf07c:	data_out=16'h9ff;
17'hf07d:	data_out=16'h9ff;
17'hf07e:	data_out=16'ha2;
17'hf07f:	data_out=16'h89cd;
17'hf080:	data_out=16'h8073;
17'hf081:	data_out=16'h4d1;
17'hf082:	data_out=16'h8a00;
17'hf083:	data_out=16'h89fd;
17'hf084:	data_out=16'h9f2;
17'hf085:	data_out=16'h8a00;
17'hf086:	data_out=16'h9fe;
17'hf087:	data_out=16'h9fb;
17'hf088:	data_out=16'h9da;
17'hf089:	data_out=16'h9fe;
17'hf08a:	data_out=16'h710;
17'hf08b:	data_out=16'ha00;
17'hf08c:	data_out=16'h9d8;
17'hf08d:	data_out=16'h8a00;
17'hf08e:	data_out=16'h866a;
17'hf08f:	data_out=16'h89fa;
17'hf090:	data_out=16'h80d9;
17'hf091:	data_out=16'ha00;
17'hf092:	data_out=16'h99f;
17'hf093:	data_out=16'h557;
17'hf094:	data_out=16'h8586;
17'hf095:	data_out=16'h89ff;
17'hf096:	data_out=16'h8a00;
17'hf097:	data_out=16'h89ba;
17'hf098:	data_out=16'h21b;
17'hf099:	data_out=16'hb0;
17'hf09a:	data_out=16'h8a00;
17'hf09b:	data_out=16'h38;
17'hf09c:	data_out=16'h8a00;
17'hf09d:	data_out=16'ha00;
17'hf09e:	data_out=16'h833e;
17'hf09f:	data_out=16'h9f5;
17'hf0a0:	data_out=16'h987;
17'hf0a1:	data_out=16'h86e7;
17'hf0a2:	data_out=16'h89fc;
17'hf0a3:	data_out=16'ha00;
17'hf0a4:	data_out=16'ha00;
17'hf0a5:	data_out=16'h80d1;
17'hf0a6:	data_out=16'h8513;
17'hf0a7:	data_out=16'ha00;
17'hf0a8:	data_out=16'h8730;
17'hf0a9:	data_out=16'h8a00;
17'hf0aa:	data_out=16'h871f;
17'hf0ab:	data_out=16'ha00;
17'hf0ac:	data_out=16'h8a00;
17'hf0ad:	data_out=16'ha00;
17'hf0ae:	data_out=16'h2f;
17'hf0af:	data_out=16'h8498;
17'hf0b0:	data_out=16'h8a00;
17'hf0b1:	data_out=16'h9e8;
17'hf0b2:	data_out=16'h8a00;
17'hf0b3:	data_out=16'h9e2;
17'hf0b4:	data_out=16'h4dc;
17'hf0b5:	data_out=16'h9f1;
17'hf0b6:	data_out=16'h896;
17'hf0b7:	data_out=16'h89e7;
17'hf0b8:	data_out=16'h9ed;
17'hf0b9:	data_out=16'h9a5;
17'hf0ba:	data_out=16'h9fb;
17'hf0bb:	data_out=16'h9fd;
17'hf0bc:	data_out=16'h8a00;
17'hf0bd:	data_out=16'h81de;
17'hf0be:	data_out=16'h872f;
17'hf0bf:	data_out=16'h8a00;
17'hf0c0:	data_out=16'h849e;
17'hf0c1:	data_out=16'h89ff;
17'hf0c2:	data_out=16'h89df;
17'hf0c3:	data_out=16'h8a00;
17'hf0c4:	data_out=16'ha00;
17'hf0c5:	data_out=16'h89ff;
17'hf0c6:	data_out=16'h89fd;
17'hf0c7:	data_out=16'ha00;
17'hf0c8:	data_out=16'h9fd;
17'hf0c9:	data_out=16'h826c;
17'hf0ca:	data_out=16'h9fa;
17'hf0cb:	data_out=16'h88d8;
17'hf0cc:	data_out=16'h89fd;
17'hf0cd:	data_out=16'h89fb;
17'hf0ce:	data_out=16'h9f6;
17'hf0cf:	data_out=16'h8206;
17'hf0d0:	data_out=16'h8a00;
17'hf0d1:	data_out=16'h8a00;
17'hf0d2:	data_out=16'h9f9;
17'hf0d3:	data_out=16'h9ec;
17'hf0d4:	data_out=16'h8f9;
17'hf0d5:	data_out=16'h89d5;
17'hf0d6:	data_out=16'h9d6;
17'hf0d7:	data_out=16'h8166;
17'hf0d8:	data_out=16'h8a00;
17'hf0d9:	data_out=16'h89fa;
17'hf0da:	data_out=16'h9f1;
17'hf0db:	data_out=16'ha00;
17'hf0dc:	data_out=16'h317;
17'hf0dd:	data_out=16'h89fd;
17'hf0de:	data_out=16'h870e;
17'hf0df:	data_out=16'h676;
17'hf0e0:	data_out=16'h8941;
17'hf0e1:	data_out=16'h87ab;
17'hf0e2:	data_out=16'h862e;
17'hf0e3:	data_out=16'h9e6;
17'hf0e4:	data_out=16'ha00;
17'hf0e5:	data_out=16'h9ff;
17'hf0e6:	data_out=16'h9fe;
17'hf0e7:	data_out=16'h89f5;
17'hf0e8:	data_out=16'h86fe;
17'hf0e9:	data_out=16'h9e3;
17'hf0ea:	data_out=16'h8639;
17'hf0eb:	data_out=16'h89fe;
17'hf0ec:	data_out=16'h89f8;
17'hf0ed:	data_out=16'h9e5;
17'hf0ee:	data_out=16'h863d;
17'hf0ef:	data_out=16'h8a00;
17'hf0f0:	data_out=16'h8654;
17'hf0f1:	data_out=16'h875;
17'hf0f2:	data_out=16'h89ff;
17'hf0f3:	data_out=16'h8a00;
17'hf0f4:	data_out=16'h8a00;
17'hf0f5:	data_out=16'h8a00;
17'hf0f6:	data_out=16'h696;
17'hf0f7:	data_out=16'h89fb;
17'hf0f8:	data_out=16'h8a00;
17'hf0f9:	data_out=16'h8a00;
17'hf0fa:	data_out=16'h73e;
17'hf0fb:	data_out=16'h8734;
17'hf0fc:	data_out=16'h9f1;
17'hf0fd:	data_out=16'h905;
17'hf0fe:	data_out=16'h9fc;
17'hf0ff:	data_out=16'h8a00;
17'hf100:	data_out=16'h89f6;
17'hf101:	data_out=16'h89ff;
17'hf102:	data_out=16'h89fd;
17'hf103:	data_out=16'h89fe;
17'hf104:	data_out=16'h9f4;
17'hf105:	data_out=16'h8a00;
17'hf106:	data_out=16'h9ff;
17'hf107:	data_out=16'h9fd;
17'hf108:	data_out=16'h84d1;
17'hf109:	data_out=16'ha00;
17'hf10a:	data_out=16'h7a0;
17'hf10b:	data_out=16'ha00;
17'hf10c:	data_out=16'h9f6;
17'hf10d:	data_out=16'h8a00;
17'hf10e:	data_out=16'h81e6;
17'hf10f:	data_out=16'h89f6;
17'hf110:	data_out=16'h59;
17'hf111:	data_out=16'h9ac;
17'hf112:	data_out=16'h350;
17'hf113:	data_out=16'h9fc;
17'hf114:	data_out=16'h89fc;
17'hf115:	data_out=16'h8a00;
17'hf116:	data_out=16'h8a00;
17'hf117:	data_out=16'h8a00;
17'hf118:	data_out=16'h897e;
17'hf119:	data_out=16'h89b8;
17'hf11a:	data_out=16'h8a00;
17'hf11b:	data_out=16'h89fa;
17'hf11c:	data_out=16'h8a00;
17'hf11d:	data_out=16'h586;
17'hf11e:	data_out=16'h89f9;
17'hf11f:	data_out=16'h7f5;
17'hf120:	data_out=16'h89fa;
17'hf121:	data_out=16'h8167;
17'hf122:	data_out=16'h89fc;
17'hf123:	data_out=16'ha00;
17'hf124:	data_out=16'ha00;
17'hf125:	data_out=16'h795;
17'hf126:	data_out=16'h9f0;
17'hf127:	data_out=16'h9e7;
17'hf128:	data_out=16'h82f2;
17'hf129:	data_out=16'h8a00;
17'hf12a:	data_out=16'h89f5;
17'hf12b:	data_out=16'ha00;
17'hf12c:	data_out=16'h8a00;
17'hf12d:	data_out=16'ha00;
17'hf12e:	data_out=16'h8529;
17'hf12f:	data_out=16'h8a00;
17'hf130:	data_out=16'h8a00;
17'hf131:	data_out=16'h89f4;
17'hf132:	data_out=16'h8a00;
17'hf133:	data_out=16'h89fd;
17'hf134:	data_out=16'h89e7;
17'hf135:	data_out=16'h9bb;
17'hf136:	data_out=16'h89f7;
17'hf137:	data_out=16'h89fa;
17'hf138:	data_out=16'h827;
17'hf139:	data_out=16'h89fc;
17'hf13a:	data_out=16'h9de;
17'hf13b:	data_out=16'ha00;
17'hf13c:	data_out=16'h8a00;
17'hf13d:	data_out=16'h89f3;
17'hf13e:	data_out=16'h8304;
17'hf13f:	data_out=16'h8a00;
17'hf140:	data_out=16'h8568;
17'hf141:	data_out=16'h8a00;
17'hf142:	data_out=16'h9fe;
17'hf143:	data_out=16'h8a00;
17'hf144:	data_out=16'h9e7;
17'hf145:	data_out=16'h8a00;
17'hf146:	data_out=16'h89ff;
17'hf147:	data_out=16'ha00;
17'hf148:	data_out=16'h974;
17'hf149:	data_out=16'h76b;
17'hf14a:	data_out=16'h2bb;
17'hf14b:	data_out=16'ha00;
17'hf14c:	data_out=16'h7d5;
17'hf14d:	data_out=16'h89fc;
17'hf14e:	data_out=16'h8851;
17'hf14f:	data_out=16'h9fd;
17'hf150:	data_out=16'h8a00;
17'hf151:	data_out=16'h8a00;
17'hf152:	data_out=16'ha00;
17'hf153:	data_out=16'h89ff;
17'hf154:	data_out=16'h89f8;
17'hf155:	data_out=16'h895f;
17'hf156:	data_out=16'h9c8;
17'hf157:	data_out=16'h614;
17'hf158:	data_out=16'h8a00;
17'hf159:	data_out=16'h89e7;
17'hf15a:	data_out=16'h8449;
17'hf15b:	data_out=16'h9f7;
17'hf15c:	data_out=16'h8a00;
17'hf15d:	data_out=16'h89ff;
17'hf15e:	data_out=16'h8a00;
17'hf15f:	data_out=16'h89fd;
17'hf160:	data_out=16'h8827;
17'hf161:	data_out=16'h8a00;
17'hf162:	data_out=16'h881a;
17'hf163:	data_out=16'h89fe;
17'hf164:	data_out=16'ha00;
17'hf165:	data_out=16'h9fb;
17'hf166:	data_out=16'h89d7;
17'hf167:	data_out=16'h89dc;
17'hf168:	data_out=16'h81c6;
17'hf169:	data_out=16'h81a;
17'hf16a:	data_out=16'h81d5;
17'hf16b:	data_out=16'h8a00;
17'hf16c:	data_out=16'h89f9;
17'hf16d:	data_out=16'h89fe;
17'hf16e:	data_out=16'h81da;
17'hf16f:	data_out=16'h8a00;
17'hf170:	data_out=16'h81ec;
17'hf171:	data_out=16'h89f9;
17'hf172:	data_out=16'h8a00;
17'hf173:	data_out=16'h8a00;
17'hf174:	data_out=16'h8a00;
17'hf175:	data_out=16'h8a00;
17'hf176:	data_out=16'h8364;
17'hf177:	data_out=16'h89f8;
17'hf178:	data_out=16'h8a00;
17'hf179:	data_out=16'h89fe;
17'hf17a:	data_out=16'h89fd;
17'hf17b:	data_out=16'h830f;
17'hf17c:	data_out=16'h85c3;
17'hf17d:	data_out=16'h806a;
17'hf17e:	data_out=16'ha00;
17'hf17f:	data_out=16'h8a00;
17'hf180:	data_out=16'h8a00;
17'hf181:	data_out=16'h8a00;
17'hf182:	data_out=16'h8a00;
17'hf183:	data_out=16'h89fb;
17'hf184:	data_out=16'h89ea;
17'hf185:	data_out=16'h8a00;
17'hf186:	data_out=16'ha00;
17'hf187:	data_out=16'h9fc;
17'hf188:	data_out=16'h8a00;
17'hf189:	data_out=16'ha00;
17'hf18a:	data_out=16'h3da;
17'hf18b:	data_out=16'ha00;
17'hf18c:	data_out=16'h9ee;
17'hf18d:	data_out=16'h8a00;
17'hf18e:	data_out=16'h89ec;
17'hf18f:	data_out=16'h89f6;
17'hf190:	data_out=16'h8002;
17'hf191:	data_out=16'h6a1;
17'hf192:	data_out=16'h8a00;
17'hf193:	data_out=16'h9b9;
17'hf194:	data_out=16'h89f5;
17'hf195:	data_out=16'h8a00;
17'hf196:	data_out=16'h8a00;
17'hf197:	data_out=16'h89fa;
17'hf198:	data_out=16'h8a00;
17'hf199:	data_out=16'h9ff;
17'hf19a:	data_out=16'h8a00;
17'hf19b:	data_out=16'h89f9;
17'hf19c:	data_out=16'h8a00;
17'hf19d:	data_out=16'h8795;
17'hf19e:	data_out=16'h89fa;
17'hf19f:	data_out=16'h213;
17'hf1a0:	data_out=16'h89fd;
17'hf1a1:	data_out=16'h89ee;
17'hf1a2:	data_out=16'h958;
17'hf1a3:	data_out=16'h9fe;
17'hf1a4:	data_out=16'h9fe;
17'hf1a5:	data_out=16'h884;
17'hf1a6:	data_out=16'h9c5;
17'hf1a7:	data_out=16'h89e7;
17'hf1a8:	data_out=16'h89fa;
17'hf1a9:	data_out=16'h8a00;
17'hf1aa:	data_out=16'h89ed;
17'hf1ab:	data_out=16'ha00;
17'hf1ac:	data_out=16'h8a00;
17'hf1ad:	data_out=16'ha00;
17'hf1ae:	data_out=16'h77;
17'hf1af:	data_out=16'h8a00;
17'hf1b0:	data_out=16'h8a00;
17'hf1b1:	data_out=16'h8a00;
17'hf1b2:	data_out=16'h8a00;
17'hf1b3:	data_out=16'h89f7;
17'hf1b4:	data_out=16'h89f6;
17'hf1b5:	data_out=16'h89f9;
17'hf1b6:	data_out=16'h89fc;
17'hf1b7:	data_out=16'h89ea;
17'hf1b8:	data_out=16'h89aa;
17'hf1b9:	data_out=16'h89fc;
17'hf1ba:	data_out=16'h9fc;
17'hf1bb:	data_out=16'h9e3;
17'hf1bc:	data_out=16'h8a00;
17'hf1bd:	data_out=16'h89f9;
17'hf1be:	data_out=16'h89fa;
17'hf1bf:	data_out=16'h8a00;
17'hf1c0:	data_out=16'h89fa;
17'hf1c1:	data_out=16'h8a00;
17'hf1c2:	data_out=16'h9ef;
17'hf1c3:	data_out=16'h8a00;
17'hf1c4:	data_out=16'h89ed;
17'hf1c5:	data_out=16'h8a00;
17'hf1c6:	data_out=16'h8a00;
17'hf1c7:	data_out=16'ha00;
17'hf1c8:	data_out=16'h9e9;
17'hf1c9:	data_out=16'h7a0;
17'hf1ca:	data_out=16'h89ee;
17'hf1cb:	data_out=16'ha00;
17'hf1cc:	data_out=16'h9e6;
17'hf1cd:	data_out=16'h765;
17'hf1ce:	data_out=16'h89dd;
17'hf1cf:	data_out=16'ha00;
17'hf1d0:	data_out=16'h89fc;
17'hf1d1:	data_out=16'h8a00;
17'hf1d2:	data_out=16'ha00;
17'hf1d3:	data_out=16'h89fd;
17'hf1d4:	data_out=16'h89fb;
17'hf1d5:	data_out=16'h89e2;
17'hf1d6:	data_out=16'h664;
17'hf1d7:	data_out=16'h88ce;
17'hf1d8:	data_out=16'h8a00;
17'hf1d9:	data_out=16'h89d4;
17'hf1da:	data_out=16'h89f1;
17'hf1db:	data_out=16'h889e;
17'hf1dc:	data_out=16'h8a00;
17'hf1dd:	data_out=16'h8a00;
17'hf1de:	data_out=16'h89ff;
17'hf1df:	data_out=16'h89f7;
17'hf1e0:	data_out=16'h9b6;
17'hf1e1:	data_out=16'h8a00;
17'hf1e2:	data_out=16'h8248;
17'hf1e3:	data_out=16'h89f8;
17'hf1e4:	data_out=16'h9f9;
17'hf1e5:	data_out=16'h9f7;
17'hf1e6:	data_out=16'h9f1;
17'hf1e7:	data_out=16'h899f;
17'hf1e8:	data_out=16'h89f1;
17'hf1e9:	data_out=16'h89fe;
17'hf1ea:	data_out=16'h89f5;
17'hf1eb:	data_out=16'h8a00;
17'hf1ec:	data_out=16'h8a00;
17'hf1ed:	data_out=16'h89f8;
17'hf1ee:	data_out=16'h89f5;
17'hf1ef:	data_out=16'h8a00;
17'hf1f0:	data_out=16'h89f2;
17'hf1f1:	data_out=16'h89fa;
17'hf1f2:	data_out=16'h89ff;
17'hf1f3:	data_out=16'h89ff;
17'hf1f4:	data_out=16'h8a00;
17'hf1f5:	data_out=16'h8a00;
17'hf1f6:	data_out=16'h9ff;
17'hf1f7:	data_out=16'h89f0;
17'hf1f8:	data_out=16'h8a00;
17'hf1f9:	data_out=16'h8a00;
17'hf1fa:	data_out=16'h89fc;
17'hf1fb:	data_out=16'h89fb;
17'hf1fc:	data_out=16'h8a00;
17'hf1fd:	data_out=16'h8a00;
17'hf1fe:	data_out=16'ha00;
17'hf1ff:	data_out=16'h8a00;
17'hf200:	data_out=16'h8a00;
17'hf201:	data_out=16'h8a00;
17'hf202:	data_out=16'h8a00;
17'hf203:	data_out=16'h89b5;
17'hf204:	data_out=16'h89de;
17'hf205:	data_out=16'h8a00;
17'hf206:	data_out=16'ha00;
17'hf207:	data_out=16'h70e;
17'hf208:	data_out=16'h8a00;
17'hf209:	data_out=16'ha00;
17'hf20a:	data_out=16'h9eb;
17'hf20b:	data_out=16'ha00;
17'hf20c:	data_out=16'h51e;
17'hf20d:	data_out=16'h8a00;
17'hf20e:	data_out=16'h8979;
17'hf20f:	data_out=16'h89d9;
17'hf210:	data_out=16'h9f7;
17'hf211:	data_out=16'h829d;
17'hf212:	data_out=16'h8a00;
17'hf213:	data_out=16'h4f0;
17'hf214:	data_out=16'h89b6;
17'hf215:	data_out=16'h8a00;
17'hf216:	data_out=16'h8a00;
17'hf217:	data_out=16'h8965;
17'hf218:	data_out=16'h8a00;
17'hf219:	data_out=16'h9fb;
17'hf21a:	data_out=16'h89e6;
17'hf21b:	data_out=16'h89d9;
17'hf21c:	data_out=16'h8a00;
17'hf21d:	data_out=16'h88c2;
17'hf21e:	data_out=16'h89da;
17'hf21f:	data_out=16'h888c;
17'hf220:	data_out=16'h89f5;
17'hf221:	data_out=16'h8981;
17'hf222:	data_out=16'ha00;
17'hf223:	data_out=16'h9ec;
17'hf224:	data_out=16'h9ed;
17'hf225:	data_out=16'h9f7;
17'hf226:	data_out=16'h7f7;
17'hf227:	data_out=16'h89ea;
17'hf228:	data_out=16'h8996;
17'hf229:	data_out=16'h8757;
17'hf22a:	data_out=16'h8999;
17'hf22b:	data_out=16'h9f3;
17'hf22c:	data_out=16'h8a00;
17'hf22d:	data_out=16'ha00;
17'hf22e:	data_out=16'h81fb;
17'hf22f:	data_out=16'h89df;
17'hf230:	data_out=16'h89bd;
17'hf231:	data_out=16'h89cd;
17'hf232:	data_out=16'h8864;
17'hf233:	data_out=16'h89dc;
17'hf234:	data_out=16'h89f0;
17'hf235:	data_out=16'h89dc;
17'hf236:	data_out=16'h8a00;
17'hf237:	data_out=16'h89e3;
17'hf238:	data_out=16'h897d;
17'hf239:	data_out=16'h89e4;
17'hf23a:	data_out=16'ha00;
17'hf23b:	data_out=16'h82c1;
17'hf23c:	data_out=16'h89cf;
17'hf23d:	data_out=16'h89ea;
17'hf23e:	data_out=16'h8999;
17'hf23f:	data_out=16'h8a00;
17'hf240:	data_out=16'h89bd;
17'hf241:	data_out=16'h8a00;
17'hf242:	data_out=16'h9e2;
17'hf243:	data_out=16'h89da;
17'hf244:	data_out=16'h896a;
17'hf245:	data_out=16'h8a00;
17'hf246:	data_out=16'h8a00;
17'hf247:	data_out=16'h9e4;
17'hf248:	data_out=16'h8b3;
17'hf249:	data_out=16'h9f3;
17'hf24a:	data_out=16'h8a00;
17'hf24b:	data_out=16'ha00;
17'hf24c:	data_out=16'h9fa;
17'hf24d:	data_out=16'ha00;
17'hf24e:	data_out=16'h8a00;
17'hf24f:	data_out=16'ha00;
17'hf250:	data_out=16'h8945;
17'hf251:	data_out=16'h8a00;
17'hf252:	data_out=16'ha00;
17'hf253:	data_out=16'h89c2;
17'hf254:	data_out=16'h89d9;
17'hf255:	data_out=16'h8924;
17'hf256:	data_out=16'h89fc;
17'hf257:	data_out=16'h837b;
17'hf258:	data_out=16'h8a00;
17'hf259:	data_out=16'h898d;
17'hf25a:	data_out=16'h89f4;
17'hf25b:	data_out=16'h899b;
17'hf25c:	data_out=16'h8a00;
17'hf25d:	data_out=16'h89db;
17'hf25e:	data_out=16'h89ce;
17'hf25f:	data_out=16'h89ef;
17'hf260:	data_out=16'h99a;
17'hf261:	data_out=16'h89ce;
17'hf262:	data_out=16'h8445;
17'hf263:	data_out=16'h89dc;
17'hf264:	data_out=16'h61a;
17'hf265:	data_out=16'h9e9;
17'hf266:	data_out=16'h9e0;
17'hf267:	data_out=16'h9fe;
17'hf268:	data_out=16'h8977;
17'hf269:	data_out=16'h8a00;
17'hf26a:	data_out=16'h897f;
17'hf26b:	data_out=16'h89fd;
17'hf26c:	data_out=16'h8a00;
17'hf26d:	data_out=16'h89db;
17'hf26e:	data_out=16'h897e;
17'hf26f:	data_out=16'h8999;
17'hf270:	data_out=16'h8979;
17'hf271:	data_out=16'h89e8;
17'hf272:	data_out=16'h89af;
17'hf273:	data_out=16'h88ee;
17'hf274:	data_out=16'h89eb;
17'hf275:	data_out=16'h8a00;
17'hf276:	data_out=16'ha00;
17'hf277:	data_out=16'h8849;
17'hf278:	data_out=16'h89e6;
17'hf279:	data_out=16'h8a00;
17'hf27a:	data_out=16'h89d6;
17'hf27b:	data_out=16'h899a;
17'hf27c:	data_out=16'h8a00;
17'hf27d:	data_out=16'h89fb;
17'hf27e:	data_out=16'ha00;
17'hf27f:	data_out=16'h8a00;
17'hf280:	data_out=16'h8a00;
17'hf281:	data_out=16'h8991;
17'hf282:	data_out=16'h8a00;
17'hf283:	data_out=16'h8859;
17'hf284:	data_out=16'h89ab;
17'hf285:	data_out=16'h899a;
17'hf286:	data_out=16'ha00;
17'hf287:	data_out=16'h89ff;
17'hf288:	data_out=16'h8a00;
17'hf289:	data_out=16'ha00;
17'hf28a:	data_out=16'ha00;
17'hf28b:	data_out=16'ha00;
17'hf28c:	data_out=16'h89fc;
17'hf28d:	data_out=16'h8a00;
17'hf28e:	data_out=16'h89ee;
17'hf28f:	data_out=16'h89f2;
17'hf290:	data_out=16'ha00;
17'hf291:	data_out=16'h71e;
17'hf292:	data_out=16'h8a00;
17'hf293:	data_out=16'h8872;
17'hf294:	data_out=16'h89af;
17'hf295:	data_out=16'h89ff;
17'hf296:	data_out=16'h89e3;
17'hf297:	data_out=16'h8952;
17'hf298:	data_out=16'h8a00;
17'hf299:	data_out=16'h9fc;
17'hf29a:	data_out=16'h897f;
17'hf29b:	data_out=16'h89f3;
17'hf29c:	data_out=16'h89f6;
17'hf29d:	data_out=16'h828a;
17'hf29e:	data_out=16'h89d3;
17'hf29f:	data_out=16'h88ae;
17'hf2a0:	data_out=16'h89f5;
17'hf2a1:	data_out=16'h89eb;
17'hf2a2:	data_out=16'ha00;
17'hf2a3:	data_out=16'h9f9;
17'hf2a4:	data_out=16'h9f9;
17'hf2a5:	data_out=16'ha00;
17'hf2a6:	data_out=16'h86d2;
17'hf2a7:	data_out=16'h89f2;
17'hf2a8:	data_out=16'h89ef;
17'hf2a9:	data_out=16'h9b8;
17'hf2aa:	data_out=16'h8911;
17'hf2ab:	data_out=16'h8362;
17'hf2ac:	data_out=16'h89d2;
17'hf2ad:	data_out=16'ha00;
17'hf2ae:	data_out=16'h8241;
17'hf2af:	data_out=16'h89ce;
17'hf2b0:	data_out=16'h891f;
17'hf2b1:	data_out=16'h83a9;
17'hf2b2:	data_out=16'h81d1;
17'hf2b3:	data_out=16'h89ed;
17'hf2b4:	data_out=16'h891b;
17'hf2b5:	data_out=16'h898c;
17'hf2b6:	data_out=16'h8a00;
17'hf2b7:	data_out=16'h8a00;
17'hf2b8:	data_out=16'h8997;
17'hf2b9:	data_out=16'h89f5;
17'hf2ba:	data_out=16'ha00;
17'hf2bb:	data_out=16'h824c;
17'hf2bc:	data_out=16'h89d0;
17'hf2bd:	data_out=16'h89be;
17'hf2be:	data_out=16'h89ef;
17'hf2bf:	data_out=16'h899d;
17'hf2c0:	data_out=16'h8899;
17'hf2c1:	data_out=16'h8a00;
17'hf2c2:	data_out=16'ha00;
17'hf2c3:	data_out=16'h2f8;
17'hf2c4:	data_out=16'h86b4;
17'hf2c5:	data_out=16'h89ff;
17'hf2c6:	data_out=16'h8a00;
17'hf2c7:	data_out=16'h69a;
17'hf2c8:	data_out=16'h24;
17'hf2c9:	data_out=16'h9fe;
17'hf2ca:	data_out=16'h8a00;
17'hf2cb:	data_out=16'ha00;
17'hf2cc:	data_out=16'ha00;
17'hf2cd:	data_out=16'ha00;
17'hf2ce:	data_out=16'h8a00;
17'hf2cf:	data_out=16'ha00;
17'hf2d0:	data_out=16'h83ed;
17'hf2d1:	data_out=16'h8a00;
17'hf2d2:	data_out=16'ha00;
17'hf2d3:	data_out=16'h89f3;
17'hf2d4:	data_out=16'h89ed;
17'hf2d5:	data_out=16'h8990;
17'hf2d6:	data_out=16'h8a00;
17'hf2d7:	data_out=16'h89d8;
17'hf2d8:	data_out=16'h8a00;
17'hf2d9:	data_out=16'h1a6;
17'hf2da:	data_out=16'h8a00;
17'hf2db:	data_out=16'h8985;
17'hf2dc:	data_out=16'h8a00;
17'hf2dd:	data_out=16'h8952;
17'hf2de:	data_out=16'h8929;
17'hf2df:	data_out=16'h89f8;
17'hf2e0:	data_out=16'h9f5;
17'hf2e1:	data_out=16'h87ef;
17'hf2e2:	data_out=16'h833c;
17'hf2e3:	data_out=16'h89f3;
17'hf2e4:	data_out=16'h5c5;
17'hf2e5:	data_out=16'ha00;
17'hf2e6:	data_out=16'h603;
17'hf2e7:	data_out=16'ha00;
17'hf2e8:	data_out=16'h89e4;
17'hf2e9:	data_out=16'h8a00;
17'hf2ea:	data_out=16'h89eb;
17'hf2eb:	data_out=16'h896d;
17'hf2ec:	data_out=16'h89fe;
17'hf2ed:	data_out=16'h89f1;
17'hf2ee:	data_out=16'h89eb;
17'hf2ef:	data_out=16'h8728;
17'hf2f0:	data_out=16'h89ee;
17'hf2f1:	data_out=16'h8a00;
17'hf2f2:	data_out=16'h80c9;
17'hf2f3:	data_out=16'h8262;
17'hf2f4:	data_out=16'h89d6;
17'hf2f5:	data_out=16'h89d5;
17'hf2f6:	data_out=16'ha00;
17'hf2f7:	data_out=16'h853c;
17'hf2f8:	data_out=16'h622;
17'hf2f9:	data_out=16'h8a00;
17'hf2fa:	data_out=16'h89de;
17'hf2fb:	data_out=16'h89ef;
17'hf2fc:	data_out=16'h8a00;
17'hf2fd:	data_out=16'h89f9;
17'hf2fe:	data_out=16'ha00;
17'hf2ff:	data_out=16'h89eb;
17'hf300:	data_out=16'h8a00;
17'hf301:	data_out=16'h89f2;
17'hf302:	data_out=16'h8a00;
17'hf303:	data_out=16'h8881;
17'hf304:	data_out=16'h8811;
17'hf305:	data_out=16'h8997;
17'hf306:	data_out=16'ha00;
17'hf307:	data_out=16'h89a3;
17'hf308:	data_out=16'h8a00;
17'hf309:	data_out=16'ha00;
17'hf30a:	data_out=16'ha00;
17'hf30b:	data_out=16'h51c;
17'hf30c:	data_out=16'h830c;
17'hf30d:	data_out=16'h8a00;
17'hf30e:	data_out=16'h8a00;
17'hf30f:	data_out=16'h8a00;
17'hf310:	data_out=16'ha00;
17'hf311:	data_out=16'ha00;
17'hf312:	data_out=16'h8a00;
17'hf313:	data_out=16'h89ff;
17'hf314:	data_out=16'h8a00;
17'hf315:	data_out=16'h89ff;
17'hf316:	data_out=16'h8982;
17'hf317:	data_out=16'h8a00;
17'hf318:	data_out=16'h8a00;
17'hf319:	data_out=16'ha00;
17'hf31a:	data_out=16'h8909;
17'hf31b:	data_out=16'h8a00;
17'hf31c:	data_out=16'h8a00;
17'hf31d:	data_out=16'h314;
17'hf31e:	data_out=16'h8a00;
17'hf31f:	data_out=16'h89c3;
17'hf320:	data_out=16'h89fc;
17'hf321:	data_out=16'h8a00;
17'hf322:	data_out=16'ha00;
17'hf323:	data_out=16'ha00;
17'hf324:	data_out=16'ha00;
17'hf325:	data_out=16'ha00;
17'hf326:	data_out=16'h89f7;
17'hf327:	data_out=16'h89ff;
17'hf328:	data_out=16'h8a00;
17'hf329:	data_out=16'h7fb;
17'hf32a:	data_out=16'h89d5;
17'hf32b:	data_out=16'h87af;
17'hf32c:	data_out=16'h8940;
17'hf32d:	data_out=16'ha00;
17'hf32e:	data_out=16'h86a0;
17'hf32f:	data_out=16'h89f3;
17'hf330:	data_out=16'h889a;
17'hf331:	data_out=16'h8028;
17'hf332:	data_out=16'h9fa;
17'hf333:	data_out=16'h8a00;
17'hf334:	data_out=16'h8888;
17'hf335:	data_out=16'h898f;
17'hf336:	data_out=16'h8a00;
17'hf337:	data_out=16'h8a00;
17'hf338:	data_out=16'h89fc;
17'hf339:	data_out=16'h8a00;
17'hf33a:	data_out=16'ha00;
17'hf33b:	data_out=16'h2a;
17'hf33c:	data_out=16'h8a00;
17'hf33d:	data_out=16'h89cc;
17'hf33e:	data_out=16'h8a00;
17'hf33f:	data_out=16'h8999;
17'hf340:	data_out=16'h8034;
17'hf341:	data_out=16'h8a00;
17'hf342:	data_out=16'ha00;
17'hf343:	data_out=16'h9fc;
17'hf344:	data_out=16'h88f2;
17'hf345:	data_out=16'h89ff;
17'hf346:	data_out=16'h8a00;
17'hf347:	data_out=16'h828d;
17'hf348:	data_out=16'h8166;
17'hf349:	data_out=16'ha00;
17'hf34a:	data_out=16'h89ec;
17'hf34b:	data_out=16'ha00;
17'hf34c:	data_out=16'ha00;
17'hf34d:	data_out=16'ha00;
17'hf34e:	data_out=16'h8a00;
17'hf34f:	data_out=16'ha00;
17'hf350:	data_out=16'h8b0;
17'hf351:	data_out=16'h8a00;
17'hf352:	data_out=16'ha00;
17'hf353:	data_out=16'h8a00;
17'hf354:	data_out=16'h89fe;
17'hf355:	data_out=16'h8a00;
17'hf356:	data_out=16'h8a00;
17'hf357:	data_out=16'h89fc;
17'hf358:	data_out=16'h8a00;
17'hf359:	data_out=16'ha00;
17'hf35a:	data_out=16'h8a00;
17'hf35b:	data_out=16'h89c0;
17'hf35c:	data_out=16'h8a00;
17'hf35d:	data_out=16'h86cf;
17'hf35e:	data_out=16'h8862;
17'hf35f:	data_out=16'h89f9;
17'hf360:	data_out=16'h9f2;
17'hf361:	data_out=16'h8847;
17'hf362:	data_out=16'h86e0;
17'hf363:	data_out=16'h8a00;
17'hf364:	data_out=16'h649;
17'hf365:	data_out=16'ha00;
17'hf366:	data_out=16'h80f5;
17'hf367:	data_out=16'ha00;
17'hf368:	data_out=16'h8a00;
17'hf369:	data_out=16'h8a00;
17'hf36a:	data_out=16'h8a00;
17'hf36b:	data_out=16'h85d5;
17'hf36c:	data_out=16'h8a00;
17'hf36d:	data_out=16'h8a00;
17'hf36e:	data_out=16'h8a00;
17'hf36f:	data_out=16'h8212;
17'hf370:	data_out=16'h8a00;
17'hf371:	data_out=16'h8a00;
17'hf372:	data_out=16'ha00;
17'hf373:	data_out=16'h8319;
17'hf374:	data_out=16'h89bc;
17'hf375:	data_out=16'h8a00;
17'hf376:	data_out=16'ha00;
17'hf377:	data_out=16'hc4;
17'hf378:	data_out=16'h9fa;
17'hf379:	data_out=16'h8a00;
17'hf37a:	data_out=16'h8a00;
17'hf37b:	data_out=16'h8a00;
17'hf37c:	data_out=16'h8a00;
17'hf37d:	data_out=16'h89ed;
17'hf37e:	data_out=16'ha00;
17'hf37f:	data_out=16'h89d3;
17'hf380:	data_out=16'h8a00;
17'hf381:	data_out=16'h8a00;
17'hf382:	data_out=16'h8a00;
17'hf383:	data_out=16'h89f1;
17'hf384:	data_out=16'h8484;
17'hf385:	data_out=16'h8495;
17'hf386:	data_out=16'ha00;
17'hf387:	data_out=16'h89e5;
17'hf388:	data_out=16'h8a00;
17'hf389:	data_out=16'ha00;
17'hf38a:	data_out=16'h9ff;
17'hf38b:	data_out=16'h897c;
17'hf38c:	data_out=16'h8961;
17'hf38d:	data_out=16'h8a00;
17'hf38e:	data_out=16'h89ff;
17'hf38f:	data_out=16'h8a00;
17'hf390:	data_out=16'ha00;
17'hf391:	data_out=16'ha00;
17'hf392:	data_out=16'h8a00;
17'hf393:	data_out=16'h8a00;
17'hf394:	data_out=16'h8a00;
17'hf395:	data_out=16'h89fe;
17'hf396:	data_out=16'h89fc;
17'hf397:	data_out=16'h8a00;
17'hf398:	data_out=16'h8a00;
17'hf399:	data_out=16'h9fe;
17'hf39a:	data_out=16'h180;
17'hf39b:	data_out=16'h8a00;
17'hf39c:	data_out=16'h8a00;
17'hf39d:	data_out=16'h8157;
17'hf39e:	data_out=16'h8a00;
17'hf39f:	data_out=16'h89cf;
17'hf3a0:	data_out=16'h89f6;
17'hf3a1:	data_out=16'h89fe;
17'hf3a2:	data_out=16'ha00;
17'hf3a3:	data_out=16'h831a;
17'hf3a4:	data_out=16'h83c2;
17'hf3a5:	data_out=16'ha00;
17'hf3a6:	data_out=16'h8a00;
17'hf3a7:	data_out=16'h89ff;
17'hf3a8:	data_out=16'h8a00;
17'hf3a9:	data_out=16'h6c6;
17'hf3aa:	data_out=16'h89b9;
17'hf3ab:	data_out=16'h89fb;
17'hf3ac:	data_out=16'h89be;
17'hf3ad:	data_out=16'ha00;
17'hf3ae:	data_out=16'h8678;
17'hf3af:	data_out=16'h89ff;
17'hf3b0:	data_out=16'h89e2;
17'hf3b1:	data_out=16'h8748;
17'hf3b2:	data_out=16'h9ff;
17'hf3b3:	data_out=16'h8a00;
17'hf3b4:	data_out=16'h8a00;
17'hf3b5:	data_out=16'h89ff;
17'hf3b6:	data_out=16'h8a00;
17'hf3b7:	data_out=16'h8a00;
17'hf3b8:	data_out=16'h89fd;
17'hf3b9:	data_out=16'h8a00;
17'hf3ba:	data_out=16'ha00;
17'hf3bb:	data_out=16'h8986;
17'hf3bc:	data_out=16'h8a00;
17'hf3bd:	data_out=16'h8722;
17'hf3be:	data_out=16'h8a00;
17'hf3bf:	data_out=16'h84a6;
17'hf3c0:	data_out=16'ha00;
17'hf3c1:	data_out=16'h8a00;
17'hf3c2:	data_out=16'ha00;
17'hf3c3:	data_out=16'h9ed;
17'hf3c4:	data_out=16'h89fb;
17'hf3c5:	data_out=16'h89fe;
17'hf3c6:	data_out=16'h8a00;
17'hf3c7:	data_out=16'h8701;
17'hf3c8:	data_out=16'ha00;
17'hf3c9:	data_out=16'ha00;
17'hf3ca:	data_out=16'h89cb;
17'hf3cb:	data_out=16'ha00;
17'hf3cc:	data_out=16'ha00;
17'hf3cd:	data_out=16'ha00;
17'hf3ce:	data_out=16'h8a00;
17'hf3cf:	data_out=16'ha00;
17'hf3d0:	data_out=16'ha00;
17'hf3d1:	data_out=16'h8a00;
17'hf3d2:	data_out=16'ha00;
17'hf3d3:	data_out=16'h8a00;
17'hf3d4:	data_out=16'h89fe;
17'hf3d5:	data_out=16'h8a00;
17'hf3d6:	data_out=16'h8a00;
17'hf3d7:	data_out=16'h89f6;
17'hf3d8:	data_out=16'h8a00;
17'hf3d9:	data_out=16'ha00;
17'hf3da:	data_out=16'h8a00;
17'hf3db:	data_out=16'h89fb;
17'hf3dc:	data_out=16'h8a00;
17'hf3dd:	data_out=16'h525;
17'hf3de:	data_out=16'h8459;
17'hf3df:	data_out=16'h8923;
17'hf3e0:	data_out=16'h86ba;
17'hf3e1:	data_out=16'h80c6;
17'hf3e2:	data_out=16'h89bd;
17'hf3e3:	data_out=16'h8a00;
17'hf3e4:	data_out=16'h830f;
17'hf3e5:	data_out=16'ha00;
17'hf3e6:	data_out=16'h89e6;
17'hf3e7:	data_out=16'ha00;
17'hf3e8:	data_out=16'h89fd;
17'hf3e9:	data_out=16'h8a00;
17'hf3ea:	data_out=16'h89fe;
17'hf3eb:	data_out=16'h47c;
17'hf3ec:	data_out=16'h8a00;
17'hf3ed:	data_out=16'h8a00;
17'hf3ee:	data_out=16'h89fe;
17'hf3ef:	data_out=16'h68b;
17'hf3f0:	data_out=16'h89fe;
17'hf3f1:	data_out=16'h8a00;
17'hf3f2:	data_out=16'ha00;
17'hf3f3:	data_out=16'h9dd;
17'hf3f4:	data_out=16'h89fc;
17'hf3f5:	data_out=16'h8a00;
17'hf3f6:	data_out=16'h8709;
17'hf3f7:	data_out=16'h420;
17'hf3f8:	data_out=16'ha00;
17'hf3f9:	data_out=16'h8a00;
17'hf3fa:	data_out=16'h8a00;
17'hf3fb:	data_out=16'h8a00;
17'hf3fc:	data_out=16'h8a00;
17'hf3fd:	data_out=16'h89a1;
17'hf3fe:	data_out=16'ha00;
17'hf3ff:	data_out=16'ha00;
17'hf400:	data_out=16'h8a00;
17'hf401:	data_out=16'h8a00;
17'hf402:	data_out=16'h8a00;
17'hf403:	data_out=16'h885e;
17'hf404:	data_out=16'h89e0;
17'hf405:	data_out=16'h5a;
17'hf406:	data_out=16'ha00;
17'hf407:	data_out=16'h8a00;
17'hf408:	data_out=16'h8a00;
17'hf409:	data_out=16'h9ff;
17'hf40a:	data_out=16'h9ff;
17'hf40b:	data_out=16'h8a00;
17'hf40c:	data_out=16'h8a00;
17'hf40d:	data_out=16'h8a00;
17'hf40e:	data_out=16'h511;
17'hf40f:	data_out=16'h8a00;
17'hf410:	data_out=16'ha00;
17'hf411:	data_out=16'ha00;
17'hf412:	data_out=16'h8a00;
17'hf413:	data_out=16'h8a00;
17'hf414:	data_out=16'h8a00;
17'hf415:	data_out=16'h89fe;
17'hf416:	data_out=16'h89fc;
17'hf417:	data_out=16'h89ff;
17'hf418:	data_out=16'h8a00;
17'hf419:	data_out=16'h89b8;
17'hf41a:	data_out=16'h5f2;
17'hf41b:	data_out=16'h8a00;
17'hf41c:	data_out=16'h8a00;
17'hf41d:	data_out=16'h85af;
17'hf41e:	data_out=16'h8a00;
17'hf41f:	data_out=16'h89b1;
17'hf420:	data_out=16'h8622;
17'hf421:	data_out=16'h534;
17'hf422:	data_out=16'ha00;
17'hf423:	data_out=16'h8a00;
17'hf424:	data_out=16'h8a00;
17'hf425:	data_out=16'ha00;
17'hf426:	data_out=16'h8a00;
17'hf427:	data_out=16'h8a00;
17'hf428:	data_out=16'h3c4;
17'hf429:	data_out=16'h9c4;
17'hf42a:	data_out=16'h8a00;
17'hf42b:	data_out=16'h8a00;
17'hf42c:	data_out=16'h8776;
17'hf42d:	data_out=16'ha00;
17'hf42e:	data_out=16'h2c7;
17'hf42f:	data_out=16'h8864;
17'hf430:	data_out=16'h8a00;
17'hf431:	data_out=16'h89fe;
17'hf432:	data_out=16'h8348;
17'hf433:	data_out=16'h8a00;
17'hf434:	data_out=16'h8a00;
17'hf435:	data_out=16'h8a00;
17'hf436:	data_out=16'h8a00;
17'hf437:	data_out=16'h8a00;
17'hf438:	data_out=16'h9e0;
17'hf439:	data_out=16'h8a00;
17'hf43a:	data_out=16'h9ff;
17'hf43b:	data_out=16'h8a00;
17'hf43c:	data_out=16'h8a00;
17'hf43d:	data_out=16'h955;
17'hf43e:	data_out=16'h39b;
17'hf43f:	data_out=16'h7b;
17'hf440:	data_out=16'h82e2;
17'hf441:	data_out=16'h8a00;
17'hf442:	data_out=16'h9f9;
17'hf443:	data_out=16'h9cd;
17'hf444:	data_out=16'h8a00;
17'hf445:	data_out=16'h89fe;
17'hf446:	data_out=16'h8a00;
17'hf447:	data_out=16'h89a5;
17'hf448:	data_out=16'h9f7;
17'hf449:	data_out=16'h9fe;
17'hf44a:	data_out=16'h8a00;
17'hf44b:	data_out=16'ha00;
17'hf44c:	data_out=16'ha00;
17'hf44d:	data_out=16'ha00;
17'hf44e:	data_out=16'h8a00;
17'hf44f:	data_out=16'ha00;
17'hf450:	data_out=16'ha00;
17'hf451:	data_out=16'h8a00;
17'hf452:	data_out=16'h89d6;
17'hf453:	data_out=16'h8a00;
17'hf454:	data_out=16'h87e0;
17'hf455:	data_out=16'h8a00;
17'hf456:	data_out=16'h8a00;
17'hf457:	data_out=16'h9f;
17'hf458:	data_out=16'h8a00;
17'hf459:	data_out=16'ha00;
17'hf45a:	data_out=16'h8a00;
17'hf45b:	data_out=16'h8a00;
17'hf45c:	data_out=16'h8a00;
17'hf45d:	data_out=16'h9ff;
17'hf45e:	data_out=16'h2c4;
17'hf45f:	data_out=16'h816f;
17'hf460:	data_out=16'h8a00;
17'hf461:	data_out=16'h22;
17'hf462:	data_out=16'h88ce;
17'hf463:	data_out=16'h8a00;
17'hf464:	data_out=16'h8536;
17'hf465:	data_out=16'ha00;
17'hf466:	data_out=16'h8a00;
17'hf467:	data_out=16'ha00;
17'hf468:	data_out=16'h532;
17'hf469:	data_out=16'h8a00;
17'hf46a:	data_out=16'h513;
17'hf46b:	data_out=16'h9fb;
17'hf46c:	data_out=16'h8901;
17'hf46d:	data_out=16'h8a00;
17'hf46e:	data_out=16'h512;
17'hf46f:	data_out=16'h87cc;
17'hf470:	data_out=16'h4ea;
17'hf471:	data_out=16'h8a00;
17'hf472:	data_out=16'ha00;
17'hf473:	data_out=16'ha00;
17'hf474:	data_out=16'h8a00;
17'hf475:	data_out=16'h8a00;
17'hf476:	data_out=16'h89f6;
17'hf477:	data_out=16'h8329;
17'hf478:	data_out=16'ha00;
17'hf479:	data_out=16'h8a00;
17'hf47a:	data_out=16'h8a00;
17'hf47b:	data_out=16'h38a;
17'hf47c:	data_out=16'h8a00;
17'hf47d:	data_out=16'h899b;
17'hf47e:	data_out=16'ha00;
17'hf47f:	data_out=16'ha00;
17'hf480:	data_out=16'h8a00;
17'hf481:	data_out=16'h8a00;
17'hf482:	data_out=16'h8a00;
17'hf483:	data_out=16'h895;
17'hf484:	data_out=16'h8a00;
17'hf485:	data_out=16'h827e;
17'hf486:	data_out=16'ha00;
17'hf487:	data_out=16'h8a00;
17'hf488:	data_out=16'h8a00;
17'hf489:	data_out=16'h981;
17'hf48a:	data_out=16'h28;
17'hf48b:	data_out=16'h8a00;
17'hf48c:	data_out=16'h8a00;
17'hf48d:	data_out=16'h8a00;
17'hf48e:	data_out=16'h3e3;
17'hf48f:	data_out=16'h8a00;
17'hf490:	data_out=16'h9f4;
17'hf491:	data_out=16'ha00;
17'hf492:	data_out=16'h880b;
17'hf493:	data_out=16'h6e4;
17'hf494:	data_out=16'h21b;
17'hf495:	data_out=16'h894a;
17'hf496:	data_out=16'h57c;
17'hf497:	data_out=16'h851c;
17'hf498:	data_out=16'h8a00;
17'hf499:	data_out=16'h8a00;
17'hf49a:	data_out=16'h705;
17'hf49b:	data_out=16'h8a00;
17'hf49c:	data_out=16'h8a00;
17'hf49d:	data_out=16'h8a00;
17'hf49e:	data_out=16'h8cc;
17'hf49f:	data_out=16'h9f2;
17'hf4a0:	data_out=16'h862;
17'hf4a1:	data_out=16'h48b;
17'hf4a2:	data_out=16'ha00;
17'hf4a3:	data_out=16'h8a00;
17'hf4a4:	data_out=16'h8a00;
17'hf4a5:	data_out=16'h9c7;
17'hf4a6:	data_out=16'h8a00;
17'hf4a7:	data_out=16'h8a00;
17'hf4a8:	data_out=16'h414;
17'hf4a9:	data_out=16'h9c8;
17'hf4aa:	data_out=16'h849b;
17'hf4ab:	data_out=16'h8a00;
17'hf4ac:	data_out=16'h904;
17'hf4ad:	data_out=16'h9e6;
17'hf4ae:	data_out=16'h9e4;
17'hf4af:	data_out=16'h749;
17'hf4b0:	data_out=16'h8a00;
17'hf4b1:	data_out=16'h8a00;
17'hf4b2:	data_out=16'h89ec;
17'hf4b3:	data_out=16'h771;
17'hf4b4:	data_out=16'h8a00;
17'hf4b5:	data_out=16'h8a00;
17'hf4b6:	data_out=16'h8a00;
17'hf4b7:	data_out=16'h8a00;
17'hf4b8:	data_out=16'ha00;
17'hf4b9:	data_out=16'h822;
17'hf4ba:	data_out=16'h912;
17'hf4bb:	data_out=16'h8a00;
17'hf4bc:	data_out=16'h8a00;
17'hf4bd:	data_out=16'h9a9;
17'hf4be:	data_out=16'h3fc;
17'hf4bf:	data_out=16'h8254;
17'hf4c0:	data_out=16'h856b;
17'hf4c1:	data_out=16'h8a00;
17'hf4c2:	data_out=16'h8533;
17'hf4c3:	data_out=16'h9d6;
17'hf4c4:	data_out=16'h8a00;
17'hf4c5:	data_out=16'h88f5;
17'hf4c6:	data_out=16'h8a00;
17'hf4c7:	data_out=16'h89e9;
17'hf4c8:	data_out=16'h9e6;
17'hf4c9:	data_out=16'h742;
17'hf4ca:	data_out=16'h8a00;
17'hf4cb:	data_out=16'h9a4;
17'hf4cc:	data_out=16'ha00;
17'hf4cd:	data_out=16'ha00;
17'hf4ce:	data_out=16'h3bf;
17'hf4cf:	data_out=16'h9fd;
17'hf4d0:	data_out=16'h9f5;
17'hf4d1:	data_out=16'h8a00;
17'hf4d2:	data_out=16'h8a00;
17'hf4d3:	data_out=16'h8a00;
17'hf4d4:	data_out=16'h7e3;
17'hf4d5:	data_out=16'h8a00;
17'hf4d6:	data_out=16'h8a00;
17'hf4d7:	data_out=16'h81d1;
17'hf4d8:	data_out=16'h8a00;
17'hf4d9:	data_out=16'ha00;
17'hf4da:	data_out=16'h8a00;
17'hf4db:	data_out=16'h8a00;
17'hf4dc:	data_out=16'h8a00;
17'hf4dd:	data_out=16'h9ee;
17'hf4de:	data_out=16'h9c4;
17'hf4df:	data_out=16'h9f9;
17'hf4e0:	data_out=16'h8a00;
17'hf4e1:	data_out=16'h857b;
17'hf4e2:	data_out=16'h81ac;
17'hf4e3:	data_out=16'h517;
17'hf4e4:	data_out=16'h8a00;
17'hf4e5:	data_out=16'h83de;
17'hf4e6:	data_out=16'h8a00;
17'hf4e7:	data_out=16'ha00;
17'hf4e8:	data_out=16'h4db;
17'hf4e9:	data_out=16'h8a00;
17'hf4ea:	data_out=16'h3a8;
17'hf4eb:	data_out=16'h9c8;
17'hf4ec:	data_out=16'h8325;
17'hf4ed:	data_out=16'h5ff;
17'hf4ee:	data_out=16'h3a7;
17'hf4ef:	data_out=16'h8953;
17'hf4f0:	data_out=16'h39c;
17'hf4f1:	data_out=16'h8a00;
17'hf4f2:	data_out=16'ha00;
17'hf4f3:	data_out=16'ha00;
17'hf4f4:	data_out=16'h8a00;
17'hf4f5:	data_out=16'h8a00;
17'hf4f6:	data_out=16'h8a00;
17'hf4f7:	data_out=16'h8d3;
17'hf4f8:	data_out=16'h9f6;
17'hf4f9:	data_out=16'h1b3;
17'hf4fa:	data_out=16'h821c;
17'hf4fb:	data_out=16'h3f1;
17'hf4fc:	data_out=16'h8a00;
17'hf4fd:	data_out=16'h9fe;
17'hf4fe:	data_out=16'ha00;
17'hf4ff:	data_out=16'ha00;
17'hf500:	data_out=16'h89e9;
17'hf501:	data_out=16'h8a00;
17'hf502:	data_out=16'h8a00;
17'hf503:	data_out=16'h961;
17'hf504:	data_out=16'h8a00;
17'hf505:	data_out=16'h8a00;
17'hf506:	data_out=16'ha00;
17'hf507:	data_out=16'h8a00;
17'hf508:	data_out=16'h8a00;
17'hf509:	data_out=16'h9bd;
17'hf50a:	data_out=16'h8a00;
17'hf50b:	data_out=16'h8a00;
17'hf50c:	data_out=16'h8a00;
17'hf50d:	data_out=16'h91f;
17'hf50e:	data_out=16'h27a;
17'hf50f:	data_out=16'h894c;
17'hf510:	data_out=16'h9d5;
17'hf511:	data_out=16'h86e0;
17'hf512:	data_out=16'h958;
17'hf513:	data_out=16'h9ea;
17'hf514:	data_out=16'h954;
17'hf515:	data_out=16'h9a0;
17'hf516:	data_out=16'h97d;
17'hf517:	data_out=16'h891;
17'hf518:	data_out=16'h8a00;
17'hf519:	data_out=16'h8a00;
17'hf51a:	data_out=16'h84b3;
17'hf51b:	data_out=16'h8a00;
17'hf51c:	data_out=16'h8a00;
17'hf51d:	data_out=16'h8a00;
17'hf51e:	data_out=16'h9bc;
17'hf51f:	data_out=16'h9ed;
17'hf520:	data_out=16'h8b5;
17'hf521:	data_out=16'h376;
17'hf522:	data_out=16'ha00;
17'hf523:	data_out=16'h8a00;
17'hf524:	data_out=16'h8a00;
17'hf525:	data_out=16'h981;
17'hf526:	data_out=16'h8a00;
17'hf527:	data_out=16'h8a00;
17'hf528:	data_out=16'h32e;
17'hf529:	data_out=16'h89cf;
17'hf52a:	data_out=16'h51a;
17'hf52b:	data_out=16'h8a00;
17'hf52c:	data_out=16'h9be;
17'hf52d:	data_out=16'h89fe;
17'hf52e:	data_out=16'h9b8;
17'hf52f:	data_out=16'h802;
17'hf530:	data_out=16'h8a00;
17'hf531:	data_out=16'h8a00;
17'hf532:	data_out=16'h8a00;
17'hf533:	data_out=16'h9bb;
17'hf534:	data_out=16'h8a00;
17'hf535:	data_out=16'h8a00;
17'hf536:	data_out=16'h8a00;
17'hf537:	data_out=16'h8a00;
17'hf538:	data_out=16'ha00;
17'hf539:	data_out=16'h9ca;
17'hf53a:	data_out=16'h983;
17'hf53b:	data_out=16'h8a00;
17'hf53c:	data_out=16'h8a00;
17'hf53d:	data_out=16'h9a7;
17'hf53e:	data_out=16'h31b;
17'hf53f:	data_out=16'h8a00;
17'hf540:	data_out=16'h8783;
17'hf541:	data_out=16'h8a00;
17'hf542:	data_out=16'h8a00;
17'hf543:	data_out=16'h788;
17'hf544:	data_out=16'h8a00;
17'hf545:	data_out=16'h9a7;
17'hf546:	data_out=16'h8a00;
17'hf547:	data_out=16'h9e5;
17'hf548:	data_out=16'h9ee;
17'hf549:	data_out=16'h84cb;
17'hf54a:	data_out=16'h8a00;
17'hf54b:	data_out=16'h82a7;
17'hf54c:	data_out=16'ha00;
17'hf54d:	data_out=16'ha00;
17'hf54e:	data_out=16'h757;
17'hf54f:	data_out=16'h38b;
17'hf550:	data_out=16'ha00;
17'hf551:	data_out=16'h898f;
17'hf552:	data_out=16'h8a00;
17'hf553:	data_out=16'h8a00;
17'hf554:	data_out=16'h804;
17'hf555:	data_out=16'h89f5;
17'hf556:	data_out=16'h8a00;
17'hf557:	data_out=16'h89a6;
17'hf558:	data_out=16'h8a00;
17'hf559:	data_out=16'h9f7;
17'hf55a:	data_out=16'h8a00;
17'hf55b:	data_out=16'h8a00;
17'hf55c:	data_out=16'h8a00;
17'hf55d:	data_out=16'h9d7;
17'hf55e:	data_out=16'h9ee;
17'hf55f:	data_out=16'h9f9;
17'hf560:	data_out=16'h8a00;
17'hf561:	data_out=16'h8a00;
17'hf562:	data_out=16'h56b;
17'hf563:	data_out=16'h98e;
17'hf564:	data_out=16'h8a00;
17'hf565:	data_out=16'h8a00;
17'hf566:	data_out=16'h8a00;
17'hf567:	data_out=16'h9d2;
17'hf568:	data_out=16'h3e1;
17'hf569:	data_out=16'h8a00;
17'hf56a:	data_out=16'h1f8;
17'hf56b:	data_out=16'h9b4;
17'hf56c:	data_out=16'h345;
17'hf56d:	data_out=16'h997;
17'hf56e:	data_out=16'h1f8;
17'hf56f:	data_out=16'h83b3;
17'hf570:	data_out=16'h21b;
17'hf571:	data_out=16'h672;
17'hf572:	data_out=16'h9fd;
17'hf573:	data_out=16'h9bb;
17'hf574:	data_out=16'h8a00;
17'hf575:	data_out=16'h8a00;
17'hf576:	data_out=16'h8a00;
17'hf577:	data_out=16'h957;
17'hf578:	data_out=16'h2c9;
17'hf579:	data_out=16'h9dd;
17'hf57a:	data_out=16'h90e;
17'hf57b:	data_out=16'h313;
17'hf57c:	data_out=16'h8a00;
17'hf57d:	data_out=16'h9ff;
17'hf57e:	data_out=16'ha00;
17'hf57f:	data_out=16'ha00;
17'hf580:	data_out=16'h8a00;
17'hf581:	data_out=16'h8a00;
17'hf582:	data_out=16'h8a00;
17'hf583:	data_out=16'h80f;
17'hf584:	data_out=16'h8a00;
17'hf585:	data_out=16'h8a00;
17'hf586:	data_out=16'h9f7;
17'hf587:	data_out=16'h8a00;
17'hf588:	data_out=16'h8a00;
17'hf589:	data_out=16'h99e;
17'hf58a:	data_out=16'h8a00;
17'hf58b:	data_out=16'h89f8;
17'hf58c:	data_out=16'h8a00;
17'hf58d:	data_out=16'h940;
17'hf58e:	data_out=16'h808;
17'hf58f:	data_out=16'h7dc;
17'hf590:	data_out=16'h9b0;
17'hf591:	data_out=16'h8a00;
17'hf592:	data_out=16'h9d6;
17'hf593:	data_out=16'h9fa;
17'hf594:	data_out=16'h968;
17'hf595:	data_out=16'h8980;
17'hf596:	data_out=16'h8a00;
17'hf597:	data_out=16'h613;
17'hf598:	data_out=16'h9f6;
17'hf599:	data_out=16'h8a00;
17'hf59a:	data_out=16'h8a00;
17'hf59b:	data_out=16'h8a00;
17'hf59c:	data_out=16'h82bb;
17'hf59d:	data_out=16'h8a00;
17'hf59e:	data_out=16'h9cd;
17'hf59f:	data_out=16'h9d9;
17'hf5a0:	data_out=16'h92f;
17'hf5a1:	data_out=16'h8bb;
17'hf5a2:	data_out=16'h9ba;
17'hf5a3:	data_out=16'h8a00;
17'hf5a4:	data_out=16'h8a00;
17'hf5a5:	data_out=16'h58f;
17'hf5a6:	data_out=16'h8a00;
17'hf5a7:	data_out=16'h8a00;
17'hf5a8:	data_out=16'h8e5;
17'hf5a9:	data_out=16'h8a00;
17'hf5aa:	data_out=16'h842c;
17'hf5ab:	data_out=16'h8a00;
17'hf5ac:	data_out=16'h87cf;
17'hf5ad:	data_out=16'h89fd;
17'hf5ae:	data_out=16'h636;
17'hf5af:	data_out=16'h8cd;
17'hf5b0:	data_out=16'h89f6;
17'hf5b1:	data_out=16'h8a00;
17'hf5b2:	data_out=16'h8a00;
17'hf5b3:	data_out=16'h9fe;
17'hf5b4:	data_out=16'h8a00;
17'hf5b5:	data_out=16'h8a00;
17'hf5b6:	data_out=16'h8a00;
17'hf5b7:	data_out=16'h8a00;
17'hf5b8:	data_out=16'ha00;
17'hf5b9:	data_out=16'ha00;
17'hf5ba:	data_out=16'h9c8;
17'hf5bb:	data_out=16'h8a00;
17'hf5bc:	data_out=16'h8a00;
17'hf5bd:	data_out=16'h988;
17'hf5be:	data_out=16'h8dc;
17'hf5bf:	data_out=16'h8a00;
17'hf5c0:	data_out=16'h8a00;
17'hf5c1:	data_out=16'h8a00;
17'hf5c2:	data_out=16'h8a00;
17'hf5c3:	data_out=16'h87ad;
17'hf5c4:	data_out=16'h8a00;
17'hf5c5:	data_out=16'h897c;
17'hf5c6:	data_out=16'h8a00;
17'hf5c7:	data_out=16'h9f7;
17'hf5c8:	data_out=16'h9eb;
17'hf5c9:	data_out=16'h849e;
17'hf5ca:	data_out=16'h8a00;
17'hf5cb:	data_out=16'h8a00;
17'hf5cc:	data_out=16'h86e;
17'hf5cd:	data_out=16'h9c8;
17'hf5ce:	data_out=16'h6b6;
17'hf5cf:	data_out=16'h1a5;
17'hf5d0:	data_out=16'h9b9;
17'hf5d1:	data_out=16'h89a2;
17'hf5d2:	data_out=16'h8a00;
17'hf5d3:	data_out=16'h8a00;
17'hf5d4:	data_out=16'h886;
17'hf5d5:	data_out=16'h89f2;
17'hf5d6:	data_out=16'h8a00;
17'hf5d7:	data_out=16'h242;
17'hf5d8:	data_out=16'h8a00;
17'hf5d9:	data_out=16'h86ef;
17'hf5da:	data_out=16'h89fe;
17'hf5db:	data_out=16'h8a00;
17'hf5dc:	data_out=16'h8a00;
17'hf5dd:	data_out=16'h9db;
17'hf5de:	data_out=16'ha00;
17'hf5df:	data_out=16'h9f4;
17'hf5e0:	data_out=16'h8a00;
17'hf5e1:	data_out=16'h8a00;
17'hf5e2:	data_out=16'h8a00;
17'hf5e3:	data_out=16'h9dd;
17'hf5e4:	data_out=16'h8a00;
17'hf5e5:	data_out=16'h8a00;
17'hf5e6:	data_out=16'h86c3;
17'hf5e7:	data_out=16'h8a00;
17'hf5e8:	data_out=16'h918;
17'hf5e9:	data_out=16'h89f5;
17'hf5ea:	data_out=16'h79a;
17'hf5eb:	data_out=16'h954;
17'hf5ec:	data_out=16'h8a00;
17'hf5ed:	data_out=16'h9e3;
17'hf5ee:	data_out=16'h79a;
17'hf5ef:	data_out=16'h8a00;
17'hf5f0:	data_out=16'h7cc;
17'hf5f1:	data_out=16'h760;
17'hf5f2:	data_out=16'h99f;
17'hf5f3:	data_out=16'h8a00;
17'hf5f4:	data_out=16'h8a00;
17'hf5f5:	data_out=16'h8a00;
17'hf5f6:	data_out=16'h8a00;
17'hf5f7:	data_out=16'h94e;
17'hf5f8:	data_out=16'h89ff;
17'hf5f9:	data_out=16'h15f;
17'hf5fa:	data_out=16'h97c;
17'hf5fb:	data_out=16'h8d6;
17'hf5fc:	data_out=16'h9f3;
17'hf5fd:	data_out=16'h9f4;
17'hf5fe:	data_out=16'h9ff;
17'hf5ff:	data_out=16'h9ee;
17'hf600:	data_out=16'h89cc;
17'hf601:	data_out=16'h8a00;
17'hf602:	data_out=16'h89db;
17'hf603:	data_out=16'h8980;
17'hf604:	data_out=16'h89c3;
17'hf605:	data_out=16'h8a00;
17'hf606:	data_out=16'h9c4;
17'hf607:	data_out=16'h89d4;
17'hf608:	data_out=16'h4de;
17'hf609:	data_out=16'h9a9;
17'hf60a:	data_out=16'h89fe;
17'hf60b:	data_out=16'h5c9;
17'hf60c:	data_out=16'h89ee;
17'hf60d:	data_out=16'h89ad;
17'hf60e:	data_out=16'h9fb;
17'hf60f:	data_out=16'h7e5;
17'hf610:	data_out=16'h996;
17'hf611:	data_out=16'h8966;
17'hf612:	data_out=16'h9e0;
17'hf613:	data_out=16'ha00;
17'hf614:	data_out=16'h928;
17'hf615:	data_out=16'h89dc;
17'hf616:	data_out=16'h89d6;
17'hf617:	data_out=16'h88d2;
17'hf618:	data_out=16'h9f9;
17'hf619:	data_out=16'h9d6;
17'hf61a:	data_out=16'h8a00;
17'hf61b:	data_out=16'h89fc;
17'hf61c:	data_out=16'h8472;
17'hf61d:	data_out=16'h89fe;
17'hf61e:	data_out=16'h9d6;
17'hf61f:	data_out=16'h687;
17'hf620:	data_out=16'h9c1;
17'hf621:	data_out=16'h9fc;
17'hf622:	data_out=16'h613;
17'hf623:	data_out=16'h89fc;
17'hf624:	data_out=16'h89fc;
17'hf625:	data_out=16'h801;
17'hf626:	data_out=16'h89f1;
17'hf627:	data_out=16'h89f8;
17'hf628:	data_out=16'h9fa;
17'hf629:	data_out=16'h8a00;
17'hf62a:	data_out=16'h86c8;
17'hf62b:	data_out=16'h89df;
17'hf62c:	data_out=16'h89bb;
17'hf62d:	data_out=16'h736;
17'hf62e:	data_out=16'h816c;
17'hf62f:	data_out=16'h46e;
17'hf630:	data_out=16'h946;
17'hf631:	data_out=16'h8a00;
17'hf632:	data_out=16'h8a00;
17'hf633:	data_out=16'h9f6;
17'hf634:	data_out=16'h8a00;
17'hf635:	data_out=16'h89fd;
17'hf636:	data_out=16'h5c3;
17'hf637:	data_out=16'h89f8;
17'hf638:	data_out=16'ha00;
17'hf639:	data_out=16'ha00;
17'hf63a:	data_out=16'h9d0;
17'hf63b:	data_out=16'h8a00;
17'hf63c:	data_out=16'h8a00;
17'hf63d:	data_out=16'h9cf;
17'hf63e:	data_out=16'h9fa;
17'hf63f:	data_out=16'h8a00;
17'hf640:	data_out=16'h825b;
17'hf641:	data_out=16'h89a8;
17'hf642:	data_out=16'h89e7;
17'hf643:	data_out=16'h89ca;
17'hf644:	data_out=16'h8a00;
17'hf645:	data_out=16'h89dc;
17'hf646:	data_out=16'h89f1;
17'hf647:	data_out=16'h9fb;
17'hf648:	data_out=16'h9d4;
17'hf649:	data_out=16'h778;
17'hf64a:	data_out=16'ha7;
17'hf64b:	data_out=16'h89db;
17'hf64c:	data_out=16'h6f0;
17'hf64d:	data_out=16'h7c4;
17'hf64e:	data_out=16'h859;
17'hf64f:	data_out=16'h7b8;
17'hf650:	data_out=16'h88a4;
17'hf651:	data_out=16'h89b9;
17'hf652:	data_out=16'h8a00;
17'hf653:	data_out=16'h89fc;
17'hf654:	data_out=16'h93d;
17'hf655:	data_out=16'h89d3;
17'hf656:	data_out=16'h8111;
17'hf657:	data_out=16'h9a1;
17'hf658:	data_out=16'h89ed;
17'hf659:	data_out=16'h8248;
17'hf65a:	data_out=16'h89bd;
17'hf65b:	data_out=16'h8a00;
17'hf65c:	data_out=16'h8a00;
17'hf65d:	data_out=16'h88e2;
17'hf65e:	data_out=16'ha00;
17'hf65f:	data_out=16'h9f7;
17'hf660:	data_out=16'h8a00;
17'hf661:	data_out=16'h8a00;
17'hf662:	data_out=16'h89ff;
17'hf663:	data_out=16'h9e1;
17'hf664:	data_out=16'h806f;
17'hf665:	data_out=16'h8a00;
17'hf666:	data_out=16'ha00;
17'hf667:	data_out=16'h8a00;
17'hf668:	data_out=16'h9fc;
17'hf669:	data_out=16'h93d;
17'hf66a:	data_out=16'h9fb;
17'hf66b:	data_out=16'h85b0;
17'hf66c:	data_out=16'h89da;
17'hf66d:	data_out=16'h9e5;
17'hf66e:	data_out=16'h9fb;
17'hf66f:	data_out=16'h8a00;
17'hf670:	data_out=16'h9fb;
17'hf671:	data_out=16'h3e6;
17'hf672:	data_out=16'h8b6;
17'hf673:	data_out=16'h89f0;
17'hf674:	data_out=16'h724;
17'hf675:	data_out=16'h8a00;
17'hf676:	data_out=16'h8a00;
17'hf677:	data_out=16'h7fa;
17'hf678:	data_out=16'h8a00;
17'hf679:	data_out=16'h5ff;
17'hf67a:	data_out=16'h981;
17'hf67b:	data_out=16'h9fa;
17'hf67c:	data_out=16'h9f7;
17'hf67d:	data_out=16'h9d4;
17'hf67e:	data_out=16'h9f5;
17'hf67f:	data_out=16'h62b;
17'hf680:	data_out=16'h899a;
17'hf681:	data_out=16'h89f8;
17'hf682:	data_out=16'h9b8;
17'hf683:	data_out=16'h8977;
17'hf684:	data_out=16'h8980;
17'hf685:	data_out=16'h8a00;
17'hf686:	data_out=16'h8ee;
17'hf687:	data_out=16'ha00;
17'hf688:	data_out=16'ha00;
17'hf689:	data_out=16'h9e1;
17'hf68a:	data_out=16'h89f6;
17'hf68b:	data_out=16'ha00;
17'hf68c:	data_out=16'h9e2;
17'hf68d:	data_out=16'h89d0;
17'hf68e:	data_out=16'h9f9;
17'hf68f:	data_out=16'h9ea;
17'hf690:	data_out=16'h84d;
17'hf691:	data_out=16'h8897;
17'hf692:	data_out=16'h9eb;
17'hf693:	data_out=16'h9fc;
17'hf694:	data_out=16'h951;
17'hf695:	data_out=16'h89e4;
17'hf696:	data_out=16'h89d4;
17'hf697:	data_out=16'h8930;
17'hf698:	data_out=16'h9fb;
17'hf699:	data_out=16'ha00;
17'hf69a:	data_out=16'h8a00;
17'hf69b:	data_out=16'h9fd;
17'hf69c:	data_out=16'h89dc;
17'hf69d:	data_out=16'h89ad;
17'hf69e:	data_out=16'h9c8;
17'hf69f:	data_out=16'h1d;
17'hf6a0:	data_out=16'h8871;
17'hf6a1:	data_out=16'h9f9;
17'hf6a2:	data_out=16'h89ee;
17'hf6a3:	data_out=16'h9dd;
17'hf6a4:	data_out=16'h9dd;
17'hf6a5:	data_out=16'h5f1;
17'hf6a6:	data_out=16'h533;
17'hf6a7:	data_out=16'ha00;
17'hf6a8:	data_out=16'h9f9;
17'hf6a9:	data_out=16'h8a00;
17'hf6aa:	data_out=16'h24e;
17'hf6ab:	data_out=16'ha00;
17'hf6ac:	data_out=16'h89dc;
17'hf6ad:	data_out=16'h9eb;
17'hf6ae:	data_out=16'h43d;
17'hf6af:	data_out=16'h8943;
17'hf6b0:	data_out=16'ha00;
17'hf6b1:	data_out=16'h89c7;
17'hf6b2:	data_out=16'h89fc;
17'hf6b3:	data_out=16'h9fb;
17'hf6b4:	data_out=16'h89d5;
17'hf6b5:	data_out=16'he8;
17'hf6b6:	data_out=16'h9ff;
17'hf6b7:	data_out=16'h3eb;
17'hf6b8:	data_out=16'h85fe;
17'hf6b9:	data_out=16'h9fb;
17'hf6ba:	data_out=16'h9ea;
17'hf6bb:	data_out=16'h835b;
17'hf6bc:	data_out=16'h8a00;
17'hf6bd:	data_out=16'h88af;
17'hf6be:	data_out=16'h9f9;
17'hf6bf:	data_out=16'h8a00;
17'hf6c0:	data_out=16'h89cb;
17'hf6c1:	data_out=16'h5f3;
17'hf6c2:	data_out=16'h89a8;
17'hf6c3:	data_out=16'h89c2;
17'hf6c4:	data_out=16'h890e;
17'hf6c5:	data_out=16'h89e5;
17'hf6c6:	data_out=16'h83a2;
17'hf6c7:	data_out=16'h9f7;
17'hf6c8:	data_out=16'h52b;
17'hf6c9:	data_out=16'h740;
17'hf6ca:	data_out=16'ha00;
17'hf6cb:	data_out=16'h89ae;
17'hf6cc:	data_out=16'h6da;
17'hf6cd:	data_out=16'h89b4;
17'hf6ce:	data_out=16'h9ff;
17'hf6cf:	data_out=16'h931;
17'hf6d0:	data_out=16'h89bc;
17'hf6d1:	data_out=16'h89e6;
17'hf6d2:	data_out=16'h83e;
17'hf6d3:	data_out=16'h3b;
17'hf6d4:	data_out=16'h8534;
17'hf6d5:	data_out=16'h8945;
17'hf6d6:	data_out=16'h9e2;
17'hf6d7:	data_out=16'h970;
17'hf6d8:	data_out=16'h82af;
17'hf6d9:	data_out=16'h89ba;
17'hf6da:	data_out=16'h697;
17'hf6db:	data_out=16'h8977;
17'hf6dc:	data_out=16'h8a00;
17'hf6dd:	data_out=16'h8965;
17'hf6de:	data_out=16'h8814;
17'hf6df:	data_out=16'h9f9;
17'hf6e0:	data_out=16'h89aa;
17'hf6e1:	data_out=16'h8a00;
17'hf6e2:	data_out=16'h8828;
17'hf6e3:	data_out=16'h9f9;
17'hf6e4:	data_out=16'h89ab;
17'hf6e5:	data_out=16'h894e;
17'hf6e6:	data_out=16'ha00;
17'hf6e7:	data_out=16'h8a00;
17'hf6e8:	data_out=16'h9f9;
17'hf6e9:	data_out=16'h9fc;
17'hf6ea:	data_out=16'h9f9;
17'hf6eb:	data_out=16'h895d;
17'hf6ec:	data_out=16'h89b8;
17'hf6ed:	data_out=16'h9fa;
17'hf6ee:	data_out=16'h9f9;
17'hf6ef:	data_out=16'h89ff;
17'hf6f0:	data_out=16'h9f9;
17'hf6f1:	data_out=16'h699;
17'hf6f2:	data_out=16'h89b9;
17'hf6f3:	data_out=16'h8a00;
17'hf6f4:	data_out=16'ha00;
17'hf6f5:	data_out=16'h8a00;
17'hf6f6:	data_out=16'h958;
17'hf6f7:	data_out=16'h913;
17'hf6f8:	data_out=16'h8a00;
17'hf6f9:	data_out=16'h9fb;
17'hf6fa:	data_out=16'h9f6;
17'hf6fb:	data_out=16'h9f9;
17'hf6fc:	data_out=16'h9f9;
17'hf6fd:	data_out=16'h862e;
17'hf6fe:	data_out=16'ha00;
17'hf6ff:	data_out=16'h8a00;
17'hf700:	data_out=16'h89ee;
17'hf701:	data_out=16'h8a00;
17'hf702:	data_out=16'h979;
17'hf703:	data_out=16'h8987;
17'hf704:	data_out=16'h88e7;
17'hf705:	data_out=16'h8a00;
17'hf706:	data_out=16'h89d9;
17'hf707:	data_out=16'ha00;
17'hf708:	data_out=16'h9ff;
17'hf709:	data_out=16'ha00;
17'hf70a:	data_out=16'h89fe;
17'hf70b:	data_out=16'ha00;
17'hf70c:	data_out=16'ha00;
17'hf70d:	data_out=16'h89d4;
17'hf70e:	data_out=16'h9f9;
17'hf70f:	data_out=16'h9f8;
17'hf710:	data_out=16'h988;
17'hf711:	data_out=16'h89f9;
17'hf712:	data_out=16'h9ed;
17'hf713:	data_out=16'h256;
17'hf714:	data_out=16'h85a9;
17'hf715:	data_out=16'h89f9;
17'hf716:	data_out=16'h89dc;
17'hf717:	data_out=16'h8921;
17'hf718:	data_out=16'h9f9;
17'hf719:	data_out=16'ha00;
17'hf71a:	data_out=16'h8a00;
17'hf71b:	data_out=16'h9fe;
17'hf71c:	data_out=16'h89e9;
17'hf71d:	data_out=16'h89f9;
17'hf71e:	data_out=16'h8563;
17'hf71f:	data_out=16'h6bd;
17'hf720:	data_out=16'h89c6;
17'hf721:	data_out=16'h9fa;
17'hf722:	data_out=16'h8760;
17'hf723:	data_out=16'ha00;
17'hf724:	data_out=16'ha00;
17'hf725:	data_out=16'h9c8;
17'hf726:	data_out=16'h8419;
17'hf727:	data_out=16'h9c6;
17'hf728:	data_out=16'h9fb;
17'hf729:	data_out=16'h89f1;
17'hf72a:	data_out=16'h9fd;
17'hf72b:	data_out=16'ha00;
17'hf72c:	data_out=16'h89e6;
17'hf72d:	data_out=16'h9c5;
17'hf72e:	data_out=16'h9da;
17'hf72f:	data_out=16'h8852;
17'hf730:	data_out=16'h794;
17'hf731:	data_out=16'h89fd;
17'hf732:	data_out=16'h89e8;
17'hf733:	data_out=16'h783;
17'hf734:	data_out=16'h89ff;
17'hf735:	data_out=16'h8447;
17'hf736:	data_out=16'ha00;
17'hf737:	data_out=16'h9b0;
17'hf738:	data_out=16'h8a00;
17'hf739:	data_out=16'h35c;
17'hf73a:	data_out=16'ha00;
17'hf73b:	data_out=16'ha00;
17'hf73c:	data_out=16'h89fd;
17'hf73d:	data_out=16'h899c;
17'hf73e:	data_out=16'h9fb;
17'hf73f:	data_out=16'h8a00;
17'hf740:	data_out=16'h87c2;
17'hf741:	data_out=16'h735;
17'hf742:	data_out=16'h89b9;
17'hf743:	data_out=16'h990;
17'hf744:	data_out=16'h89dc;
17'hf745:	data_out=16'h89f9;
17'hf746:	data_out=16'h89bc;
17'hf747:	data_out=16'ha00;
17'hf748:	data_out=16'h71a;
17'hf749:	data_out=16'h9f5;
17'hf74a:	data_out=16'ha00;
17'hf74b:	data_out=16'h89d0;
17'hf74c:	data_out=16'h82b;
17'hf74d:	data_out=16'h85d4;
17'hf74e:	data_out=16'h9ff;
17'hf74f:	data_out=16'h9f3;
17'hf750:	data_out=16'h89ab;
17'hf751:	data_out=16'h89cd;
17'hf752:	data_out=16'ha00;
17'hf753:	data_out=16'h949;
17'hf754:	data_out=16'h819c;
17'hf755:	data_out=16'h54f;
17'hf756:	data_out=16'h8647;
17'hf757:	data_out=16'h872f;
17'hf758:	data_out=16'h8984;
17'hf759:	data_out=16'h89c5;
17'hf75a:	data_out=16'h809c;
17'hf75b:	data_out=16'h89ec;
17'hf75c:	data_out=16'h8a00;
17'hf75d:	data_out=16'h89b1;
17'hf75e:	data_out=16'h87a1;
17'hf75f:	data_out=16'h9f9;
17'hf760:	data_out=16'h880c;
17'hf761:	data_out=16'h8a00;
17'hf762:	data_out=16'h806c;
17'hf763:	data_out=16'h88e;
17'hf764:	data_out=16'h89e0;
17'hf765:	data_out=16'h886a;
17'hf766:	data_out=16'ha00;
17'hf767:	data_out=16'h9b1;
17'hf768:	data_out=16'h9fb;
17'hf769:	data_out=16'h9fc;
17'hf76a:	data_out=16'h9f8;
17'hf76b:	data_out=16'h89ce;
17'hf76c:	data_out=16'h89f8;
17'hf76d:	data_out=16'h85a;
17'hf76e:	data_out=16'h9f8;
17'hf76f:	data_out=16'h89ff;
17'hf770:	data_out=16'h9f9;
17'hf771:	data_out=16'h9f2;
17'hf772:	data_out=16'h8a00;
17'hf773:	data_out=16'h8a00;
17'hf774:	data_out=16'h774;
17'hf775:	data_out=16'h8a00;
17'hf776:	data_out=16'ha00;
17'hf777:	data_out=16'ha00;
17'hf778:	data_out=16'h8a00;
17'hf779:	data_out=16'h9f6;
17'hf77a:	data_out=16'h695;
17'hf77b:	data_out=16'h9fb;
17'hf77c:	data_out=16'h9f7;
17'hf77d:	data_out=16'h6ac;
17'hf77e:	data_out=16'h840;
17'hf77f:	data_out=16'h8a00;
17'hf780:	data_out=16'h8a00;
17'hf781:	data_out=16'h8a00;
17'hf782:	data_out=16'h8403;
17'hf783:	data_out=16'h8988;
17'hf784:	data_out=16'h9f2;
17'hf785:	data_out=16'h8a00;
17'hf786:	data_out=16'h8995;
17'hf787:	data_out=16'ha00;
17'hf788:	data_out=16'h9b4;
17'hf789:	data_out=16'ha00;
17'hf78a:	data_out=16'h8a00;
17'hf78b:	data_out=16'ha00;
17'hf78c:	data_out=16'ha00;
17'hf78d:	data_out=16'h89d0;
17'hf78e:	data_out=16'h701;
17'hf78f:	data_out=16'h9ee;
17'hf790:	data_out=16'h99e;
17'hf791:	data_out=16'h89fe;
17'hf792:	data_out=16'h89ee;
17'hf793:	data_out=16'h88bb;
17'hf794:	data_out=16'h8940;
17'hf795:	data_out=16'h89f9;
17'hf796:	data_out=16'h89cb;
17'hf797:	data_out=16'h89a0;
17'hf798:	data_out=16'h841;
17'hf799:	data_out=16'ha00;
17'hf79a:	data_out=16'h2aa;
17'hf79b:	data_out=16'h9db;
17'hf79c:	data_out=16'h8a00;
17'hf79d:	data_out=16'h89ff;
17'hf79e:	data_out=16'h8989;
17'hf79f:	data_out=16'h4d2;
17'hf7a0:	data_out=16'h89f7;
17'hf7a1:	data_out=16'h922;
17'hf7a2:	data_out=16'h8713;
17'hf7a3:	data_out=16'ha00;
17'hf7a4:	data_out=16'ha00;
17'hf7a5:	data_out=16'h81d7;
17'hf7a6:	data_out=16'h865f;
17'hf7a7:	data_out=16'h194;
17'hf7a8:	data_out=16'h9f3;
17'hf7a9:	data_out=16'h89de;
17'hf7aa:	data_out=16'h9f8;
17'hf7ab:	data_out=16'ha00;
17'hf7ac:	data_out=16'h89d5;
17'hf7ad:	data_out=16'h89bf;
17'hf7ae:	data_out=16'h3b6;
17'hf7af:	data_out=16'h83f3;
17'hf7b0:	data_out=16'ha00;
17'hf7b1:	data_out=16'h8a00;
17'hf7b2:	data_out=16'h9c4;
17'hf7b3:	data_out=16'h89d5;
17'hf7b4:	data_out=16'h8a00;
17'hf7b5:	data_out=16'h70f;
17'hf7b6:	data_out=16'h9ef;
17'hf7b7:	data_out=16'h178;
17'hf7b8:	data_out=16'h8a00;
17'hf7b9:	data_out=16'h89e4;
17'hf7ba:	data_out=16'h9ff;
17'hf7bb:	data_out=16'ha00;
17'hf7bc:	data_out=16'h89f9;
17'hf7bd:	data_out=16'h89e5;
17'hf7be:	data_out=16'h9f3;
17'hf7bf:	data_out=16'h8a00;
17'hf7c0:	data_out=16'h84a;
17'hf7c1:	data_out=16'h924;
17'hf7c2:	data_out=16'h86f1;
17'hf7c3:	data_out=16'ha00;
17'hf7c4:	data_out=16'h89ed;
17'hf7c5:	data_out=16'h89f8;
17'hf7c6:	data_out=16'h89f7;
17'hf7c7:	data_out=16'h9ff;
17'hf7c8:	data_out=16'h207;
17'hf7c9:	data_out=16'h87;
17'hf7ca:	data_out=16'ha00;
17'hf7cb:	data_out=16'h822c;
17'hf7cc:	data_out=16'h81f6;
17'hf7cd:	data_out=16'h879d;
17'hf7ce:	data_out=16'ha00;
17'hf7cf:	data_out=16'h241;
17'hf7d0:	data_out=16'h8812;
17'hf7d1:	data_out=16'h8a00;
17'hf7d2:	data_out=16'ha00;
17'hf7d3:	data_out=16'h95e;
17'hf7d4:	data_out=16'h8834;
17'hf7d5:	data_out=16'h24e;
17'hf7d6:	data_out=16'h871b;
17'hf7d7:	data_out=16'h89d1;
17'hf7d8:	data_out=16'h89ff;
17'hf7d9:	data_out=16'h8951;
17'hf7da:	data_out=16'h89a3;
17'hf7db:	data_out=16'h89f3;
17'hf7dc:	data_out=16'h8a00;
17'hf7dd:	data_out=16'h860a;
17'hf7de:	data_out=16'h82ed;
17'hf7df:	data_out=16'h88f0;
17'hf7e0:	data_out=16'h89ae;
17'hf7e1:	data_out=16'h8a00;
17'hf7e2:	data_out=16'h48d;
17'hf7e3:	data_out=16'h89c9;
17'hf7e4:	data_out=16'h8a00;
17'hf7e5:	data_out=16'h4bd;
17'hf7e6:	data_out=16'ha00;
17'hf7e7:	data_out=16'ha00;
17'hf7e8:	data_out=16'h9f4;
17'hf7e9:	data_out=16'h9be;
17'hf7ea:	data_out=16'h544;
17'hf7eb:	data_out=16'h89d5;
17'hf7ec:	data_out=16'h8a00;
17'hf7ed:	data_out=16'h89cb;
17'hf7ee:	data_out=16'h54f;
17'hf7ef:	data_out=16'h1d0;
17'hf7f0:	data_out=16'h65e;
17'hf7f1:	data_out=16'h9ee;
17'hf7f2:	data_out=16'h8a00;
17'hf7f3:	data_out=16'h8a00;
17'hf7f4:	data_out=16'h9f6;
17'hf7f5:	data_out=16'h8a00;
17'hf7f6:	data_out=16'ha00;
17'hf7f7:	data_out=16'ha00;
17'hf7f8:	data_out=16'h881b;
17'hf7f9:	data_out=16'h9ba;
17'hf7fa:	data_out=16'h88ca;
17'hf7fb:	data_out=16'h9f3;
17'hf7fc:	data_out=16'h99c;
17'hf7fd:	data_out=16'h80a8;
17'hf7fe:	data_out=16'h89d3;
17'hf7ff:	data_out=16'h8a00;
17'hf800:	data_out=16'h8a00;
17'hf801:	data_out=16'h8a00;
17'hf802:	data_out=16'h81da;
17'hf803:	data_out=16'h89be;
17'hf804:	data_out=16'h9ff;
17'hf805:	data_out=16'h89ee;
17'hf806:	data_out=16'h8971;
17'hf807:	data_out=16'ha00;
17'hf808:	data_out=16'h9a2;
17'hf809:	data_out=16'hd9;
17'hf80a:	data_out=16'h8a00;
17'hf80b:	data_out=16'h809a;
17'hf80c:	data_out=16'h9ff;
17'hf80d:	data_out=16'h89d5;
17'hf80e:	data_out=16'hd4;
17'hf80f:	data_out=16'h9f9;
17'hf810:	data_out=16'h8591;
17'hf811:	data_out=16'h89ff;
17'hf812:	data_out=16'h89ec;
17'hf813:	data_out=16'h89c7;
17'hf814:	data_out=16'h89be;
17'hf815:	data_out=16'h89f6;
17'hf816:	data_out=16'h893b;
17'hf817:	data_out=16'h89be;
17'hf818:	data_out=16'h85ea;
17'hf819:	data_out=16'ha00;
17'hf81a:	data_out=16'h96d;
17'hf81b:	data_out=16'h83ca;
17'hf81c:	data_out=16'h8a00;
17'hf81d:	data_out=16'h8a00;
17'hf81e:	data_out=16'h89cc;
17'hf81f:	data_out=16'h8657;
17'hf820:	data_out=16'h89f4;
17'hf821:	data_out=16'h21c;
17'hf822:	data_out=16'h8745;
17'hf823:	data_out=16'h9ff;
17'hf824:	data_out=16'h9ff;
17'hf825:	data_out=16'h825d;
17'hf826:	data_out=16'h8763;
17'hf827:	data_out=16'h903;
17'hf828:	data_out=16'h41f;
17'hf829:	data_out=16'h8a00;
17'hf82a:	data_out=16'ha00;
17'hf82b:	data_out=16'ha00;
17'hf82c:	data_out=16'h89dc;
17'hf82d:	data_out=16'h8a00;
17'hf82e:	data_out=16'h2fa;
17'hf82f:	data_out=16'h8123;
17'hf830:	data_out=16'h9ff;
17'hf831:	data_out=16'h8a00;
17'hf832:	data_out=16'h9ec;
17'hf833:	data_out=16'h89e0;
17'hf834:	data_out=16'h8a00;
17'hf835:	data_out=16'h919;
17'hf836:	data_out=16'h9e3;
17'hf837:	data_out=16'h81b2;
17'hf838:	data_out=16'h8a00;
17'hf839:	data_out=16'h89ee;
17'hf83a:	data_out=16'h5e2;
17'hf83b:	data_out=16'ha00;
17'hf83c:	data_out=16'h8a00;
17'hf83d:	data_out=16'h89f4;
17'hf83e:	data_out=16'h42f;
17'hf83f:	data_out=16'h89f0;
17'hf840:	data_out=16'h9fb;
17'hf841:	data_out=16'h96b;
17'hf842:	data_out=16'h8490;
17'hf843:	data_out=16'h9ec;
17'hf844:	data_out=16'h8256;
17'hf845:	data_out=16'h89f5;
17'hf846:	data_out=16'h8a00;
17'hf847:	data_out=16'ha00;
17'hf848:	data_out=16'h8555;
17'hf849:	data_out=16'h8160;
17'hf84a:	data_out=16'ha00;
17'hf84b:	data_out=16'h9eb;
17'hf84c:	data_out=16'h8153;
17'hf84d:	data_out=16'h87c7;
17'hf84e:	data_out=16'ha00;
17'hf84f:	data_out=16'h58a;
17'hf850:	data_out=16'h85dd;
17'hf851:	data_out=16'h89dd;
17'hf852:	data_out=16'h9ff;
17'hf853:	data_out=16'h972;
17'hf854:	data_out=16'h883b;
17'hf855:	data_out=16'h8216;
17'hf856:	data_out=16'h936;
17'hf857:	data_out=16'h898d;
17'hf858:	data_out=16'h89f2;
17'hf859:	data_out=16'h85d0;
17'hf85a:	data_out=16'h89de;
17'hf85b:	data_out=16'h82f3;
17'hf85c:	data_out=16'h8a00;
17'hf85d:	data_out=16'h24;
17'hf85e:	data_out=16'h80a2;
17'hf85f:	data_out=16'h886d;
17'hf860:	data_out=16'h89dd;
17'hf861:	data_out=16'h89ff;
17'hf862:	data_out=16'h127;
17'hf863:	data_out=16'h89d8;
17'hf864:	data_out=16'h8a00;
17'hf865:	data_out=16'h970;
17'hf866:	data_out=16'ha00;
17'hf867:	data_out=16'ha00;
17'hf868:	data_out=16'h2de;
17'hf869:	data_out=16'h9b4;
17'hf86a:	data_out=16'h8073;
17'hf86b:	data_out=16'h8909;
17'hf86c:	data_out=16'h8a00;
17'hf86d:	data_out=16'h89da;
17'hf86e:	data_out=16'h806a;
17'hf86f:	data_out=16'h9aa;
17'hf870:	data_out=16'h67;
17'hf871:	data_out=16'h9f9;
17'hf872:	data_out=16'h89fd;
17'hf873:	data_out=16'h8a00;
17'hf874:	data_out=16'h9a1;
17'hf875:	data_out=16'h8a00;
17'hf876:	data_out=16'ha00;
17'hf877:	data_out=16'ha00;
17'hf878:	data_out=16'h8258;
17'hf879:	data_out=16'h9e6;
17'hf87a:	data_out=16'h89c8;
17'hf87b:	data_out=16'h438;
17'hf87c:	data_out=16'h87a;
17'hf87d:	data_out=16'h8659;
17'hf87e:	data_out=16'h89f3;
17'hf87f:	data_out=16'h89ff;
17'hf880:	data_out=16'h85af;
17'hf881:	data_out=16'h8a00;
17'hf882:	data_out=16'h12d;
17'hf883:	data_out=16'h89a3;
17'hf884:	data_out=16'ha00;
17'hf885:	data_out=16'h8806;
17'hf886:	data_out=16'h89eb;
17'hf887:	data_out=16'ha00;
17'hf888:	data_out=16'h9ce;
17'hf889:	data_out=16'h8127;
17'hf88a:	data_out=16'h89e1;
17'hf88b:	data_out=16'h9f7;
17'hf88c:	data_out=16'h9ee;
17'hf88d:	data_out=16'h89d5;
17'hf88e:	data_out=16'h826d;
17'hf88f:	data_out=16'ha00;
17'hf890:	data_out=16'h89f2;
17'hf891:	data_out=16'h9b3;
17'hf892:	data_out=16'h88fd;
17'hf893:	data_out=16'h89cb;
17'hf894:	data_out=16'h894f;
17'hf895:	data_out=16'h85d5;
17'hf896:	data_out=16'h8279;
17'hf897:	data_out=16'h8953;
17'hf898:	data_out=16'h868f;
17'hf899:	data_out=16'h9ff;
17'hf89a:	data_out=16'h9e4;
17'hf89b:	data_out=16'h85bc;
17'hf89c:	data_out=16'h8a00;
17'hf89d:	data_out=16'h8257;
17'hf89e:	data_out=16'h8731;
17'hf89f:	data_out=16'h1d5;
17'hf8a0:	data_out=16'h105;
17'hf8a1:	data_out=16'h81e2;
17'hf8a2:	data_out=16'h8992;
17'hf8a3:	data_out=16'h22a;
17'hf8a4:	data_out=16'h257;
17'hf8a5:	data_out=16'h8495;
17'hf8a6:	data_out=16'h86aa;
17'hf8a7:	data_out=16'h9dc;
17'hf8a8:	data_out=16'h80ff;
17'hf8a9:	data_out=16'h89c3;
17'hf8aa:	data_out=16'ha00;
17'hf8ab:	data_out=16'ha00;
17'hf8ac:	data_out=16'h8455;
17'hf8ad:	data_out=16'h8a00;
17'hf8ae:	data_out=16'h79c;
17'hf8af:	data_out=16'h3e2;
17'hf8b0:	data_out=16'h8390;
17'hf8b1:	data_out=16'h89f5;
17'hf8b2:	data_out=16'h79;
17'hf8b3:	data_out=16'h89ec;
17'hf8b4:	data_out=16'h8a00;
17'hf8b5:	data_out=16'h9e5;
17'hf8b6:	data_out=16'h9e7;
17'hf8b7:	data_out=16'h1f7;
17'hf8b8:	data_out=16'h8a00;
17'hf8b9:	data_out=16'h89f5;
17'hf8ba:	data_out=16'h18d;
17'hf8bb:	data_out=16'ha00;
17'hf8bc:	data_out=16'h89f8;
17'hf8bd:	data_out=16'h8308;
17'hf8be:	data_out=16'h80f4;
17'hf8bf:	data_out=16'h8848;
17'hf8c0:	data_out=16'ha00;
17'hf8c1:	data_out=16'h9ca;
17'hf8c2:	data_out=16'h82f0;
17'hf8c3:	data_out=16'h9fb;
17'hf8c4:	data_out=16'ha00;
17'hf8c5:	data_out=16'h8595;
17'hf8c6:	data_out=16'h8a00;
17'hf8c7:	data_out=16'h9f9;
17'hf8c8:	data_out=16'h47e;
17'hf8c9:	data_out=16'h8527;
17'hf8ca:	data_out=16'ha00;
17'hf8cb:	data_out=16'h9d5;
17'hf8cc:	data_out=16'h8533;
17'hf8cd:	data_out=16'h89f7;
17'hf8ce:	data_out=16'ha00;
17'hf8cf:	data_out=16'h556;
17'hf8d0:	data_out=16'h87a1;
17'hf8d1:	data_out=16'h89c8;
17'hf8d2:	data_out=16'h80c4;
17'hf8d3:	data_out=16'h9e3;
17'hf8d4:	data_out=16'h27c;
17'hf8d5:	data_out=16'h82e8;
17'hf8d6:	data_out=16'h9ec;
17'hf8d7:	data_out=16'h8778;
17'hf8d8:	data_out=16'h89ed;
17'hf8d9:	data_out=16'h8052;
17'hf8da:	data_out=16'h89eb;
17'hf8db:	data_out=16'ha00;
17'hf8dc:	data_out=16'h89fb;
17'hf8dd:	data_out=16'h988;
17'hf8de:	data_out=16'h4b7;
17'hf8df:	data_out=16'h8609;
17'hf8e0:	data_out=16'h898e;
17'hf8e1:	data_out=16'h789;
17'hf8e2:	data_out=16'h15a;
17'hf8e3:	data_out=16'h89b5;
17'hf8e4:	data_out=16'h8a00;
17'hf8e5:	data_out=16'h9ea;
17'hf8e6:	data_out=16'ha00;
17'hf8e7:	data_out=16'ha00;
17'hf8e8:	data_out=16'h8191;
17'hf8e9:	data_out=16'h9e3;
17'hf8ea:	data_out=16'h8326;
17'hf8eb:	data_out=16'h972;
17'hf8ec:	data_out=16'h834a;
17'hf8ed:	data_out=16'h89c3;
17'hf8ee:	data_out=16'h8321;
17'hf8ef:	data_out=16'h6c2;
17'hf8f0:	data_out=16'h82a9;
17'hf8f1:	data_out=16'ha00;
17'hf8f2:	data_out=16'h89f2;
17'hf8f3:	data_out=16'h89cb;
17'hf8f4:	data_out=16'h86d6;
17'hf8f5:	data_out=16'h89fe;
17'hf8f6:	data_out=16'ha00;
17'hf8f7:	data_out=16'ha00;
17'hf8f8:	data_out=16'h8202;
17'hf8f9:	data_out=16'h9f5;
17'hf8fa:	data_out=16'h891e;
17'hf8fb:	data_out=16'h80ef;
17'hf8fc:	data_out=16'h8085;
17'hf8fd:	data_out=16'h73e;
17'hf8fe:	data_out=16'h8a00;
17'hf8ff:	data_out=16'h89fe;
17'hf900:	data_out=16'h89f3;
17'hf901:	data_out=16'h7a1;
17'hf902:	data_out=16'h89e4;
17'hf903:	data_out=16'h89f9;
17'hf904:	data_out=16'ha00;
17'hf905:	data_out=16'h8583;
17'hf906:	data_out=16'h89fd;
17'hf907:	data_out=16'h9f0;
17'hf908:	data_out=16'h47d;
17'hf909:	data_out=16'h851e;
17'hf90a:	data_out=16'h9ef;
17'hf90b:	data_out=16'h9e7;
17'hf90c:	data_out=16'h9c7;
17'hf90d:	data_out=16'h89ff;
17'hf90e:	data_out=16'h89f5;
17'hf90f:	data_out=16'h84c9;
17'hf910:	data_out=16'h89fa;
17'hf911:	data_out=16'h9e1;
17'hf912:	data_out=16'h89fd;
17'hf913:	data_out=16'h89f8;
17'hf914:	data_out=16'h89e9;
17'hf915:	data_out=16'h89b5;
17'hf916:	data_out=16'h8941;
17'hf917:	data_out=16'h89f0;
17'hf918:	data_out=16'h89fb;
17'hf919:	data_out=16'ha00;
17'hf91a:	data_out=16'ha00;
17'hf91b:	data_out=16'h89e7;
17'hf91c:	data_out=16'h8a00;
17'hf91d:	data_out=16'h8e8;
17'hf91e:	data_out=16'h89f2;
17'hf91f:	data_out=16'h81dd;
17'hf920:	data_out=16'h8335;
17'hf921:	data_out=16'h89f5;
17'hf922:	data_out=16'h840f;
17'hf923:	data_out=16'h894b;
17'hf924:	data_out=16'h893e;
17'hf925:	data_out=16'h89f0;
17'hf926:	data_out=16'h89c9;
17'hf927:	data_out=16'h9ef;
17'hf928:	data_out=16'h89f5;
17'hf929:	data_out=16'h89fa;
17'hf92a:	data_out=16'h207;
17'hf92b:	data_out=16'ha00;
17'hf92c:	data_out=16'h8982;
17'hf92d:	data_out=16'h8a00;
17'hf92e:	data_out=16'h8369;
17'hf92f:	data_out=16'h8460;
17'hf930:	data_out=16'h83c6;
17'hf931:	data_out=16'h88b;
17'hf932:	data_out=16'h160;
17'hf933:	data_out=16'h89f2;
17'hf934:	data_out=16'h8a00;
17'hf935:	data_out=16'h9e7;
17'hf936:	data_out=16'h8527;
17'hf937:	data_out=16'h89e1;
17'hf938:	data_out=16'h8a00;
17'hf939:	data_out=16'h89fa;
17'hf93a:	data_out=16'h81df;
17'hf93b:	data_out=16'h9ff;
17'hf93c:	data_out=16'h89f6;
17'hf93d:	data_out=16'h895c;
17'hf93e:	data_out=16'h89f5;
17'hf93f:	data_out=16'h8609;
17'hf940:	data_out=16'ha00;
17'hf941:	data_out=16'h84b7;
17'hf942:	data_out=16'h9ce;
17'hf943:	data_out=16'h801;
17'hf944:	data_out=16'ha00;
17'hf945:	data_out=16'h89a2;
17'hf946:	data_out=16'h8a00;
17'hf947:	data_out=16'h9cf;
17'hf948:	data_out=16'h781;
17'hf949:	data_out=16'h89f0;
17'hf94a:	data_out=16'h9fc;
17'hf94b:	data_out=16'h9c4;
17'hf94c:	data_out=16'h674;
17'hf94d:	data_out=16'h8502;
17'hf94e:	data_out=16'h569;
17'hf94f:	data_out=16'h872;
17'hf950:	data_out=16'h89f0;
17'hf951:	data_out=16'h89e4;
17'hf952:	data_out=16'h8536;
17'hf953:	data_out=16'ha00;
17'hf954:	data_out=16'h84a4;
17'hf955:	data_out=16'h899d;
17'hf956:	data_out=16'h8803;
17'hf957:	data_out=16'h89db;
17'hf958:	data_out=16'h89f9;
17'hf959:	data_out=16'h667;
17'hf95a:	data_out=16'h89f5;
17'hf95b:	data_out=16'ha00;
17'hf95c:	data_out=16'h239;
17'hf95d:	data_out=16'h82eb;
17'hf95e:	data_out=16'h8307;
17'hf95f:	data_out=16'h88c0;
17'hf960:	data_out=16'h89e9;
17'hf961:	data_out=16'h9fb;
17'hf962:	data_out=16'h8641;
17'hf963:	data_out=16'h89ee;
17'hf964:	data_out=16'h2dc;
17'hf965:	data_out=16'h9e8;
17'hf966:	data_out=16'ha00;
17'hf967:	data_out=16'ha00;
17'hf968:	data_out=16'h89f4;
17'hf969:	data_out=16'h8ad;
17'hf96a:	data_out=16'h89f5;
17'hf96b:	data_out=16'h9c6;
17'hf96c:	data_out=16'h89f3;
17'hf96d:	data_out=16'h89f0;
17'hf96e:	data_out=16'h89f5;
17'hf96f:	data_out=16'h7bf;
17'hf970:	data_out=16'h89f5;
17'hf971:	data_out=16'h824c;
17'hf972:	data_out=16'h89f8;
17'hf973:	data_out=16'h8563;
17'hf974:	data_out=16'h8861;
17'hf975:	data_out=16'h89e3;
17'hf976:	data_out=16'ha00;
17'hf977:	data_out=16'h8499;
17'hf978:	data_out=16'h88eb;
17'hf979:	data_out=16'h661;
17'hf97a:	data_out=16'h89ed;
17'hf97b:	data_out=16'h89f5;
17'hf97c:	data_out=16'h89e4;
17'hf97d:	data_out=16'h14;
17'hf97e:	data_out=16'h8a00;
17'hf97f:	data_out=16'h89ff;
17'hf980:	data_out=16'h89ed;
17'hf981:	data_out=16'h88c;
17'hf982:	data_out=16'h89ef;
17'hf983:	data_out=16'h8a00;
17'hf984:	data_out=16'ha00;
17'hf985:	data_out=16'h422;
17'hf986:	data_out=16'h89fd;
17'hf987:	data_out=16'h9de;
17'hf988:	data_out=16'h89ec;
17'hf989:	data_out=16'h87eb;
17'hf98a:	data_out=16'h9ff;
17'hf98b:	data_out=16'h9c9;
17'hf98c:	data_out=16'h283;
17'hf98d:	data_out=16'h89ff;
17'hf98e:	data_out=16'h8460;
17'hf98f:	data_out=16'h89ed;
17'hf990:	data_out=16'h8a00;
17'hf991:	data_out=16'h9f3;
17'hf992:	data_out=16'h89ff;
17'hf993:	data_out=16'h89f3;
17'hf994:	data_out=16'h8a00;
17'hf995:	data_out=16'h8595;
17'hf996:	data_out=16'h89fc;
17'hf997:	data_out=16'h8a00;
17'hf998:	data_out=16'h89f5;
17'hf999:	data_out=16'ha00;
17'hf99a:	data_out=16'ha00;
17'hf99b:	data_out=16'h8a00;
17'hf99c:	data_out=16'h8a00;
17'hf99d:	data_out=16'h986;
17'hf99e:	data_out=16'h89ff;
17'hf99f:	data_out=16'h845a;
17'hf9a0:	data_out=16'h7bf;
17'hf9a1:	data_out=16'h84d1;
17'hf9a2:	data_out=16'h8af;
17'hf9a3:	data_out=16'h7bf;
17'hf9a4:	data_out=16'h7dd;
17'hf9a5:	data_out=16'h89e7;
17'hf9a6:	data_out=16'h89fc;
17'hf9a7:	data_out=16'h9f1;
17'hf9a8:	data_out=16'h85a9;
17'hf9a9:	data_out=16'h8a00;
17'hf9aa:	data_out=16'h89e1;
17'hf9ab:	data_out=16'ha00;
17'hf9ac:	data_out=16'h89fb;
17'hf9ad:	data_out=16'h8a00;
17'hf9ae:	data_out=16'h89f2;
17'hf9af:	data_out=16'h89ff;
17'hf9b0:	data_out=16'h8042;
17'hf9b1:	data_out=16'h9e1;
17'hf9b2:	data_out=16'h5c7;
17'hf9b3:	data_out=16'h8a00;
17'hf9b4:	data_out=16'h53d;
17'hf9b5:	data_out=16'h9ff;
17'hf9b6:	data_out=16'h89ec;
17'hf9b7:	data_out=16'h89ee;
17'hf9b8:	data_out=16'h26b;
17'hf9b9:	data_out=16'h8a00;
17'hf9ba:	data_out=16'h8279;
17'hf9bb:	data_out=16'ha00;
17'hf9bc:	data_out=16'h89f8;
17'hf9bd:	data_out=16'h188;
17'hf9be:	data_out=16'h85b2;
17'hf9bf:	data_out=16'h3f8;
17'hf9c0:	data_out=16'ha00;
17'hf9c1:	data_out=16'h89f4;
17'hf9c2:	data_out=16'h9c7;
17'hf9c3:	data_out=16'h8704;
17'hf9c4:	data_out=16'ha00;
17'hf9c5:	data_out=16'h866c;
17'hf9c6:	data_out=16'h8a00;
17'hf9c7:	data_out=16'h369;
17'hf9c8:	data_out=16'h84c4;
17'hf9c9:	data_out=16'h89e9;
17'hf9ca:	data_out=16'h9e5;
17'hf9cb:	data_out=16'h9cb;
17'hf9cc:	data_out=16'h868a;
17'hf9cd:	data_out=16'h852;
17'hf9ce:	data_out=16'h1ab;
17'hf9cf:	data_out=16'h8722;
17'hf9d0:	data_out=16'h89f7;
17'hf9d1:	data_out=16'h89f6;
17'hf9d2:	data_out=16'h9d9;
17'hf9d3:	data_out=16'h9f6;
17'hf9d4:	data_out=16'h881a;
17'hf9d5:	data_out=16'h89f6;
17'hf9d6:	data_out=16'h89f2;
17'hf9d7:	data_out=16'h89cf;
17'hf9d8:	data_out=16'h8a00;
17'hf9d9:	data_out=16'ha00;
17'hf9da:	data_out=16'h8a00;
17'hf9db:	data_out=16'ha00;
17'hf9dc:	data_out=16'h3ce;
17'hf9dd:	data_out=16'h89ee;
17'hf9de:	data_out=16'h8a00;
17'hf9df:	data_out=16'h8920;
17'hf9e0:	data_out=16'h89fe;
17'hf9e1:	data_out=16'h9ff;
17'hf9e2:	data_out=16'h8a00;
17'hf9e3:	data_out=16'h8a00;
17'hf9e4:	data_out=16'h9bb;
17'hf9e5:	data_out=16'h9e9;
17'hf9e6:	data_out=16'ha00;
17'hf9e7:	data_out=16'ha00;
17'hf9e8:	data_out=16'h8515;
17'hf9e9:	data_out=16'h89fd;
17'hf9ea:	data_out=16'h841a;
17'hf9eb:	data_out=16'h961;
17'hf9ec:	data_out=16'h89ea;
17'hf9ed:	data_out=16'h8a00;
17'hf9ee:	data_out=16'h841c;
17'hf9ef:	data_out=16'h8370;
17'hf9f0:	data_out=16'h8447;
17'hf9f1:	data_out=16'h89d9;
17'hf9f2:	data_out=16'h8df;
17'hf9f3:	data_out=16'h9d8;
17'hf9f4:	data_out=16'h8499;
17'hf9f5:	data_out=16'h89dc;
17'hf9f6:	data_out=16'ha00;
17'hf9f7:	data_out=16'h89f7;
17'hf9f8:	data_out=16'h89e3;
17'hf9f9:	data_out=16'h8534;
17'hf9fa:	data_out=16'h8a00;
17'hf9fb:	data_out=16'h85b5;
17'hf9fc:	data_out=16'h89e5;
17'hf9fd:	data_out=16'h174;
17'hf9fe:	data_out=16'h8a00;
17'hf9ff:	data_out=16'h89df;
17'hfa00:	data_out=16'ha00;
17'hfa01:	data_out=16'h9fb;
17'hfa02:	data_out=16'h8a00;
17'hfa03:	data_out=16'h8a00;
17'hfa04:	data_out=16'ha00;
17'hfa05:	data_out=16'h8d4;
17'hfa06:	data_out=16'h89fc;
17'hfa07:	data_out=16'h8a00;
17'hfa08:	data_out=16'h8a00;
17'hfa09:	data_out=16'h86b;
17'hfa0a:	data_out=16'ha00;
17'hfa0b:	data_out=16'h8629;
17'hfa0c:	data_out=16'h8a00;
17'hfa0d:	data_out=16'h8a00;
17'hfa0e:	data_out=16'h838f;
17'hfa0f:	data_out=16'h8a00;
17'hfa10:	data_out=16'h934;
17'hfa11:	data_out=16'ha00;
17'hfa12:	data_out=16'h8a00;
17'hfa13:	data_out=16'h89f7;
17'hfa14:	data_out=16'h8a00;
17'hfa15:	data_out=16'ha00;
17'hfa16:	data_out=16'h81c9;
17'hfa17:	data_out=16'h8a00;
17'hfa18:	data_out=16'h89ec;
17'hfa19:	data_out=16'ha00;
17'hfa1a:	data_out=16'ha00;
17'hfa1b:	data_out=16'h8a00;
17'hfa1c:	data_out=16'h273;
17'hfa1d:	data_out=16'ha00;
17'hfa1e:	data_out=16'h8a00;
17'hfa1f:	data_out=16'h870f;
17'hfa20:	data_out=16'ha00;
17'hfa21:	data_out=16'h8423;
17'hfa22:	data_out=16'h9f1;
17'hfa23:	data_out=16'h8796;
17'hfa24:	data_out=16'h877c;
17'hfa25:	data_out=16'h8b;
17'hfa26:	data_out=16'h8a00;
17'hfa27:	data_out=16'ha00;
17'hfa28:	data_out=16'h852a;
17'hfa29:	data_out=16'h8a00;
17'hfa2a:	data_out=16'h89ff;
17'hfa2b:	data_out=16'ha00;
17'hfa2c:	data_out=16'h975;
17'hfa2d:	data_out=16'h84d7;
17'hfa2e:	data_out=16'h8a00;
17'hfa2f:	data_out=16'h8ff;
17'hfa30:	data_out=16'h838f;
17'hfa31:	data_out=16'ha00;
17'hfa32:	data_out=16'h655;
17'hfa33:	data_out=16'h8a00;
17'hfa34:	data_out=16'h9ee;
17'hfa35:	data_out=16'ha00;
17'hfa36:	data_out=16'h89fe;
17'hfa37:	data_out=16'h8a00;
17'hfa38:	data_out=16'ha00;
17'hfa39:	data_out=16'h89fd;
17'hfa3a:	data_out=16'h9cc;
17'hfa3b:	data_out=16'h7a1;
17'hfa3c:	data_out=16'h8a00;
17'hfa3d:	data_out=16'ha00;
17'hfa3e:	data_out=16'h8536;
17'hfa3f:	data_out=16'h8e4;
17'hfa40:	data_out=16'ha00;
17'hfa41:	data_out=16'h8a00;
17'hfa42:	data_out=16'h82e2;
17'hfa43:	data_out=16'h89f4;
17'hfa44:	data_out=16'ha00;
17'hfa45:	data_out=16'ha00;
17'hfa46:	data_out=16'h8a00;
17'hfa47:	data_out=16'h9e4;
17'hfa48:	data_out=16'h89e7;
17'hfa49:	data_out=16'h463;
17'hfa4a:	data_out=16'h8748;
17'hfa4b:	data_out=16'h1c;
17'hfa4c:	data_out=16'h837e;
17'hfa4d:	data_out=16'h9fd;
17'hfa4e:	data_out=16'h859e;
17'hfa4f:	data_out=16'h3ae;
17'hfa50:	data_out=16'h948;
17'hfa51:	data_out=16'h8a00;
17'hfa52:	data_out=16'h869;
17'hfa53:	data_out=16'h83c6;
17'hfa54:	data_out=16'ha00;
17'hfa55:	data_out=16'h8a00;
17'hfa56:	data_out=16'h1a2;
17'hfa57:	data_out=16'ha00;
17'hfa58:	data_out=16'h8a00;
17'hfa59:	data_out=16'ha00;
17'hfa5a:	data_out=16'h8a00;
17'hfa5b:	data_out=16'ha00;
17'hfa5c:	data_out=16'h1fc;
17'hfa5d:	data_out=16'h606;
17'hfa5e:	data_out=16'h877;
17'hfa5f:	data_out=16'h85d;
17'hfa60:	data_out=16'h8a00;
17'hfa61:	data_out=16'h9ff;
17'hfa62:	data_out=16'h8a00;
17'hfa63:	data_out=16'h8a00;
17'hfa64:	data_out=16'ha00;
17'hfa65:	data_out=16'ha00;
17'hfa66:	data_out=16'ha00;
17'hfa67:	data_out=16'h9fe;
17'hfa68:	data_out=16'h8477;
17'hfa69:	data_out=16'h8a00;
17'hfa6a:	data_out=16'h832c;
17'hfa6b:	data_out=16'ha00;
17'hfa6c:	data_out=16'ha00;
17'hfa6d:	data_out=16'h8a00;
17'hfa6e:	data_out=16'h832f;
17'hfa6f:	data_out=16'h8945;
17'hfa70:	data_out=16'h836f;
17'hfa71:	data_out=16'h8a00;
17'hfa72:	data_out=16'ha00;
17'hfa73:	data_out=16'ha00;
17'hfa74:	data_out=16'h886e;
17'hfa75:	data_out=16'h89fb;
17'hfa76:	data_out=16'ha00;
17'hfa77:	data_out=16'h619;
17'hfa78:	data_out=16'h89cd;
17'hfa79:	data_out=16'h8969;
17'hfa7a:	data_out=16'h8a00;
17'hfa7b:	data_out=16'h853c;
17'hfa7c:	data_out=16'h806e;
17'hfa7d:	data_out=16'h7d;
17'hfa7e:	data_out=16'h66a;
17'hfa7f:	data_out=16'ha00;
17'hfa80:	data_out=16'ha00;
17'hfa81:	data_out=16'ha00;
17'hfa82:	data_out=16'h8a00;
17'hfa83:	data_out=16'h93d;
17'hfa84:	data_out=16'ha00;
17'hfa85:	data_out=16'h9aa;
17'hfa86:	data_out=16'ha00;
17'hfa87:	data_out=16'h8a00;
17'hfa88:	data_out=16'h8a00;
17'hfa89:	data_out=16'ha00;
17'hfa8a:	data_out=16'ha00;
17'hfa8b:	data_out=16'h83db;
17'hfa8c:	data_out=16'h8a00;
17'hfa8d:	data_out=16'h8a00;
17'hfa8e:	data_out=16'h8563;
17'hfa8f:	data_out=16'h8a00;
17'hfa90:	data_out=16'ha00;
17'hfa91:	data_out=16'ha00;
17'hfa92:	data_out=16'h8a00;
17'hfa93:	data_out=16'h9b6;
17'hfa94:	data_out=16'h589;
17'hfa95:	data_out=16'ha00;
17'hfa96:	data_out=16'h5cc;
17'hfa97:	data_out=16'h8a00;
17'hfa98:	data_out=16'h845a;
17'hfa99:	data_out=16'ha00;
17'hfa9a:	data_out=16'ha00;
17'hfa9b:	data_out=16'h8a00;
17'hfa9c:	data_out=16'h8e2;
17'hfa9d:	data_out=16'ha00;
17'hfa9e:	data_out=16'h8c4;
17'hfa9f:	data_out=16'ha00;
17'hfaa0:	data_out=16'ha00;
17'hfaa1:	data_out=16'h857b;
17'hfaa2:	data_out=16'ha00;
17'hfaa3:	data_out=16'h8a00;
17'hfaa4:	data_out=16'h8a00;
17'hfaa5:	data_out=16'ha00;
17'hfaa6:	data_out=16'h8a00;
17'hfaa7:	data_out=16'ha00;
17'hfaa8:	data_out=16'h858d;
17'hfaa9:	data_out=16'h83b8;
17'hfaaa:	data_out=16'h8a00;
17'hfaab:	data_out=16'ha00;
17'hfaac:	data_out=16'ha00;
17'hfaad:	data_out=16'h8e8;
17'hfaae:	data_out=16'h8a00;
17'hfaaf:	data_out=16'ha00;
17'hfab0:	data_out=16'h8a00;
17'hfab1:	data_out=16'ha00;
17'hfab2:	data_out=16'h8518;
17'hfab3:	data_out=16'ha00;
17'hfab4:	data_out=16'ha00;
17'hfab5:	data_out=16'ha00;
17'hfab6:	data_out=16'h8777;
17'hfab7:	data_out=16'h8a00;
17'hfab8:	data_out=16'ha00;
17'hfab9:	data_out=16'ha00;
17'hfaba:	data_out=16'ha00;
17'hfabb:	data_out=16'h8207;
17'hfabc:	data_out=16'h8a00;
17'hfabd:	data_out=16'ha00;
17'hfabe:	data_out=16'h8590;
17'hfabf:	data_out=16'h9b0;
17'hfac0:	data_out=16'ha00;
17'hfac1:	data_out=16'h8a00;
17'hfac2:	data_out=16'h898a;
17'hfac3:	data_out=16'ha00;
17'hfac4:	data_out=16'ha00;
17'hfac5:	data_out=16'ha00;
17'hfac6:	data_out=16'h8a00;
17'hfac7:	data_out=16'ha00;
17'hfac8:	data_out=16'ha00;
17'hfac9:	data_out=16'ha00;
17'hfaca:	data_out=16'h8792;
17'hfacb:	data_out=16'h8944;
17'hfacc:	data_out=16'h4f2;
17'hfacd:	data_out=16'ha00;
17'hface:	data_out=16'h8a00;
17'hfacf:	data_out=16'h9fd;
17'hfad0:	data_out=16'ha00;
17'hfad1:	data_out=16'h8a00;
17'hfad2:	data_out=16'h8797;
17'hfad3:	data_out=16'ha00;
17'hfad4:	data_out=16'ha00;
17'hfad5:	data_out=16'h8a00;
17'hfad6:	data_out=16'h93c;
17'hfad7:	data_out=16'ha00;
17'hfad8:	data_out=16'h8a00;
17'hfad9:	data_out=16'ha00;
17'hfada:	data_out=16'h8a00;
17'hfadb:	data_out=16'ha00;
17'hfadc:	data_out=16'h60c;
17'hfadd:	data_out=16'ha00;
17'hfade:	data_out=16'ha00;
17'hfadf:	data_out=16'ha00;
17'hfae0:	data_out=16'h8a00;
17'hfae1:	data_out=16'ha00;
17'hfae2:	data_out=16'h89ff;
17'hfae3:	data_out=16'ha00;
17'hfae4:	data_out=16'ha00;
17'hfae5:	data_out=16'ha00;
17'hfae6:	data_out=16'ha00;
17'hfae7:	data_out=16'ha00;
17'hfae8:	data_out=16'h8578;
17'hfae9:	data_out=16'h8a00;
17'hfaea:	data_out=16'h8551;
17'hfaeb:	data_out=16'ha00;
17'hfaec:	data_out=16'ha00;
17'hfaed:	data_out=16'ha00;
17'hfaee:	data_out=16'h8553;
17'hfaef:	data_out=16'h857;
17'hfaf0:	data_out=16'h8566;
17'hfaf1:	data_out=16'h8a00;
17'hfaf2:	data_out=16'ha00;
17'hfaf3:	data_out=16'ha00;
17'hfaf4:	data_out=16'h8a00;
17'hfaf5:	data_out=16'h8a00;
17'hfaf6:	data_out=16'ha00;
17'hfaf7:	data_out=16'h9f9;
17'hfaf8:	data_out=16'h9e1;
17'hfaf9:	data_out=16'h8a00;
17'hfafa:	data_out=16'h9f2;
17'hfafb:	data_out=16'h8592;
17'hfafc:	data_out=16'he2;
17'hfafd:	data_out=16'ha00;
17'hfafe:	data_out=16'ha00;
17'hfaff:	data_out=16'ha00;
17'hfb00:	data_out=16'ha00;
17'hfb01:	data_out=16'ha00;
17'hfb02:	data_out=16'h89ed;
17'hfb03:	data_out=16'h7b6;
17'hfb04:	data_out=16'ha00;
17'hfb05:	data_out=16'h8fe;
17'hfb06:	data_out=16'h8102;
17'hfb07:	data_out=16'h82d0;
17'hfb08:	data_out=16'h88e5;
17'hfb09:	data_out=16'ha00;
17'hfb0a:	data_out=16'ha00;
17'hfb0b:	data_out=16'h865f;
17'hfb0c:	data_out=16'h8a00;
17'hfb0d:	data_out=16'h84a8;
17'hfb0e:	data_out=16'h8229;
17'hfb0f:	data_out=16'h8832;
17'hfb10:	data_out=16'ha00;
17'hfb11:	data_out=16'ha00;
17'hfb12:	data_out=16'h829e;
17'hfb13:	data_out=16'h33e;
17'hfb14:	data_out=16'h65e;
17'hfb15:	data_out=16'h696;
17'hfb16:	data_out=16'h35;
17'hfb17:	data_out=16'h77;
17'hfb18:	data_out=16'h80b3;
17'hfb19:	data_out=16'h56f;
17'hfb1a:	data_out=16'h6a0;
17'hfb1b:	data_out=16'h2a4;
17'hfb1c:	data_out=16'h9b0;
17'hfb1d:	data_out=16'ha00;
17'hfb1e:	data_out=16'h781;
17'hfb1f:	data_out=16'h534;
17'hfb20:	data_out=16'ha00;
17'hfb21:	data_out=16'h8237;
17'hfb22:	data_out=16'ha00;
17'hfb23:	data_out=16'h8839;
17'hfb24:	data_out=16'h8834;
17'hfb25:	data_out=16'h247;
17'hfb26:	data_out=16'h8155;
17'hfb27:	data_out=16'ha00;
17'hfb28:	data_out=16'h8235;
17'hfb29:	data_out=16'h7a7;
17'hfb2a:	data_out=16'h8978;
17'hfb2b:	data_out=16'ha00;
17'hfb2c:	data_out=16'h2c3;
17'hfb2d:	data_out=16'h2ff;
17'hfb2e:	data_out=16'h85bc;
17'hfb2f:	data_out=16'ha00;
17'hfb30:	data_out=16'h8a00;
17'hfb31:	data_out=16'ha00;
17'hfb32:	data_out=16'h8a00;
17'hfb33:	data_out=16'ha00;
17'hfb34:	data_out=16'ha00;
17'hfb35:	data_out=16'h844c;
17'hfb36:	data_out=16'h18;
17'hfb37:	data_out=16'h89eb;
17'hfb38:	data_out=16'ha00;
17'hfb39:	data_out=16'ha00;
17'hfb3a:	data_out=16'ha00;
17'hfb3b:	data_out=16'h3bb;
17'hfb3c:	data_out=16'h8a00;
17'hfb3d:	data_out=16'ha00;
17'hfb3e:	data_out=16'h823f;
17'hfb3f:	data_out=16'h87b;
17'hfb40:	data_out=16'h4f0;
17'hfb41:	data_out=16'h8a00;
17'hfb42:	data_out=16'h88b2;
17'hfb43:	data_out=16'h8123;
17'hfb44:	data_out=16'ha00;
17'hfb45:	data_out=16'h67f;
17'hfb46:	data_out=16'h81d5;
17'hfb47:	data_out=16'h4de;
17'hfb48:	data_out=16'h325;
17'hfb49:	data_out=16'h326;
17'hfb4a:	data_out=16'h856a;
17'hfb4b:	data_out=16'h8a00;
17'hfb4c:	data_out=16'h846e;
17'hfb4d:	data_out=16'ha00;
17'hfb4e:	data_out=16'h86fa;
17'hfb4f:	data_out=16'h81bb;
17'hfb50:	data_out=16'h50f;
17'hfb51:	data_out=16'h8a00;
17'hfb52:	data_out=16'h8648;
17'hfb53:	data_out=16'ha00;
17'hfb54:	data_out=16'ha00;
17'hfb55:	data_out=16'h8a00;
17'hfb56:	data_out=16'h5fb;
17'hfb57:	data_out=16'h8ec;
17'hfb58:	data_out=16'h8a00;
17'hfb59:	data_out=16'h647;
17'hfb5a:	data_out=16'h84ce;
17'hfb5b:	data_out=16'ha00;
17'hfb5c:	data_out=16'h943;
17'hfb5d:	data_out=16'h31c;
17'hfb5e:	data_out=16'ha00;
17'hfb5f:	data_out=16'h345;
17'hfb60:	data_out=16'h83a0;
17'hfb61:	data_out=16'h9f1;
17'hfb62:	data_out=16'h8a00;
17'hfb63:	data_out=16'ha00;
17'hfb64:	data_out=16'ha00;
17'hfb65:	data_out=16'ha00;
17'hfb66:	data_out=16'h551;
17'hfb67:	data_out=16'h4f1;
17'hfb68:	data_out=16'h8239;
17'hfb69:	data_out=16'h8a00;
17'hfb6a:	data_out=16'h8222;
17'hfb6b:	data_out=16'ha00;
17'hfb6c:	data_out=16'h804;
17'hfb6d:	data_out=16'ha00;
17'hfb6e:	data_out=16'h8223;
17'hfb6f:	data_out=16'h90;
17'hfb70:	data_out=16'h8228;
17'hfb71:	data_out=16'h89a8;
17'hfb72:	data_out=16'ha00;
17'hfb73:	data_out=16'ha00;
17'hfb74:	data_out=16'h8a00;
17'hfb75:	data_out=16'h8a00;
17'hfb76:	data_out=16'ha00;
17'hfb77:	data_out=16'h4d2;
17'hfb78:	data_out=16'h8170;
17'hfb79:	data_out=16'h8a00;
17'hfb7a:	data_out=16'h7b5;
17'hfb7b:	data_out=16'h822b;
17'hfb7c:	data_out=16'hc1;
17'hfb7d:	data_out=16'h195;
17'hfb7e:	data_out=16'ha00;
17'hfb7f:	data_out=16'h6a6;
17'hfb80:	data_out=16'h48e;
17'hfb81:	data_out=16'h217;
17'hfb82:	data_out=16'h832f;
17'hfb83:	data_out=16'h8249;
17'hfb84:	data_out=16'h8033;
17'hfb85:	data_out=16'h81b2;
17'hfb86:	data_out=16'h8253;
17'hfb87:	data_out=16'h8133;
17'hfb88:	data_out=16'h53;
17'hfb89:	data_out=16'h187;
17'hfb8a:	data_out=16'h312;
17'hfb8b:	data_out=16'h812b;
17'hfb8c:	data_out=16'h81f5;
17'hfb8d:	data_out=16'h82a4;
17'hfb8e:	data_out=16'h80b2;
17'hfb8f:	data_out=16'h82a8;
17'hfb90:	data_out=16'h808c;
17'hfb91:	data_out=16'h28a;
17'hfb92:	data_out=16'h82e9;
17'hfb93:	data_out=16'h81b4;
17'hfb94:	data_out=16'h8292;
17'hfb95:	data_out=16'h11c;
17'hfb96:	data_out=16'h29;
17'hfb97:	data_out=16'h834e;
17'hfb98:	data_out=16'h80cc;
17'hfb99:	data_out=16'h208;
17'hfb9a:	data_out=16'h80f3;
17'hfb9b:	data_out=16'h8179;
17'hfb9c:	data_out=16'h54;
17'hfb9d:	data_out=16'h258;
17'hfb9e:	data_out=16'h81ce;
17'hfb9f:	data_out=16'h827e;
17'hfba0:	data_out=16'h175;
17'hfba1:	data_out=16'h80b6;
17'hfba2:	data_out=16'h812b;
17'hfba3:	data_out=16'h22;
17'hfba4:	data_out=16'h17;
17'hfba5:	data_out=16'h80b6;
17'hfba6:	data_out=16'h15e;
17'hfba7:	data_out=16'h22c;
17'hfba8:	data_out=16'h80bd;
17'hfba9:	data_out=16'h81c9;
17'hfbaa:	data_out=16'h8241;
17'hfbab:	data_out=16'h676;
17'hfbac:	data_out=16'h80be;
17'hfbad:	data_out=16'h115;
17'hfbae:	data_out=16'h83a2;
17'hfbaf:	data_out=16'h8069;
17'hfbb0:	data_out=16'h81d9;
17'hfbb1:	data_out=16'h588;
17'hfbb2:	data_out=16'h81bd;
17'hfbb3:	data_out=16'h81fd;
17'hfbb4:	data_out=16'h50f;
17'hfbb5:	data_out=16'h807d;
17'hfbb6:	data_out=16'h8169;
17'hfbb7:	data_out=16'h8376;
17'hfbb8:	data_out=16'h365;
17'hfbb9:	data_out=16'h806e;
17'hfbba:	data_out=16'h80a8;
17'hfbbb:	data_out=16'h26c;
17'hfbbc:	data_out=16'h8272;
17'hfbbd:	data_out=16'h336;
17'hfbbe:	data_out=16'h80c1;
17'hfbbf:	data_out=16'h818e;
17'hfbc0:	data_out=16'h81d4;
17'hfbc1:	data_out=16'h8297;
17'hfbc2:	data_out=16'h80d4;
17'hfbc3:	data_out=16'h82f1;
17'hfbc4:	data_out=16'h14f;
17'hfbc5:	data_out=16'h116;
17'hfbc6:	data_out=16'h8163;
17'hfbc7:	data_out=16'h8125;
17'hfbc8:	data_out=16'h827d;
17'hfbc9:	data_out=16'h80c0;
17'hfbca:	data_out=16'h8219;
17'hfbcb:	data_out=16'h828c;
17'hfbcc:	data_out=16'h820f;
17'hfbcd:	data_out=16'h808c;
17'hfbce:	data_out=16'h8180;
17'hfbcf:	data_out=16'h8181;
17'hfbd0:	data_out=16'h826e;
17'hfbd1:	data_out=16'h81bc;
17'hfbd2:	data_out=16'h26;
17'hfbd3:	data_out=16'h11;
17'hfbd4:	data_out=16'h59;
17'hfbd5:	data_out=16'h8393;
17'hfbd6:	data_out=16'h820d;
17'hfbd7:	data_out=16'h81c4;
17'hfbd8:	data_out=16'h8309;
17'hfbd9:	data_out=16'h8162;
17'hfbda:	data_out=16'h82d8;
17'hfbdb:	data_out=16'h48;
17'hfbdc:	data_out=16'h6d;
17'hfbdd:	data_out=16'h8183;
17'hfbde:	data_out=16'h810f;
17'hfbdf:	data_out=16'h808f;
17'hfbe0:	data_out=16'h14e;
17'hfbe1:	data_out=16'hbd;
17'hfbe2:	data_out=16'h8372;
17'hfbe3:	data_out=16'h8223;
17'hfbe4:	data_out=16'h533;
17'hfbe5:	data_out=16'hdf;
17'hfbe6:	data_out=16'h18d;
17'hfbe7:	data_out=16'h8250;
17'hfbe8:	data_out=16'h80c0;
17'hfbe9:	data_out=16'h8131;
17'hfbea:	data_out=16'h80b8;
17'hfbeb:	data_out=16'he5;
17'hfbec:	data_out=16'h1ca;
17'hfbed:	data_out=16'h81fa;
17'hfbee:	data_out=16'h80bc;
17'hfbef:	data_out=16'h826b;
17'hfbf0:	data_out=16'h80bf;
17'hfbf1:	data_out=16'h835a;
17'hfbf2:	data_out=16'h80df;
17'hfbf3:	data_out=16'h8066;
17'hfbf4:	data_out=16'h81ec;
17'hfbf5:	data_out=16'h82e3;
17'hfbf6:	data_out=16'h381;
17'hfbf7:	data_out=16'h823b;
17'hfbf8:	data_out=16'h8117;
17'hfbf9:	data_out=16'h841b;
17'hfbfa:	data_out=16'h8271;
17'hfbfb:	data_out=16'h80bb;
17'hfbfc:	data_out=16'h8128;
17'hfbfd:	data_out=16'h825c;
17'hfbfe:	data_out=16'h15e;
17'hfbff:	data_out=16'h81d0;
17'hfc00:	data_out=16'h8023;
17'hfc01:	data_out=16'h800c;
17'hfc02:	data_out=16'h49;
17'hfc03:	data_out=16'h8001;
17'hfc04:	data_out=16'h8049;
17'hfc05:	data_out=16'h8039;
17'hfc06:	data_out=16'h802a;
17'hfc07:	data_out=16'h8037;
17'hfc08:	data_out=16'h6;
17'hfc09:	data_out=16'h8019;
17'hfc0a:	data_out=16'h8005;
17'hfc0b:	data_out=16'h8000;
17'hfc0c:	data_out=16'h8039;
17'hfc0d:	data_out=16'h8031;
17'hfc0e:	data_out=16'h8012;
17'hfc0f:	data_out=16'h801a;
17'hfc10:	data_out=16'h36;
17'hfc11:	data_out=16'h8047;
17'hfc12:	data_out=16'h17;
17'hfc13:	data_out=16'h8019;
17'hfc14:	data_out=16'h19;
17'hfc15:	data_out=16'h803a;
17'hfc16:	data_out=16'h8021;
17'hfc17:	data_out=16'h1c;
17'hfc18:	data_out=16'h801f;
17'hfc19:	data_out=16'h8048;
17'hfc1a:	data_out=16'h8067;
17'hfc1b:	data_out=16'h8009;
17'hfc1c:	data_out=16'h8012;
17'hfc1d:	data_out=16'h3a;
17'hfc1e:	data_out=16'ha;
17'hfc1f:	data_out=16'h803f;
17'hfc20:	data_out=16'h800f;
17'hfc21:	data_out=16'h8005;
17'hfc22:	data_out=16'h3b;
17'hfc23:	data_out=16'h803d;
17'hfc24:	data_out=16'h804e;
17'hfc25:	data_out=16'h15;
17'hfc26:	data_out=16'ha;
17'hfc27:	data_out=16'h2b;
17'hfc28:	data_out=16'h800b;
17'hfc29:	data_out=16'h1;
17'hfc2a:	data_out=16'h8;
17'hfc2b:	data_out=16'h8005;
17'hfc2c:	data_out=16'h801d;
17'hfc2d:	data_out=16'h49;
17'hfc2e:	data_out=16'h30;
17'hfc2f:	data_out=16'h1e;
17'hfc30:	data_out=16'h8053;
17'hfc31:	data_out=16'h803b;
17'hfc32:	data_out=16'h8056;
17'hfc33:	data_out=16'h20;
17'hfc34:	data_out=16'h8043;
17'hfc35:	data_out=16'h804c;
17'hfc36:	data_out=16'h18;
17'hfc37:	data_out=16'h31;
17'hfc38:	data_out=16'h8062;
17'hfc39:	data_out=16'h8013;
17'hfc3a:	data_out=16'h37;
17'hfc3b:	data_out=16'h8044;
17'hfc3c:	data_out=16'h69;
17'hfc3d:	data_out=16'h8033;
17'hfc3e:	data_out=16'h800b;
17'hfc3f:	data_out=16'h804b;
17'hfc40:	data_out=16'h8015;
17'hfc41:	data_out=16'h3c;
17'hfc42:	data_out=16'h13;
17'hfc43:	data_out=16'h801c;
17'hfc44:	data_out=16'h801f;
17'hfc45:	data_out=16'h8021;
17'hfc46:	data_out=16'h7d;
17'hfc47:	data_out=16'h801f;
17'hfc48:	data_out=16'h2f;
17'hfc49:	data_out=16'h2a;
17'hfc4a:	data_out=16'h8056;
17'hfc4b:	data_out=16'h8014;
17'hfc4c:	data_out=16'h8013;
17'hfc4d:	data_out=16'h24;
17'hfc4e:	data_out=16'h801d;
17'hfc4f:	data_out=16'h802c;
17'hfc50:	data_out=16'h8022;
17'hfc51:	data_out=16'h8040;
17'hfc52:	data_out=16'h8049;
17'hfc53:	data_out=16'h21;
17'hfc54:	data_out=16'h7;
17'hfc55:	data_out=16'h16;
17'hfc56:	data_out=16'h21;
17'hfc57:	data_out=16'h4b;
17'hfc58:	data_out=16'h63;
17'hfc59:	data_out=16'h2b;
17'hfc5a:	data_out=16'h4a;
17'hfc5b:	data_out=16'h8060;
17'hfc5c:	data_out=16'h8005;
17'hfc5d:	data_out=16'h13;
17'hfc5e:	data_out=16'h8001;
17'hfc5f:	data_out=16'h2;
17'hfc60:	data_out=16'h800b;
17'hfc61:	data_out=16'h8059;
17'hfc62:	data_out=16'h8;
17'hfc63:	data_out=16'h1b;
17'hfc64:	data_out=16'h803d;
17'hfc65:	data_out=16'h8001;
17'hfc66:	data_out=16'h803c;
17'hfc67:	data_out=16'h38;
17'hfc68:	data_out=16'h800e;
17'hfc69:	data_out=16'h1d;
17'hfc6a:	data_out=16'h8011;
17'hfc6b:	data_out=16'h8051;
17'hfc6c:	data_out=16'h5e;
17'hfc6d:	data_out=16'h13;
17'hfc6e:	data_out=16'h8012;
17'hfc6f:	data_out=16'h8002;
17'hfc70:	data_out=16'h8008;
17'hfc71:	data_out=16'h8023;
17'hfc72:	data_out=16'h8012;
17'hfc73:	data_out=16'h8041;
17'hfc74:	data_out=16'h8052;
17'hfc75:	data_out=16'h8036;
17'hfc76:	data_out=16'h8014;
17'hfc77:	data_out=16'h8029;
17'hfc78:	data_out=16'h803c;
17'hfc79:	data_out=16'h18;
17'hfc7a:	data_out=16'h19;
17'hfc7b:	data_out=16'h8011;
17'hfc7c:	data_out=16'h8009;
17'hfc7d:	data_out=16'h8061;
17'hfc7e:	data_out=16'h5;
17'hfc7f:	data_out=16'h8033;
17'hfc80:	data_out=16'h8001;
17'hfc81:	data_out=16'h18;
17'hfc82:	data_out=16'h2a;
17'hfc83:	data_out=16'h2a;
17'hfc84:	data_out=16'h15;
17'hfc85:	data_out=16'h34;
17'hfc86:	data_out=16'h47;
17'hfc87:	data_out=16'h33;
17'hfc88:	data_out=16'h2a;
17'hfc89:	data_out=16'hd;
17'hfc8a:	data_out=16'h24;
17'hfc8b:	data_out=16'h58;
17'hfc8c:	data_out=16'h30;
17'hfc8d:	data_out=16'h1b;
17'hfc8e:	data_out=16'h17;
17'hfc8f:	data_out=16'h28;
17'hfc90:	data_out=16'h19;
17'hfc91:	data_out=16'h1d;
17'hfc92:	data_out=16'h50;
17'hfc93:	data_out=16'h28;
17'hfc94:	data_out=16'h50;
17'hfc95:	data_out=16'hb;
17'hfc96:	data_out=16'h19;
17'hfc97:	data_out=16'h5c;
17'hfc98:	data_out=16'h11;
17'hfc99:	data_out=16'hd;
17'hfc9a:	data_out=16'h1a;
17'hfc9b:	data_out=16'h47;
17'hfc9c:	data_out=16'h40;
17'hfc9d:	data_out=16'h31;
17'hfc9e:	data_out=16'h47;
17'hfc9f:	data_out=16'h3f;
17'hfca0:	data_out=16'h2f;
17'hfca1:	data_out=16'he;
17'hfca2:	data_out=16'h2d;
17'hfca3:	data_out=16'h8011;
17'hfca4:	data_out=16'h8002;
17'hfca5:	data_out=16'h24;
17'hfca6:	data_out=16'h2b;
17'hfca7:	data_out=16'h34;
17'hfca8:	data_out=16'h17;
17'hfca9:	data_out=16'h3a;
17'hfcaa:	data_out=16'h37;
17'hfcab:	data_out=16'h1e;
17'hfcac:	data_out=16'h28;
17'hfcad:	data_out=16'h18;
17'hfcae:	data_out=16'h49;
17'hfcaf:	data_out=16'h35;
17'hfcb0:	data_out=16'h37;
17'hfcb1:	data_out=16'h1b;
17'hfcb2:	data_out=16'h36;
17'hfcb3:	data_out=16'h3c;
17'hfcb4:	data_out=16'h19;
17'hfcb5:	data_out=16'h3d;
17'hfcb6:	data_out=16'h3b;
17'hfcb7:	data_out=16'h3b;
17'hfcb8:	data_out=16'h2e;
17'hfcb9:	data_out=16'h2c;
17'hfcba:	data_out=16'h12;
17'hfcbb:	data_out=16'h1c;
17'hfcbc:	data_out=16'h48;
17'hfcbd:	data_out=16'h6;
17'hfcbe:	data_out=16'h9;
17'hfcbf:	data_out=16'h23;
17'hfcc0:	data_out=16'h12;
17'hfcc1:	data_out=16'h51;
17'hfcc2:	data_out=16'h21;
17'hfcc3:	data_out=16'h2d;
17'hfcc4:	data_out=16'h1d;
17'hfcc5:	data_out=16'h8;
17'hfcc6:	data_out=16'h30;
17'hfcc7:	data_out=16'h19;
17'hfcc8:	data_out=16'h4e;
17'hfcc9:	data_out=16'h27;
17'hfcca:	data_out=16'h37;
17'hfccb:	data_out=16'h4e;
17'hfccc:	data_out=16'h2b;
17'hfccd:	data_out=16'h1a;
17'hfcce:	data_out=16'h28;
17'hfccf:	data_out=16'h31;
17'hfcd0:	data_out=16'hf;
17'hfcd1:	data_out=16'h22;
17'hfcd2:	data_out=16'h8009;
17'hfcd3:	data_out=16'h47;
17'hfcd4:	data_out=16'h31;
17'hfcd5:	data_out=16'h49;
17'hfcd6:	data_out=16'h2c;
17'hfcd7:	data_out=16'h17;
17'hfcd8:	data_out=16'h34;
17'hfcd9:	data_out=16'h14;
17'hfcda:	data_out=16'h4e;
17'hfcdb:	data_out=16'h31;
17'hfcdc:	data_out=16'h2e;
17'hfcdd:	data_out=16'h22;
17'hfcde:	data_out=16'h40;
17'hfcdf:	data_out=16'h1b;
17'hfce0:	data_out=16'h27;
17'hfce1:	data_out=16'h26;
17'hfce2:	data_out=16'h5a;
17'hfce3:	data_out=16'h4d;
17'hfce4:	data_out=16'h1d;
17'hfce5:	data_out=16'h33;
17'hfce6:	data_out=16'h14;
17'hfce7:	data_out=16'h37;
17'hfce8:	data_out=16'h13;
17'hfce9:	data_out=16'h37;
17'hfcea:	data_out=16'h14;
17'hfceb:	data_out=16'h2a;
17'hfcec:	data_out=16'ha;
17'hfced:	data_out=16'h4c;
17'hfcee:	data_out=16'h11;
17'hfcef:	data_out=16'h2c;
17'hfcf0:	data_out=16'hd;
17'hfcf1:	data_out=16'h41;
17'hfcf2:	data_out=16'h2d;
17'hfcf3:	data_out=16'h28;
17'hfcf4:	data_out=16'h2f;
17'hfcf5:	data_out=16'h48;
17'hfcf6:	data_out=16'h22;
17'hfcf7:	data_out=16'h1f;
17'hfcf8:	data_out=16'h24;
17'hfcf9:	data_out=16'h4c;
17'hfcfa:	data_out=16'h57;
17'hfcfb:	data_out=16'hf;
17'hfcfc:	data_out=16'h14;
17'hfcfd:	data_out=16'h3f;
17'hfcfe:	data_out=16'h28;
17'hfcff:	data_out=16'h9;
17'hfd00:	data_out=16'h863a;
17'hfd01:	data_out=16'h27;
17'hfd02:	data_out=16'h357;
17'hfd03:	data_out=16'h3e;
17'hfd04:	data_out=16'h81df;
17'hfd05:	data_out=16'h390;
17'hfd06:	data_out=16'h42c;
17'hfd07:	data_out=16'h207;
17'hfd08:	data_out=16'h1be;
17'hfd09:	data_out=16'h8117;
17'hfd0a:	data_out=16'h8488;
17'hfd0b:	data_out=16'h52f;
17'hfd0c:	data_out=16'h2d5;
17'hfd0d:	data_out=16'h1b7;
17'hfd0e:	data_out=16'h48;
17'hfd0f:	data_out=16'h57f;
17'hfd10:	data_out=16'h81f4;
17'hfd11:	data_out=16'h80c1;
17'hfd12:	data_out=16'h627;
17'hfd13:	data_out=16'h97;
17'hfd14:	data_out=16'h385;
17'hfd15:	data_out=16'h8253;
17'hfd16:	data_out=16'h821c;
17'hfd17:	data_out=16'h459;
17'hfd18:	data_out=16'h8049;
17'hfd19:	data_out=16'h8020;
17'hfd1a:	data_out=16'h8183;
17'hfd1b:	data_out=16'h772;
17'hfd1c:	data_out=16'h29a;
17'hfd1d:	data_out=16'h1b1;
17'hfd1e:	data_out=16'h507;
17'hfd1f:	data_out=16'h38b;
17'hfd20:	data_out=16'h28b;
17'hfd21:	data_out=16'h5a;
17'hfd22:	data_out=16'h80d3;
17'hfd23:	data_out=16'h82ba;
17'hfd24:	data_out=16'h82bb;
17'hfd25:	data_out=16'h8199;
17'hfd26:	data_out=16'h8047;
17'hfd27:	data_out=16'h2f0;
17'hfd28:	data_out=16'ha1;
17'hfd29:	data_out=16'h13c;
17'hfd2a:	data_out=16'h45a;
17'hfd2b:	data_out=16'h40d;
17'hfd2c:	data_out=16'h81e1;
17'hfd2d:	data_out=16'h8538;
17'hfd2e:	data_out=16'h56e;
17'hfd2f:	data_out=16'h41a;
17'hfd30:	data_out=16'h8271;
17'hfd31:	data_out=16'h8028;
17'hfd32:	data_out=16'h8282;
17'hfd33:	data_out=16'h44d;
17'hfd34:	data_out=16'h10f;
17'hfd35:	data_out=16'h1e6;
17'hfd36:	data_out=16'h323;
17'hfd37:	data_out=16'h3a5;
17'hfd38:	data_out=16'h263;
17'hfd39:	data_out=16'h4d7;
17'hfd3a:	data_out=16'h81a3;
17'hfd3b:	data_out=16'h8130;
17'hfd3c:	data_out=16'h1bd;
17'hfd3d:	data_out=16'h82af;
17'hfd3e:	data_out=16'haa;
17'hfd3f:	data_out=16'h37a;
17'hfd40:	data_out=16'h8165;
17'hfd41:	data_out=16'h583;
17'hfd42:	data_out=16'h8374;
17'hfd43:	data_out=16'h31c;
17'hfd44:	data_out=16'h8158;
17'hfd45:	data_out=16'h8256;
17'hfd46:	data_out=16'h139;
17'hfd47:	data_out=16'h8049;
17'hfd48:	data_out=16'h5ca;
17'hfd49:	data_out=16'h81dd;
17'hfd4a:	data_out=16'h27c;
17'hfd4b:	data_out=16'h115;
17'hfd4c:	data_out=16'ha7;
17'hfd4d:	data_out=16'h80f7;
17'hfd4e:	data_out=16'h3fd;
17'hfd4f:	data_out=16'h8035;
17'hfd50:	data_out=16'h813c;
17'hfd51:	data_out=16'h22a;
17'hfd52:	data_out=16'h844d;
17'hfd53:	data_out=16'h5b2;
17'hfd54:	data_out=16'h227;
17'hfd55:	data_out=16'h213;
17'hfd56:	data_out=16'h803d;
17'hfd57:	data_out=16'h80b1;
17'hfd58:	data_out=16'h1cd;
17'hfd59:	data_out=16'h818e;
17'hfd5a:	data_out=16'h45e;
17'hfd5b:	data_out=16'h226;
17'hfd5c:	data_out=16'h3b4;
17'hfd5d:	data_out=16'h806f;
17'hfd5e:	data_out=16'h3ef;
17'hfd5f:	data_out=16'hb6;
17'hfd60:	data_out=16'h81dd;
17'hfd61:	data_out=16'hac;
17'hfd62:	data_out=16'h62e;
17'hfd63:	data_out=16'h488;
17'hfd64:	data_out=16'h1e8;
17'hfd65:	data_out=16'h80b0;
17'hfd66:	data_out=16'h800a;
17'hfd67:	data_out=16'h3c4;
17'hfd68:	data_out=16'h6f;
17'hfd69:	data_out=16'h12c;
17'hfd6a:	data_out=16'h2c;
17'hfd6b:	data_out=16'h7b;
17'hfd6c:	data_out=16'h87b4;
17'hfd6d:	data_out=16'h49a;
17'hfd6e:	data_out=16'h38;
17'hfd6f:	data_out=16'h80ed;
17'hfd70:	data_out=16'h40;
17'hfd71:	data_out=16'h5cf;
17'hfd72:	data_out=16'h8228;
17'hfd73:	data_out=16'h5e;
17'hfd74:	data_out=16'h826e;
17'hfd75:	data_out=16'h340;
17'hfd76:	data_out=16'h2ad;
17'hfd77:	data_out=16'h8122;
17'hfd78:	data_out=16'h2f6;
17'hfd79:	data_out=16'h6be;
17'hfd7a:	data_out=16'h3d5;
17'hfd7b:	data_out=16'hab;
17'hfd7c:	data_out=16'h88;
17'hfd7d:	data_out=16'h569;
17'hfd7e:	data_out=16'h1e;
17'hfd7f:	data_out=16'h828c;
17'hfd80:	data_out=16'h89fa;
17'hfd81:	data_out=16'h81fd;
17'hfd82:	data_out=16'h56a;
17'hfd83:	data_out=16'h856e;
17'hfd84:	data_out=16'h651;
17'hfd85:	data_out=16'h9f7;
17'hfd86:	data_out=16'h87d;
17'hfd87:	data_out=16'h89ff;
17'hfd88:	data_out=16'h8478;
17'hfd89:	data_out=16'h89ff;
17'hfd8a:	data_out=16'h8a00;
17'hfd8b:	data_out=16'h976;
17'hfd8c:	data_out=16'h8a00;
17'hfd8d:	data_out=16'h2ab;
17'hfd8e:	data_out=16'he4;
17'hfd8f:	data_out=16'h8375;
17'hfd90:	data_out=16'h89ea;
17'hfd91:	data_out=16'ha00;
17'hfd92:	data_out=16'h51f;
17'hfd93:	data_out=16'h879c;
17'hfd94:	data_out=16'ha00;
17'hfd95:	data_out=16'h85d5;
17'hfd96:	data_out=16'h8a00;
17'hfd97:	data_out=16'h9ff;
17'hfd98:	data_out=16'h19;
17'hfd99:	data_out=16'ha00;
17'hfd9a:	data_out=16'h948;
17'hfd9b:	data_out=16'ha00;
17'hfd9c:	data_out=16'h9fb;
17'hfd9d:	data_out=16'h989;
17'hfd9e:	data_out=16'h9f2;
17'hfd9f:	data_out=16'ha00;
17'hfda0:	data_out=16'ha00;
17'hfda1:	data_out=16'h146;
17'hfda2:	data_out=16'h89f7;
17'hfda3:	data_out=16'h8a00;
17'hfda4:	data_out=16'h8a00;
17'hfda5:	data_out=16'h8a00;
17'hfda6:	data_out=16'h8a00;
17'hfda7:	data_out=16'ha00;
17'hfda8:	data_out=16'h212;
17'hfda9:	data_out=16'h8a00;
17'hfdaa:	data_out=16'h89fb;
17'hfdab:	data_out=16'ha00;
17'hfdac:	data_out=16'h8a00;
17'hfdad:	data_out=16'h8a00;
17'hfdae:	data_out=16'h84cb;
17'hfdaf:	data_out=16'ha00;
17'hfdb0:	data_out=16'h8a00;
17'hfdb1:	data_out=16'h63a;
17'hfdb2:	data_out=16'h89ff;
17'hfdb3:	data_out=16'ha00;
17'hfdb4:	data_out=16'h86a0;
17'hfdb5:	data_out=16'h9d3;
17'hfdb6:	data_out=16'h1ac;
17'hfdb7:	data_out=16'h67d;
17'hfdb8:	data_out=16'ha00;
17'hfdb9:	data_out=16'ha00;
17'hfdba:	data_out=16'h89fd;
17'hfdbb:	data_out=16'h89c9;
17'hfdbc:	data_out=16'h673;
17'hfdbd:	data_out=16'h6c1;
17'hfdbe:	data_out=16'h217;
17'hfdbf:	data_out=16'h9f7;
17'hfdc0:	data_out=16'h8982;
17'hfdc1:	data_out=16'h9fa;
17'hfdc2:	data_out=16'h8a00;
17'hfdc3:	data_out=16'h9f7;
17'hfdc4:	data_out=16'ha00;
17'hfdc5:	data_out=16'h86b7;
17'hfdc6:	data_out=16'h89a6;
17'hfdc7:	data_out=16'h89fd;
17'hfdc8:	data_out=16'ha00;
17'hfdc9:	data_out=16'h8a00;
17'hfdca:	data_out=16'hf3;
17'hfdcb:	data_out=16'h8a00;
17'hfdcc:	data_out=16'h8a00;
17'hfdcd:	data_out=16'h89f6;
17'hfdce:	data_out=16'h87dc;
17'hfdcf:	data_out=16'h8a00;
17'hfdd0:	data_out=16'h875b;
17'hfdd1:	data_out=16'h9eb;
17'hfdd2:	data_out=16'h8a00;
17'hfdd3:	data_out=16'ha00;
17'hfdd4:	data_out=16'ha00;
17'hfdd5:	data_out=16'h863;
17'hfdd6:	data_out=16'h89fb;
17'hfdd7:	data_out=16'h89f4;
17'hfdd8:	data_out=16'h7cc;
17'hfdd9:	data_out=16'h89e6;
17'hfdda:	data_out=16'ha00;
17'hfddb:	data_out=16'ha00;
17'hfddc:	data_out=16'ha00;
17'hfddd:	data_out=16'h89f5;
17'hfdde:	data_out=16'h9ff;
17'hfddf:	data_out=16'h801d;
17'hfde0:	data_out=16'h8a00;
17'hfde1:	data_out=16'h9f5;
17'hfde2:	data_out=16'h772;
17'hfde3:	data_out=16'ha00;
17'hfde4:	data_out=16'h89d;
17'hfde5:	data_out=16'h79c;
17'hfde6:	data_out=16'ha00;
17'hfde7:	data_out=16'h89dd;
17'hfde8:	data_out=16'h18d;
17'hfde9:	data_out=16'h8917;
17'hfdea:	data_out=16'ha7;
17'hfdeb:	data_out=16'h9fd;
17'hfdec:	data_out=16'h8a00;
17'hfded:	data_out=16'ha00;
17'hfdee:	data_out=16'ha7;
17'hfdef:	data_out=16'h895e;
17'hfdf0:	data_out=16'hca;
17'hfdf1:	data_out=16'h7fb;
17'hfdf2:	data_out=16'h89f3;
17'hfdf3:	data_out=16'h771;
17'hfdf4:	data_out=16'h8a00;
17'hfdf5:	data_out=16'h9f2;
17'hfdf6:	data_out=16'h9ff;
17'hfdf7:	data_out=16'h89fc;
17'hfdf8:	data_out=16'h9fa;
17'hfdf9:	data_out=16'h8956;
17'hfdfa:	data_out=16'ha00;
17'hfdfb:	data_out=16'h218;
17'hfdfc:	data_out=16'h6c6;
17'hfdfd:	data_out=16'ha00;
17'hfdfe:	data_out=16'h89fc;
17'hfdff:	data_out=16'h87ec;
17'hfe00:	data_out=16'h944;
17'hfe01:	data_out=16'h9f8;
17'hfe02:	data_out=16'h49a;
17'hfe03:	data_out=16'h89ff;
17'hfe04:	data_out=16'ha00;
17'hfe05:	data_out=16'h8c8;
17'hfe06:	data_out=16'h678;
17'hfe07:	data_out=16'h89e9;
17'hfe08:	data_out=16'h9fa;
17'hfe09:	data_out=16'h89fd;
17'hfe0a:	data_out=16'h743;
17'hfe0b:	data_out=16'h871;
17'hfe0c:	data_out=16'h8a00;
17'hfe0d:	data_out=16'h8a00;
17'hfe0e:	data_out=16'h106;
17'hfe0f:	data_out=16'h859a;
17'hfe10:	data_out=16'h8397;
17'hfe11:	data_out=16'ha00;
17'hfe12:	data_out=16'h9ef;
17'hfe13:	data_out=16'h843f;
17'hfe14:	data_out=16'h9bd;
17'hfe15:	data_out=16'h9f5;
17'hfe16:	data_out=16'h8a00;
17'hfe17:	data_out=16'h31f;
17'hfe18:	data_out=16'h9fe;
17'hfe19:	data_out=16'ha00;
17'hfe1a:	data_out=16'h9e3;
17'hfe1b:	data_out=16'h9e0;
17'hfe1c:	data_out=16'h826;
17'hfe1d:	data_out=16'h9ff;
17'hfe1e:	data_out=16'h7d8;
17'hfe1f:	data_out=16'h9fd;
17'hfe20:	data_out=16'ha00;
17'hfe21:	data_out=16'h10d;
17'hfe22:	data_out=16'h89fc;
17'hfe23:	data_out=16'h8515;
17'hfe24:	data_out=16'h84e8;
17'hfe25:	data_out=16'h89fc;
17'hfe26:	data_out=16'h8a00;
17'hfe27:	data_out=16'ha00;
17'hfe28:	data_out=16'h1af;
17'hfe29:	data_out=16'h8a00;
17'hfe2a:	data_out=16'h89fb;
17'hfe2b:	data_out=16'ha00;
17'hfe2c:	data_out=16'h89ff;
17'hfe2d:	data_out=16'h89fe;
17'hfe2e:	data_out=16'h8438;
17'hfe2f:	data_out=16'h9eb;
17'hfe30:	data_out=16'h8a00;
17'hfe31:	data_out=16'h9fe;
17'hfe32:	data_out=16'h89fe;
17'hfe33:	data_out=16'h9f7;
17'hfe34:	data_out=16'h817;
17'hfe35:	data_out=16'ha00;
17'hfe36:	data_out=16'h9f2;
17'hfe37:	data_out=16'h4d4;
17'hfe38:	data_out=16'ha00;
17'hfe39:	data_out=16'h9f5;
17'hfe3a:	data_out=16'h89ef;
17'hfe3b:	data_out=16'h9fe;
17'hfe3c:	data_out=16'h2e0;
17'hfe3d:	data_out=16'h9e5;
17'hfe3e:	data_out=16'h1b4;
17'hfe3f:	data_out=16'h8b6;
17'hfe40:	data_out=16'h251;
17'hfe41:	data_out=16'h9d1;
17'hfe42:	data_out=16'h8a00;
17'hfe43:	data_out=16'h86bb;
17'hfe44:	data_out=16'ha00;
17'hfe45:	data_out=16'h8cd;
17'hfe46:	data_out=16'h88ff;
17'hfe47:	data_out=16'h89eb;
17'hfe48:	data_out=16'h913;
17'hfe49:	data_out=16'h89fc;
17'hfe4a:	data_out=16'ha00;
17'hfe4b:	data_out=16'h8a00;
17'hfe4c:	data_out=16'h89fe;
17'hfe4d:	data_out=16'h89fb;
17'hfe4e:	data_out=16'h8165;
17'hfe4f:	data_out=16'h8a00;
17'hfe50:	data_out=16'h89fd;
17'hfe51:	data_out=16'h542;
17'hfe52:	data_out=16'h8a00;
17'hfe53:	data_out=16'ha00;
17'hfe54:	data_out=16'h9f6;
17'hfe55:	data_out=16'h89fd;
17'hfe56:	data_out=16'h3c1;
17'hfe57:	data_out=16'h845a;
17'hfe58:	data_out=16'h9cd;
17'hfe59:	data_out=16'h83c3;
17'hfe5a:	data_out=16'h9fa;
17'hfe5b:	data_out=16'ha00;
17'hfe5c:	data_out=16'h9dd;
17'hfe5d:	data_out=16'h89fa;
17'hfe5e:	data_out=16'h950;
17'hfe5f:	data_out=16'h9fd;
17'hfe60:	data_out=16'h8a00;
17'hfe61:	data_out=16'h8b2;
17'hfe62:	data_out=16'h88c6;
17'hfe63:	data_out=16'h9f8;
17'hfe64:	data_out=16'ha00;
17'hfe65:	data_out=16'ha00;
17'hfe66:	data_out=16'ha00;
17'hfe67:	data_out=16'h89c6;
17'hfe68:	data_out=16'h138;
17'hfe69:	data_out=16'h114;
17'hfe6a:	data_out=16'hf1;
17'hfe6b:	data_out=16'h9e8;
17'hfe6c:	data_out=16'h89f8;
17'hfe6d:	data_out=16'h9f8;
17'hfe6e:	data_out=16'hee;
17'hfe6f:	data_out=16'h8a00;
17'hfe70:	data_out=16'hff;
17'hfe71:	data_out=16'h9cb;
17'hfe72:	data_out=16'h89dc;
17'hfe73:	data_out=16'h1b3;
17'hfe74:	data_out=16'h8a00;
17'hfe75:	data_out=16'h350;
17'hfe76:	data_out=16'h9fa;
17'hfe77:	data_out=16'h89fc;
17'hfe78:	data_out=16'h8a00;
17'hfe79:	data_out=16'h8150;
17'hfe7a:	data_out=16'h9ee;
17'hfe7b:	data_out=16'h1b2;
17'hfe7c:	data_out=16'ha00;
17'hfe7d:	data_out=16'ha00;
17'hfe7e:	data_out=16'h89f3;
17'hfe7f:	data_out=16'h36c;
17'hfe80:	data_out=16'h85af;
17'hfe81:	data_out=16'h992;
17'hfe82:	data_out=16'h611;
17'hfe83:	data_out=16'h8a00;
17'hfe84:	data_out=16'h9ed;
17'hfe85:	data_out=16'h8605;
17'hfe86:	data_out=16'h9fb;
17'hfe87:	data_out=16'h9e0;
17'hfe88:	data_out=16'h9db;
17'hfe89:	data_out=16'h89f5;
17'hfe8a:	data_out=16'ha00;
17'hfe8b:	data_out=16'ha00;
17'hfe8c:	data_out=16'h8797;
17'hfe8d:	data_out=16'h8a00;
17'hfe8e:	data_out=16'h9f9;
17'hfe8f:	data_out=16'h879a;
17'hfe90:	data_out=16'h89fa;
17'hfe91:	data_out=16'ha00;
17'hfe92:	data_out=16'h9a1;
17'hfe93:	data_out=16'h398;
17'hfe94:	data_out=16'h6e0;
17'hfe95:	data_out=16'h53a;
17'hfe96:	data_out=16'h8a00;
17'hfe97:	data_out=16'h8634;
17'hfe98:	data_out=16'h950;
17'hfe99:	data_out=16'h9fd;
17'hfe9a:	data_out=16'h7c3;
17'hfe9b:	data_out=16'h905;
17'hfe9c:	data_out=16'h8891;
17'hfe9d:	data_out=16'ha00;
17'hfe9e:	data_out=16'h45;
17'hfe9f:	data_out=16'ha00;
17'hfea0:	data_out=16'h9d2;
17'hfea1:	data_out=16'h9f8;
17'hfea2:	data_out=16'h89fd;
17'hfea3:	data_out=16'h9fd;
17'hfea4:	data_out=16'h9fe;
17'hfea5:	data_out=16'h8995;
17'hfea6:	data_out=16'h89e5;
17'hfea7:	data_out=16'ha00;
17'hfea8:	data_out=16'h9f7;
17'hfea9:	data_out=16'h8a00;
17'hfeaa:	data_out=16'h89f7;
17'hfeab:	data_out=16'ha00;
17'hfeac:	data_out=16'h89ff;
17'hfead:	data_out=16'h8809;
17'hfeae:	data_out=16'h42c;
17'hfeaf:	data_out=16'h91;
17'hfeb0:	data_out=16'h8a00;
17'hfeb1:	data_out=16'h9ff;
17'hfeb2:	data_out=16'h8a00;
17'hfeb3:	data_out=16'h9e4;
17'hfeb4:	data_out=16'h7be;
17'hfeb5:	data_out=16'ha00;
17'hfeb6:	data_out=16'h9d3;
17'hfeb7:	data_out=16'h9d9;
17'hfeb8:	data_out=16'h9fb;
17'hfeb9:	data_out=16'h9bd;
17'hfeba:	data_out=16'h8370;
17'hfebb:	data_out=16'ha00;
17'hfebc:	data_out=16'h81fa;
17'hfebd:	data_out=16'h618;
17'hfebe:	data_out=16'h9f7;
17'hfebf:	data_out=16'h8654;
17'hfec0:	data_out=16'h8da;
17'hfec1:	data_out=16'h89ff;
17'hfec2:	data_out=16'h8a00;
17'hfec3:	data_out=16'h8a00;
17'hfec4:	data_out=16'ha00;
17'hfec5:	data_out=16'h4b2;
17'hfec6:	data_out=16'h8923;
17'hfec7:	data_out=16'h300;
17'hfec8:	data_out=16'h9ed;
17'hfec9:	data_out=16'h8790;
17'hfeca:	data_out=16'h9fb;
17'hfecb:	data_out=16'h89f8;
17'hfecc:	data_out=16'h89fb;
17'hfecd:	data_out=16'h89fe;
17'hfece:	data_out=16'h9fc;
17'hfecf:	data_out=16'h89fc;
17'hfed0:	data_out=16'h8a00;
17'hfed1:	data_out=16'h87bf;
17'hfed2:	data_out=16'h780;
17'hfed3:	data_out=16'h9fa;
17'hfed4:	data_out=16'h9ca;
17'hfed5:	data_out=16'h89d1;
17'hfed6:	data_out=16'h9da;
17'hfed7:	data_out=16'h9c9;
17'hfed8:	data_out=16'h89ff;
17'hfed9:	data_out=16'h51d;
17'hfeda:	data_out=16'ha00;
17'hfedb:	data_out=16'ha00;
17'hfedc:	data_out=16'h988;
17'hfedd:	data_out=16'h89fb;
17'hfede:	data_out=16'h8698;
17'hfedf:	data_out=16'h851;
17'hfee0:	data_out=16'h89cc;
17'hfee1:	data_out=16'h858;
17'hfee2:	data_out=16'h89ae;
17'hfee3:	data_out=16'h9e8;
17'hfee4:	data_out=16'ha00;
17'hfee5:	data_out=16'ha00;
17'hfee6:	data_out=16'ha00;
17'hfee7:	data_out=16'h89f6;
17'hfee8:	data_out=16'h9f8;
17'hfee9:	data_out=16'h9d9;
17'hfeea:	data_out=16'h9f9;
17'hfeeb:	data_out=16'h2a9;
17'hfeec:	data_out=16'h89f5;
17'hfeed:	data_out=16'h9e7;
17'hfeee:	data_out=16'h9f9;
17'hfeef:	data_out=16'h8a00;
17'hfef0:	data_out=16'h9f9;
17'hfef1:	data_out=16'h9a7;
17'hfef2:	data_out=16'h84b8;
17'hfef3:	data_out=16'h5bc;
17'hfef4:	data_out=16'h8a00;
17'hfef5:	data_out=16'h89dc;
17'hfef6:	data_out=16'h7df;
17'hfef7:	data_out=16'h89fc;
17'hfef8:	data_out=16'h8a00;
17'hfef9:	data_out=16'h89fd;
17'hfefa:	data_out=16'h98e;
17'hfefb:	data_out=16'h9f7;
17'hfefc:	data_out=16'h9fb;
17'hfefd:	data_out=16'h9e3;
17'hfefe:	data_out=16'h9f4;
17'hfeff:	data_out=16'h8a00;
17'hff00:	data_out=16'h89dc;
17'hff01:	data_out=16'h3e4;
17'hff02:	data_out=16'h8031;
17'hff03:	data_out=16'h89f9;
17'hff04:	data_out=16'h9fc;
17'hff05:	data_out=16'h8a00;
17'hff06:	data_out=16'h9f9;
17'hff07:	data_out=16'h9e2;
17'hff08:	data_out=16'h53b;
17'hff09:	data_out=16'h89bf;
17'hff0a:	data_out=16'ha00;
17'hff0b:	data_out=16'ha00;
17'hff0c:	data_out=16'h8910;
17'hff0d:	data_out=16'h8a00;
17'hff0e:	data_out=16'h9f7;
17'hff0f:	data_out=16'h89c9;
17'hff10:	data_out=16'h89fa;
17'hff11:	data_out=16'ha00;
17'hff12:	data_out=16'hfd;
17'hff13:	data_out=16'ha00;
17'hff14:	data_out=16'h89dd;
17'hff15:	data_out=16'h1fb;
17'hff16:	data_out=16'h89fc;
17'hff17:	data_out=16'h89f9;
17'hff18:	data_out=16'h8017;
17'hff19:	data_out=16'h8482;
17'hff1a:	data_out=16'h55e;
17'hff1b:	data_out=16'h89a6;
17'hff1c:	data_out=16'h89fe;
17'hff1d:	data_out=16'ha00;
17'hff1e:	data_out=16'h89f2;
17'hff1f:	data_out=16'ha00;
17'hff20:	data_out=16'h3e3;
17'hff21:	data_out=16'h9f6;
17'hff22:	data_out=16'h89fb;
17'hff23:	data_out=16'ha00;
17'hff24:	data_out=16'ha00;
17'hff25:	data_out=16'h847;
17'hff26:	data_out=16'h80c;
17'hff27:	data_out=16'ha00;
17'hff28:	data_out=16'h9f5;
17'hff29:	data_out=16'h8a00;
17'hff2a:	data_out=16'h89ad;
17'hff2b:	data_out=16'ha00;
17'hff2c:	data_out=16'h89fc;
17'hff2d:	data_out=16'ha00;
17'hff2e:	data_out=16'h8865;
17'hff2f:	data_out=16'h89fa;
17'hff30:	data_out=16'h811b;
17'hff31:	data_out=16'h9ef;
17'hff32:	data_out=16'h956;
17'hff33:	data_out=16'h89e6;
17'hff34:	data_out=16'h1de;
17'hff35:	data_out=16'ha00;
17'hff36:	data_out=16'h898b;
17'hff37:	data_out=16'h9d7;
17'hff38:	data_out=16'h9ca;
17'hff39:	data_out=16'h89f7;
17'hff3a:	data_out=16'h11;
17'hff3b:	data_out=16'ha00;
17'hff3c:	data_out=16'h89dc;
17'hff3d:	data_out=16'h8488;
17'hff3e:	data_out=16'h9f5;
17'hff3f:	data_out=16'h8a00;
17'hff40:	data_out=16'h9b2;
17'hff41:	data_out=16'h89fb;
17'hff42:	data_out=16'h89e9;
17'hff43:	data_out=16'h8a00;
17'hff44:	data_out=16'ha00;
17'hff45:	data_out=16'h14e;
17'hff46:	data_out=16'h86d5;
17'hff47:	data_out=16'h595;
17'hff48:	data_out=16'h80e6;
17'hff49:	data_out=16'h811;
17'hff4a:	data_out=16'h282;
17'hff4b:	data_out=16'h89b4;
17'hff4c:	data_out=16'h85dd;
17'hff4d:	data_out=16'h89fe;
17'hff4e:	data_out=16'h5fc;
17'hff4f:	data_out=16'h219;
17'hff50:	data_out=16'h8a00;
17'hff51:	data_out=16'h89fb;
17'hff52:	data_out=16'h9f1;
17'hff53:	data_out=16'h85b;
17'hff54:	data_out=16'h87f5;
17'hff55:	data_out=16'h89aa;
17'hff56:	data_out=16'h9e9;
17'hff57:	data_out=16'h9b2;
17'hff58:	data_out=16'h89ff;
17'hff59:	data_out=16'h993;
17'hff5a:	data_out=16'h9f4;
17'hff5b:	data_out=16'ha00;
17'hff5c:	data_out=16'h8240;
17'hff5d:	data_out=16'h89f9;
17'hff5e:	data_out=16'h89fa;
17'hff5f:	data_out=16'h89f7;
17'hff60:	data_out=16'h89b6;
17'hff61:	data_out=16'h9a9;
17'hff62:	data_out=16'h894d;
17'hff63:	data_out=16'h89d6;
17'hff64:	data_out=16'ha00;
17'hff65:	data_out=16'h9fe;
17'hff66:	data_out=16'h891c;
17'hff67:	data_out=16'h89fb;
17'hff68:	data_out=16'h9f6;
17'hff69:	data_out=16'h67d;
17'hff6a:	data_out=16'h9f7;
17'hff6b:	data_out=16'h89fb;
17'hff6c:	data_out=16'h89f6;
17'hff6d:	data_out=16'h89da;
17'hff6e:	data_out=16'h9f7;
17'hff6f:	data_out=16'h8a00;
17'hff70:	data_out=16'h9f7;
17'hff71:	data_out=16'h89a0;
17'hff72:	data_out=16'h71;
17'hff73:	data_out=16'h9b2;
17'hff74:	data_out=16'h82ef;
17'hff75:	data_out=16'h8a00;
17'hff76:	data_out=16'h89c5;
17'hff77:	data_out=16'h89f7;
17'hff78:	data_out=16'h8a00;
17'hff79:	data_out=16'h89fa;
17'hff7a:	data_out=16'h89dc;
17'hff7b:	data_out=16'h9f5;
17'hff7c:	data_out=16'h39a;
17'hff7d:	data_out=16'h735;
17'hff7e:	data_out=16'h9fa;
17'hff7f:	data_out=16'h8a00;
17'hff80:	data_out=16'h89fa;
17'hff81:	data_out=16'h8a00;
17'hff82:	data_out=16'h8a00;
17'hff83:	data_out=16'h89f9;
17'hff84:	data_out=16'h9bc;
17'hff85:	data_out=16'h8a00;
17'hff86:	data_out=16'h9fe;
17'hff87:	data_out=16'h8081;
17'hff88:	data_out=16'h8a00;
17'hff89:	data_out=16'h6e3;
17'hff8a:	data_out=16'h9f9;
17'hff8b:	data_out=16'ha00;
17'hff8c:	data_out=16'h8901;
17'hff8d:	data_out=16'h8a00;
17'hff8e:	data_out=16'h5c3;
17'hff8f:	data_out=16'h89fe;
17'hff90:	data_out=16'h89f0;
17'hff91:	data_out=16'ha00;
17'hff92:	data_out=16'h8a00;
17'hff93:	data_out=16'h9f8;
17'hff94:	data_out=16'h89ea;
17'hff95:	data_out=16'h89ff;
17'hff96:	data_out=16'h89ff;
17'hff97:	data_out=16'h89e5;
17'hff98:	data_out=16'h8a00;
17'hff99:	data_out=16'h9a3;
17'hff9a:	data_out=16'h89ff;
17'hff9b:	data_out=16'h89f0;
17'hff9c:	data_out=16'h8a00;
17'hff9d:	data_out=16'h9fc;
17'hff9e:	data_out=16'h89f9;
17'hff9f:	data_out=16'h8995;
17'hffa0:	data_out=16'h89f9;
17'hffa1:	data_out=16'h44e;
17'hffa2:	data_out=16'h85d6;
17'hffa3:	data_out=16'h9f6;
17'hffa4:	data_out=16'h9f7;
17'hffa5:	data_out=16'h9b6;
17'hffa6:	data_out=16'h8024;
17'hffa7:	data_out=16'h8571;
17'hffa8:	data_out=16'h251;
17'hffa9:	data_out=16'h8a00;
17'hffaa:	data_out=16'h89f8;
17'hffab:	data_out=16'h9ff;
17'hffac:	data_out=16'h89fe;
17'hffad:	data_out=16'ha00;
17'hffae:	data_out=16'h8900;
17'hffaf:	data_out=16'h8a00;
17'hffb0:	data_out=16'h6bc;
17'hffb1:	data_out=16'h781;
17'hffb2:	data_out=16'h993;
17'hffb3:	data_out=16'h89f1;
17'hffb4:	data_out=16'h8059;
17'hffb5:	data_out=16'h723;
17'hffb6:	data_out=16'h89fe;
17'hffb7:	data_out=16'h89e2;
17'hffb8:	data_out=16'h889;
17'hffb9:	data_out=16'h89fb;
17'hffba:	data_out=16'h44d;
17'hffbb:	data_out=16'h9f8;
17'hffbc:	data_out=16'h89ff;
17'hffbd:	data_out=16'h89ef;
17'hffbe:	data_out=16'h240;
17'hffbf:	data_out=16'h8a00;
17'hffc0:	data_out=16'h6c7;
17'hffc1:	data_out=16'h8a00;
17'hffc2:	data_out=16'h971;
17'hffc3:	data_out=16'h89fd;
17'hffc4:	data_out=16'h9ec;
17'hffc5:	data_out=16'h89ff;
17'hffc6:	data_out=16'h89ff;
17'hffc7:	data_out=16'h8589;
17'hffc8:	data_out=16'h83fd;
17'hffc9:	data_out=16'h975;
17'hffca:	data_out=16'h89e6;
17'hffcb:	data_out=16'h365;
17'hffcc:	data_out=16'h9d3;
17'hffcd:	data_out=16'h89db;
17'hffce:	data_out=16'h89c1;
17'hffcf:	data_out=16'h9f3;
17'hffd0:	data_out=16'h89fc;
17'hffd1:	data_out=16'h8a00;
17'hffd2:	data_out=16'h9e0;
17'hffd3:	data_out=16'h89e3;
17'hffd4:	data_out=16'h89fb;
17'hffd5:	data_out=16'h89f5;
17'hffd6:	data_out=16'h9db;
17'hffd7:	data_out=16'h2ad;
17'hffd8:	data_out=16'h8a00;
17'hffd9:	data_out=16'h994;
17'hffda:	data_out=16'h89e0;
17'hffdb:	data_out=16'ha00;
17'hffdc:	data_out=16'h8a00;
17'hffdd:	data_out=16'h89fc;
17'hffde:	data_out=16'h89fd;
17'hffdf:	data_out=16'h89fe;
17'hffe0:	data_out=16'h8690;
17'hffe1:	data_out=16'hba;
17'hffe2:	data_out=16'h8922;
17'hffe3:	data_out=16'h89eb;
17'hffe4:	data_out=16'ha00;
17'hffe5:	data_out=16'ha00;
17'hffe6:	data_out=16'h8310;
17'hffe7:	data_out=16'h89f6;
17'hffe8:	data_out=16'h398;
17'hffe9:	data_out=16'h8a00;
17'hffea:	data_out=16'h6a5;
17'hffeb:	data_out=16'h89fe;
17'hffec:	data_out=16'h89fc;
17'hffed:	data_out=16'h89ec;
17'hffee:	data_out=16'h6a1;
17'hffef:	data_out=16'h8669;
17'hfff0:	data_out=16'h626;
17'hfff1:	data_out=16'h89fe;
17'hfff2:	data_out=16'h8146;
17'hfff3:	data_out=16'h663;
17'hfff4:	data_out=16'h716;
17'hfff5:	data_out=16'h8a00;
17'hfff6:	data_out=16'h823b;
17'hfff7:	data_out=16'h89f5;
17'hfff8:	data_out=16'h8a00;
17'hfff9:	data_out=16'h8a00;
17'hfffa:	data_out=16'h89f0;
17'hfffb:	data_out=16'h236;
17'hfffc:	data_out=16'h8a00;
17'hfffd:	data_out=16'h89ff;
17'hfffe:	data_out=16'h9fd;
17'hffff:	data_out=16'h8a00;
17'h10000:	data_out=16'h89fb;
17'h10001:	data_out=16'h8786;
17'h10002:	data_out=16'h8a00;
17'h10003:	data_out=16'h89dd;
17'h10004:	data_out=16'h349;
17'h10005:	data_out=16'h89fb;
17'h10006:	data_out=16'ha00;
17'h10007:	data_out=16'h8a00;
17'h10008:	data_out=16'h8a00;
17'h10009:	data_out=16'h83fb;
17'h1000a:	data_out=16'ha00;
17'h1000b:	data_out=16'h88bf;
17'h1000c:	data_out=16'h89fe;
17'h1000d:	data_out=16'h8a00;
17'h1000e:	data_out=16'h87bc;
17'h1000f:	data_out=16'h8a00;
17'h10010:	data_out=16'h8961;
17'h10011:	data_out=16'ha00;
17'h10012:	data_out=16'h8a00;
17'h10013:	data_out=16'h704;
17'h10014:	data_out=16'h89d2;
17'h10015:	data_out=16'h89fe;
17'h10016:	data_out=16'h89fc;
17'h10017:	data_out=16'h89c7;
17'h10018:	data_out=16'h8a00;
17'h10019:	data_out=16'h9df;
17'h1001a:	data_out=16'h879f;
17'h1001b:	data_out=16'h89e4;
17'h1001c:	data_out=16'h8a00;
17'h1001d:	data_out=16'h9f6;
17'h1001e:	data_out=16'h89f4;
17'h1001f:	data_out=16'h89b9;
17'h10020:	data_out=16'h89f7;
17'h10021:	data_out=16'h8913;
17'h10022:	data_out=16'h9fc;
17'h10023:	data_out=16'h9f9;
17'h10024:	data_out=16'h9fa;
17'h10025:	data_out=16'h9f1;
17'h10026:	data_out=16'h89e4;
17'h10027:	data_out=16'h89e4;
17'h10028:	data_out=16'h898d;
17'h10029:	data_out=16'h8a00;
17'h1002a:	data_out=16'h89fb;
17'h1002b:	data_out=16'h67e;
17'h1002c:	data_out=16'h89fb;
17'h1002d:	data_out=16'ha00;
17'h1002e:	data_out=16'h8872;
17'h1002f:	data_out=16'h89e6;
17'h10030:	data_out=16'h88e;
17'h10031:	data_out=16'h9cf;
17'h10032:	data_out=16'h9da;
17'h10033:	data_out=16'h89e8;
17'h10034:	data_out=16'h9c2;
17'h10035:	data_out=16'h89f3;
17'h10036:	data_out=16'h8a00;
17'h10037:	data_out=16'h89fc;
17'h10038:	data_out=16'h868;
17'h10039:	data_out=16'h89f6;
17'h1003a:	data_out=16'h84d6;
17'h1003b:	data_out=16'h9f1;
17'h1003c:	data_out=16'h89cc;
17'h1003d:	data_out=16'h89f2;
17'h1003e:	data_out=16'h8991;
17'h1003f:	data_out=16'h89fc;
17'h10040:	data_out=16'h6a8;
17'h10041:	data_out=16'h8a00;
17'h10042:	data_out=16'h9c8;
17'h10043:	data_out=16'h89ed;
17'h10044:	data_out=16'h87f9;
17'h10045:	data_out=16'h89fe;
17'h10046:	data_out=16'h89ff;
17'h10047:	data_out=16'h89dd;
17'h10048:	data_out=16'h87cd;
17'h10049:	data_out=16'h9f1;
17'h1004a:	data_out=16'h8a00;
17'h1004b:	data_out=16'h9fe;
17'h1004c:	data_out=16'h9eb;
17'h1004d:	data_out=16'ha00;
17'h1004e:	data_out=16'h8a00;
17'h1004f:	data_out=16'h9fd;
17'h10050:	data_out=16'h89bc;
17'h10051:	data_out=16'h8a00;
17'h10052:	data_out=16'h9ed;
17'h10053:	data_out=16'h89dc;
17'h10054:	data_out=16'h89f4;
17'h10055:	data_out=16'h89e4;
17'h10056:	data_out=16'h89db;
17'h10057:	data_out=16'h89eb;
17'h10058:	data_out=16'h8a00;
17'h10059:	data_out=16'h9e7;
17'h1005a:	data_out=16'h89ed;
17'h1005b:	data_out=16'ha00;
17'h1005c:	data_out=16'h89f0;
17'h1005d:	data_out=16'h89f3;
17'h1005e:	data_out=16'h89df;
17'h1005f:	data_out=16'h89fd;
17'h10060:	data_out=16'h59b;
17'h10061:	data_out=16'h520;
17'h10062:	data_out=16'h8863;
17'h10063:	data_out=16'h89e4;
17'h10064:	data_out=16'h9be;
17'h10065:	data_out=16'ha00;
17'h10066:	data_out=16'h89bf;
17'h10067:	data_out=16'h89b8;
17'h10068:	data_out=16'h8940;
17'h10069:	data_out=16'h8a00;
17'h1006a:	data_out=16'h869b;
17'h1006b:	data_out=16'h89e5;
17'h1006c:	data_out=16'h89fb;
17'h1006d:	data_out=16'h89e5;
17'h1006e:	data_out=16'h869b;
17'h1006f:	data_out=16'h44c;
17'h10070:	data_out=16'h873c;
17'h10071:	data_out=16'h8a00;
17'h10072:	data_out=16'h858;
17'h10073:	data_out=16'h9e6;
17'h10074:	data_out=16'h874;
17'h10075:	data_out=16'h89eb;
17'h10076:	data_out=16'h9fd;
17'h10077:	data_out=16'h89cd;
17'h10078:	data_out=16'h89f5;
17'h10079:	data_out=16'h8a00;
17'h1007a:	data_out=16'h89df;
17'h1007b:	data_out=16'h8992;
17'h1007c:	data_out=16'h8a00;
17'h1007d:	data_out=16'h8a00;
17'h1007e:	data_out=16'h9fe;
17'h1007f:	data_out=16'h89fe;
17'h10080:	data_out=16'h89f7;
17'h10081:	data_out=16'h8861;
17'h10082:	data_out=16'h8a00;
17'h10083:	data_out=16'h8996;
17'h10084:	data_out=16'h5dd;
17'h10085:	data_out=16'h89c1;
17'h10086:	data_out=16'ha00;
17'h10087:	data_out=16'h8a00;
17'h10088:	data_out=16'h8a00;
17'h10089:	data_out=16'ha00;
17'h1008a:	data_out=16'ha00;
17'h1008b:	data_out=16'h852d;
17'h1008c:	data_out=16'h89ff;
17'h1008d:	data_out=16'h8a00;
17'h1008e:	data_out=16'h89f0;
17'h1008f:	data_out=16'h8a00;
17'h10090:	data_out=16'ha00;
17'h10091:	data_out=16'ha00;
17'h10092:	data_out=16'h8a00;
17'h10093:	data_out=16'h3e;
17'h10094:	data_out=16'h89e2;
17'h10095:	data_out=16'h89fd;
17'h10096:	data_out=16'h89f4;
17'h10097:	data_out=16'h89d6;
17'h10098:	data_out=16'h8a00;
17'h10099:	data_out=16'h9fd;
17'h1009a:	data_out=16'h4ea;
17'h1009b:	data_out=16'h8a00;
17'h1009c:	data_out=16'h8a00;
17'h1009d:	data_out=16'ha00;
17'h1009e:	data_out=16'h89f9;
17'h1009f:	data_out=16'h89a8;
17'h100a0:	data_out=16'h89f7;
17'h100a1:	data_out=16'h89f1;
17'h100a2:	data_out=16'ha00;
17'h100a3:	data_out=16'ha00;
17'h100a4:	data_out=16'ha00;
17'h100a5:	data_out=16'ha00;
17'h100a6:	data_out=16'h89dd;
17'h100a7:	data_out=16'h89fb;
17'h100a8:	data_out=16'h89f3;
17'h100a9:	data_out=16'h8a00;
17'h100aa:	data_out=16'h89f2;
17'h100ab:	data_out=16'h86e3;
17'h100ac:	data_out=16'h89ce;
17'h100ad:	data_out=16'ha00;
17'h100ae:	data_out=16'h876e;
17'h100af:	data_out=16'h89e5;
17'h100b0:	data_out=16'h9ec;
17'h100b1:	data_out=16'h9f9;
17'h100b2:	data_out=16'h9fc;
17'h100b3:	data_out=16'h8a00;
17'h100b4:	data_out=16'h9d4;
17'h100b5:	data_out=16'h895d;
17'h100b6:	data_out=16'h8a00;
17'h100b7:	data_out=16'h8a00;
17'h100b8:	data_out=16'h8937;
17'h100b9:	data_out=16'h8a00;
17'h100ba:	data_out=16'ha00;
17'h100bb:	data_out=16'h9db;
17'h100bc:	data_out=16'h89e9;
17'h100bd:	data_out=16'h89c8;
17'h100be:	data_out=16'h89f3;
17'h100bf:	data_out=16'h89c3;
17'h100c0:	data_out=16'ha00;
17'h100c1:	data_out=16'h8a00;
17'h100c2:	data_out=16'ha00;
17'h100c3:	data_out=16'h89d6;
17'h100c4:	data_out=16'h8711;
17'h100c5:	data_out=16'h89fd;
17'h100c6:	data_out=16'h8a00;
17'h100c7:	data_out=16'h88c4;
17'h100c8:	data_out=16'h8153;
17'h100c9:	data_out=16'ha00;
17'h100ca:	data_out=16'h8a00;
17'h100cb:	data_out=16'ha00;
17'h100cc:	data_out=16'ha00;
17'h100cd:	data_out=16'ha00;
17'h100ce:	data_out=16'h8a00;
17'h100cf:	data_out=16'ha00;
17'h100d0:	data_out=16'h8505;
17'h100d1:	data_out=16'h8a00;
17'h100d2:	data_out=16'ha00;
17'h100d3:	data_out=16'h8a00;
17'h100d4:	data_out=16'h89fb;
17'h100d5:	data_out=16'h89fb;
17'h100d6:	data_out=16'h8a00;
17'h100d7:	data_out=16'h89e1;
17'h100d8:	data_out=16'h8a00;
17'h100d9:	data_out=16'ha00;
17'h100da:	data_out=16'h8a00;
17'h100db:	data_out=16'h88f6;
17'h100dc:	data_out=16'h8a00;
17'h100dd:	data_out=16'h887d;
17'h100de:	data_out=16'h88f4;
17'h100df:	data_out=16'h89e7;
17'h100e0:	data_out=16'h9ea;
17'h100e1:	data_out=16'h4ec;
17'h100e2:	data_out=16'h8725;
17'h100e3:	data_out=16'h8a00;
17'h100e4:	data_out=16'h98e;
17'h100e5:	data_out=16'ha00;
17'h100e6:	data_out=16'h8999;
17'h100e7:	data_out=16'h86bf;
17'h100e8:	data_out=16'h89f1;
17'h100e9:	data_out=16'h8a00;
17'h100ea:	data_out=16'h89ef;
17'h100eb:	data_out=16'h88d7;
17'h100ec:	data_out=16'h89b2;
17'h100ed:	data_out=16'h8a00;
17'h100ee:	data_out=16'h89ef;
17'h100ef:	data_out=16'h9f9;
17'h100f0:	data_out=16'h89f0;
17'h100f1:	data_out=16'h8a00;
17'h100f2:	data_out=16'ha00;
17'h100f3:	data_out=16'ha00;
17'h100f4:	data_out=16'h924;
17'h100f5:	data_out=16'h89e0;
17'h100f6:	data_out=16'ha00;
17'h100f7:	data_out=16'h8875;
17'h100f8:	data_out=16'h83a9;
17'h100f9:	data_out=16'h8a00;
17'h100fa:	data_out=16'h89fe;
17'h100fb:	data_out=16'h89f3;
17'h100fc:	data_out=16'h8a00;
17'h100fd:	data_out=16'h8a00;
17'h100fe:	data_out=16'ha00;
17'h100ff:	data_out=16'h89e8;
17'h10100:	data_out=16'h89f9;
17'h10101:	data_out=16'h8966;
17'h10102:	data_out=16'h8a00;
17'h10103:	data_out=16'h89fb;
17'h10104:	data_out=16'h9f9;
17'h10105:	data_out=16'h89e8;
17'h10106:	data_out=16'ha00;
17'h10107:	data_out=16'h8a00;
17'h10108:	data_out=16'h8a00;
17'h10109:	data_out=16'ha00;
17'h1010a:	data_out=16'ha00;
17'h1010b:	data_out=16'h8338;
17'h1010c:	data_out=16'h871d;
17'h1010d:	data_out=16'h8a00;
17'h1010e:	data_out=16'h89ff;
17'h1010f:	data_out=16'h8a00;
17'h10110:	data_out=16'ha00;
17'h10111:	data_out=16'ha00;
17'h10112:	data_out=16'h8a00;
17'h10113:	data_out=16'h89ff;
17'h10114:	data_out=16'h8a00;
17'h10115:	data_out=16'h89ff;
17'h10116:	data_out=16'h89fc;
17'h10117:	data_out=16'h8a00;
17'h10118:	data_out=16'h8a00;
17'h10119:	data_out=16'ha00;
17'h1011a:	data_out=16'h6d3;
17'h1011b:	data_out=16'h8a00;
17'h1011c:	data_out=16'h8a00;
17'h1011d:	data_out=16'ha00;
17'h1011e:	data_out=16'h8a00;
17'h1011f:	data_out=16'h8a00;
17'h10120:	data_out=16'h89f9;
17'h10121:	data_out=16'h89ff;
17'h10122:	data_out=16'ha00;
17'h10123:	data_out=16'ha00;
17'h10124:	data_out=16'ha00;
17'h10125:	data_out=16'ha00;
17'h10126:	data_out=16'h89ff;
17'h10127:	data_out=16'h89fd;
17'h10128:	data_out=16'h8a00;
17'h10129:	data_out=16'h8a00;
17'h1012a:	data_out=16'h8a00;
17'h1012b:	data_out=16'h8801;
17'h1012c:	data_out=16'h89f8;
17'h1012d:	data_out=16'ha00;
17'h1012e:	data_out=16'h8949;
17'h1012f:	data_out=16'h8a00;
17'h10130:	data_out=16'h9a3;
17'h10131:	data_out=16'h9eb;
17'h10132:	data_out=16'ha00;
17'h10133:	data_out=16'h8a00;
17'h10134:	data_out=16'h9c2;
17'h10135:	data_out=16'h89f7;
17'h10136:	data_out=16'h8a00;
17'h10137:	data_out=16'h8a00;
17'h10138:	data_out=16'h89fd;
17'h10139:	data_out=16'h8a00;
17'h1013a:	data_out=16'ha00;
17'h1013b:	data_out=16'h806e;
17'h1013c:	data_out=16'h8a00;
17'h1013d:	data_out=16'h89da;
17'h1013e:	data_out=16'h8a00;
17'h1013f:	data_out=16'h89e9;
17'h10140:	data_out=16'ha00;
17'h10141:	data_out=16'h8a00;
17'h10142:	data_out=16'ha00;
17'h10143:	data_out=16'h89fc;
17'h10144:	data_out=16'h89f7;
17'h10145:	data_out=16'h89ff;
17'h10146:	data_out=16'h8a00;
17'h10147:	data_out=16'h8655;
17'h10148:	data_out=16'h503;
17'h10149:	data_out=16'ha00;
17'h1014a:	data_out=16'h8a00;
17'h1014b:	data_out=16'ha00;
17'h1014c:	data_out=16'ha00;
17'h1014d:	data_out=16'ha00;
17'h1014e:	data_out=16'h8a00;
17'h1014f:	data_out=16'ha00;
17'h10150:	data_out=16'h519;
17'h10151:	data_out=16'h8a00;
17'h10152:	data_out=16'ha00;
17'h10153:	data_out=16'h8a00;
17'h10154:	data_out=16'h89fe;
17'h10155:	data_out=16'h8a00;
17'h10156:	data_out=16'h8a00;
17'h10157:	data_out=16'h8a00;
17'h10158:	data_out=16'h8a00;
17'h10159:	data_out=16'ha00;
17'h1015a:	data_out=16'h8a00;
17'h1015b:	data_out=16'h89f9;
17'h1015c:	data_out=16'h8a00;
17'h1015d:	data_out=16'h8693;
17'h1015e:	data_out=16'h8936;
17'h1015f:	data_out=16'h89ef;
17'h10160:	data_out=16'h9df;
17'h10161:	data_out=16'h8997;
17'h10162:	data_out=16'h8962;
17'h10163:	data_out=16'h8a00;
17'h10164:	data_out=16'h97d;
17'h10165:	data_out=16'ha00;
17'h10166:	data_out=16'h89f8;
17'h10167:	data_out=16'h8518;
17'h10168:	data_out=16'h89ff;
17'h10169:	data_out=16'h8a00;
17'h1016a:	data_out=16'h89ff;
17'h1016b:	data_out=16'h87e9;
17'h1016c:	data_out=16'h89b8;
17'h1016d:	data_out=16'h8a00;
17'h1016e:	data_out=16'h89fe;
17'h1016f:	data_out=16'h9d9;
17'h10170:	data_out=16'h89ff;
17'h10171:	data_out=16'h8a00;
17'h10172:	data_out=16'ha00;
17'h10173:	data_out=16'h9d7;
17'h10174:	data_out=16'h7f8;
17'h10175:	data_out=16'h8a00;
17'h10176:	data_out=16'h9f7;
17'h10177:	data_out=16'h855a;
17'h10178:	data_out=16'h9cf;
17'h10179:	data_out=16'h8a00;
17'h1017a:	data_out=16'h8a00;
17'h1017b:	data_out=16'h8a00;
17'h1017c:	data_out=16'h8a00;
17'h1017d:	data_out=16'h89ff;
17'h1017e:	data_out=16'ha00;
17'h1017f:	data_out=16'h89cb;
17'h10180:	data_out=16'h8a00;
17'h10181:	data_out=16'h8a00;
17'h10182:	data_out=16'h8a00;
17'h10183:	data_out=16'h89fc;
17'h10184:	data_out=16'h9fa;
17'h10185:	data_out=16'h89e8;
17'h10186:	data_out=16'ha00;
17'h10187:	data_out=16'h8a00;
17'h10188:	data_out=16'h8a00;
17'h10189:	data_out=16'ha00;
17'h1018a:	data_out=16'ha00;
17'h1018b:	data_out=16'h89f4;
17'h1018c:	data_out=16'h898d;
17'h1018d:	data_out=16'h8a00;
17'h1018e:	data_out=16'h89ff;
17'h1018f:	data_out=16'h8a00;
17'h10190:	data_out=16'ha00;
17'h10191:	data_out=16'ha00;
17'h10192:	data_out=16'h8a00;
17'h10193:	data_out=16'h8a00;
17'h10194:	data_out=16'h8a00;
17'h10195:	data_out=16'h89ff;
17'h10196:	data_out=16'h89fb;
17'h10197:	data_out=16'h8a00;
17'h10198:	data_out=16'h8a00;
17'h10199:	data_out=16'h5ec;
17'h1019a:	data_out=16'h93c;
17'h1019b:	data_out=16'h8a00;
17'h1019c:	data_out=16'h8a00;
17'h1019d:	data_out=16'h9f8;
17'h1019e:	data_out=16'h8a00;
17'h1019f:	data_out=16'h8a00;
17'h101a0:	data_out=16'h89fa;
17'h101a1:	data_out=16'h89ff;
17'h101a2:	data_out=16'ha00;
17'h101a3:	data_out=16'h8336;
17'h101a4:	data_out=16'h83e2;
17'h101a5:	data_out=16'ha00;
17'h101a6:	data_out=16'h8a00;
17'h101a7:	data_out=16'h8a00;
17'h101a8:	data_out=16'h8a00;
17'h101a9:	data_out=16'h8a00;
17'h101aa:	data_out=16'h8a00;
17'h101ab:	data_out=16'h89ff;
17'h101ac:	data_out=16'h89f7;
17'h101ad:	data_out=16'ha00;
17'h101ae:	data_out=16'h89ba;
17'h101af:	data_out=16'h8a00;
17'h101b0:	data_out=16'h8041;
17'h101b1:	data_out=16'h890d;
17'h101b2:	data_out=16'ha00;
17'h101b3:	data_out=16'h8a00;
17'h101b4:	data_out=16'h957;
17'h101b5:	data_out=16'h8a00;
17'h101b6:	data_out=16'h8a00;
17'h101b7:	data_out=16'h8a00;
17'h101b8:	data_out=16'h875a;
17'h101b9:	data_out=16'h8a00;
17'h101ba:	data_out=16'ha00;
17'h101bb:	data_out=16'h89ee;
17'h101bc:	data_out=16'h8a00;
17'h101bd:	data_out=16'h88a1;
17'h101be:	data_out=16'h8a00;
17'h101bf:	data_out=16'h89e7;
17'h101c0:	data_out=16'ha00;
17'h101c1:	data_out=16'h8a00;
17'h101c2:	data_out=16'ha00;
17'h101c3:	data_out=16'h89fd;
17'h101c4:	data_out=16'h89ff;
17'h101c5:	data_out=16'h89ff;
17'h101c6:	data_out=16'h8a00;
17'h101c7:	data_out=16'h87cc;
17'h101c8:	data_out=16'ha00;
17'h101c9:	data_out=16'ha00;
17'h101ca:	data_out=16'h89fb;
17'h101cb:	data_out=16'ha00;
17'h101cc:	data_out=16'ha00;
17'h101cd:	data_out=16'ha00;
17'h101ce:	data_out=16'h8a00;
17'h101cf:	data_out=16'ha00;
17'h101d0:	data_out=16'ha00;
17'h101d1:	data_out=16'h8a00;
17'h101d2:	data_out=16'ha00;
17'h101d3:	data_out=16'h8a00;
17'h101d4:	data_out=16'h8a00;
17'h101d5:	data_out=16'h8a00;
17'h101d6:	data_out=16'h8a00;
17'h101d7:	data_out=16'h8a00;
17'h101d8:	data_out=16'h8a00;
17'h101d9:	data_out=16'ha00;
17'h101da:	data_out=16'h8a00;
17'h101db:	data_out=16'h89ff;
17'h101dc:	data_out=16'h8a00;
17'h101dd:	data_out=16'h582;
17'h101de:	data_out=16'h8895;
17'h101df:	data_out=16'h8936;
17'h101e0:	data_out=16'h89ff;
17'h101e1:	data_out=16'h8992;
17'h101e2:	data_out=16'h8a00;
17'h101e3:	data_out=16'h8a00;
17'h101e4:	data_out=16'h7c5;
17'h101e5:	data_out=16'ha00;
17'h101e6:	data_out=16'h8a00;
17'h101e7:	data_out=16'h8003;
17'h101e8:	data_out=16'h89ff;
17'h101e9:	data_out=16'h8a00;
17'h101ea:	data_out=16'h89ff;
17'h101eb:	data_out=16'h243;
17'h101ec:	data_out=16'h8271;
17'h101ed:	data_out=16'h8a00;
17'h101ee:	data_out=16'h89ff;
17'h101ef:	data_out=16'h716;
17'h101f0:	data_out=16'h89ff;
17'h101f1:	data_out=16'h8a00;
17'h101f2:	data_out=16'ha00;
17'h101f3:	data_out=16'h9e8;
17'h101f4:	data_out=16'h83f2;
17'h101f5:	data_out=16'h8a00;
17'h101f6:	data_out=16'h89f5;
17'h101f7:	data_out=16'h82a8;
17'h101f8:	data_out=16'h9f8;
17'h101f9:	data_out=16'h8a00;
17'h101fa:	data_out=16'h8a00;
17'h101fb:	data_out=16'h8a00;
17'h101fc:	data_out=16'h8a00;
17'h101fd:	data_out=16'h89fc;
17'h101fe:	data_out=16'ha00;
17'h101ff:	data_out=16'ha00;
17'h10200:	data_out=16'h32;
17'h10201:	data_out=16'h8a00;
17'h10202:	data_out=16'h8a00;
17'h10203:	data_out=16'h89ff;
17'h10204:	data_out=16'h82fa;
17'h10205:	data_out=16'h8a00;
17'h10206:	data_out=16'ha00;
17'h10207:	data_out=16'h8a00;
17'h10208:	data_out=16'h8a00;
17'h10209:	data_out=16'h9fc;
17'h1020a:	data_out=16'ha00;
17'h1020b:	data_out=16'h8a00;
17'h1020c:	data_out=16'h8a00;
17'h1020d:	data_out=16'h8a00;
17'h1020e:	data_out=16'h89f6;
17'h1020f:	data_out=16'h8a00;
17'h10210:	data_out=16'ha00;
17'h10211:	data_out=16'ha00;
17'h10212:	data_out=16'h8a00;
17'h10213:	data_out=16'h8a00;
17'h10214:	data_out=16'h8a00;
17'h10215:	data_out=16'h89ff;
17'h10216:	data_out=16'h89fe;
17'h10217:	data_out=16'h8a00;
17'h10218:	data_out=16'h8a00;
17'h10219:	data_out=16'h8a00;
17'h1021a:	data_out=16'h7cb;
17'h1021b:	data_out=16'h8a00;
17'h1021c:	data_out=16'h8a00;
17'h1021d:	data_out=16'h866a;
17'h1021e:	data_out=16'h8a00;
17'h1021f:	data_out=16'h8a00;
17'h10220:	data_out=16'h28b;
17'h10221:	data_out=16'h89f6;
17'h10222:	data_out=16'ha00;
17'h10223:	data_out=16'h8a00;
17'h10224:	data_out=16'h8a00;
17'h10225:	data_out=16'h9ff;
17'h10226:	data_out=16'h8a00;
17'h10227:	data_out=16'h8a00;
17'h10228:	data_out=16'h89fc;
17'h10229:	data_out=16'h8a00;
17'h1022a:	data_out=16'h8a00;
17'h1022b:	data_out=16'h8a00;
17'h1022c:	data_out=16'h86c9;
17'h1022d:	data_out=16'h9f0;
17'h1022e:	data_out=16'h8a00;
17'h1022f:	data_out=16'h898e;
17'h10230:	data_out=16'h8a00;
17'h10231:	data_out=16'h89ff;
17'h10232:	data_out=16'h83b4;
17'h10233:	data_out=16'h8a00;
17'h10234:	data_out=16'h8a00;
17'h10235:	data_out=16'h8a00;
17'h10236:	data_out=16'h8a00;
17'h10237:	data_out=16'h8a00;
17'h10238:	data_out=16'h9ce;
17'h10239:	data_out=16'h8a00;
17'h1023a:	data_out=16'h9ff;
17'h1023b:	data_out=16'h8a00;
17'h1023c:	data_out=16'h8a00;
17'h1023d:	data_out=16'h866;
17'h1023e:	data_out=16'h89fd;
17'h1023f:	data_out=16'h8a00;
17'h10240:	data_out=16'h863;
17'h10241:	data_out=16'h8a00;
17'h10242:	data_out=16'h9fe;
17'h10243:	data_out=16'h8a00;
17'h10244:	data_out=16'h8a00;
17'h10245:	data_out=16'h89ff;
17'h10246:	data_out=16'h8a00;
17'h10247:	data_out=16'h886e;
17'h10248:	data_out=16'h9fd;
17'h10249:	data_out=16'h9eb;
17'h1024a:	data_out=16'h8a00;
17'h1024b:	data_out=16'ha00;
17'h1024c:	data_out=16'ha00;
17'h1024d:	data_out=16'ha00;
17'h1024e:	data_out=16'h8a00;
17'h1024f:	data_out=16'ha00;
17'h10250:	data_out=16'h9ef;
17'h10251:	data_out=16'h8a00;
17'h10252:	data_out=16'h89bd;
17'h10253:	data_out=16'h8a00;
17'h10254:	data_out=16'h103;
17'h10255:	data_out=16'h8a00;
17'h10256:	data_out=16'h8a00;
17'h10257:	data_out=16'h8a00;
17'h10258:	data_out=16'h8a00;
17'h10259:	data_out=16'ha00;
17'h1025a:	data_out=16'h8a00;
17'h1025b:	data_out=16'h8a00;
17'h1025c:	data_out=16'h8a00;
17'h1025d:	data_out=16'h9fc;
17'h1025e:	data_out=16'h69f;
17'h1025f:	data_out=16'h912;
17'h10260:	data_out=16'h8a00;
17'h10261:	data_out=16'h89bf;
17'h10262:	data_out=16'h8a00;
17'h10263:	data_out=16'h8a00;
17'h10264:	data_out=16'h5ae;
17'h10265:	data_out=16'ha00;
17'h10266:	data_out=16'h8a00;
17'h10267:	data_out=16'h7cd;
17'h10268:	data_out=16'h89f7;
17'h10269:	data_out=16'h8a00;
17'h1026a:	data_out=16'h89f6;
17'h1026b:	data_out=16'h7bc;
17'h1026c:	data_out=16'h945;
17'h1026d:	data_out=16'h8a00;
17'h1026e:	data_out=16'h89f6;
17'h1026f:	data_out=16'h84ed;
17'h10270:	data_out=16'h89f6;
17'h10271:	data_out=16'h8a00;
17'h10272:	data_out=16'ha00;
17'h10273:	data_out=16'h9e4;
17'h10274:	data_out=16'h8a00;
17'h10275:	data_out=16'h8a00;
17'h10276:	data_out=16'h8a00;
17'h10277:	data_out=16'h8844;
17'h10278:	data_out=16'h8046;
17'h10279:	data_out=16'h8a00;
17'h1027a:	data_out=16'h8a00;
17'h1027b:	data_out=16'h89fd;
17'h1027c:	data_out=16'h8a00;
17'h1027d:	data_out=16'h8a00;
17'h1027e:	data_out=16'h9ff;
17'h1027f:	data_out=16'ha00;
17'h10280:	data_out=16'h73a;
17'h10281:	data_out=16'h8a00;
17'h10282:	data_out=16'h8a00;
17'h10283:	data_out=16'h652;
17'h10284:	data_out=16'h89d6;
17'h10285:	data_out=16'h89ff;
17'h10286:	data_out=16'ha00;
17'h10287:	data_out=16'h8a00;
17'h10288:	data_out=16'h8a00;
17'h10289:	data_out=16'h9e1;
17'h1028a:	data_out=16'h2a8;
17'h1028b:	data_out=16'h8a00;
17'h1028c:	data_out=16'h8a00;
17'h1028d:	data_out=16'h8a00;
17'h1028e:	data_out=16'h89f8;
17'h1028f:	data_out=16'h8a00;
17'h10290:	data_out=16'ha00;
17'h10291:	data_out=16'h51a;
17'h10292:	data_out=16'h8a00;
17'h10293:	data_out=16'h719;
17'h10294:	data_out=16'h8a00;
17'h10295:	data_out=16'h6a8;
17'h10296:	data_out=16'h8c6;
17'h10297:	data_out=16'h8a00;
17'h10298:	data_out=16'h8a00;
17'h10299:	data_out=16'h8a00;
17'h1029a:	data_out=16'h880f;
17'h1029b:	data_out=16'h8a00;
17'h1029c:	data_out=16'h8a00;
17'h1029d:	data_out=16'h8a00;
17'h1029e:	data_out=16'h390;
17'h1029f:	data_out=16'h89fb;
17'h102a0:	data_out=16'h6c6;
17'h102a1:	data_out=16'h89f8;
17'h102a2:	data_out=16'ha00;
17'h102a3:	data_out=16'h8a00;
17'h102a4:	data_out=16'h8a00;
17'h102a5:	data_out=16'h9bf;
17'h102a6:	data_out=16'h8a00;
17'h102a7:	data_out=16'h8a00;
17'h102a8:	data_out=16'h89fc;
17'h102a9:	data_out=16'h8a00;
17'h102aa:	data_out=16'h8a00;
17'h102ab:	data_out=16'h8a00;
17'h102ac:	data_out=16'h931;
17'h102ad:	data_out=16'h64f;
17'h102ae:	data_out=16'h8a00;
17'h102af:	data_out=16'h530;
17'h102b0:	data_out=16'h8a00;
17'h102b1:	data_out=16'h8a00;
17'h102b2:	data_out=16'h89fe;
17'h102b3:	data_out=16'h89ba;
17'h102b4:	data_out=16'h8a00;
17'h102b5:	data_out=16'h8a00;
17'h102b6:	data_out=16'h8a00;
17'h102b7:	data_out=16'h8a00;
17'h102b8:	data_out=16'ha00;
17'h102b9:	data_out=16'hde;
17'h102ba:	data_out=16'h9c6;
17'h102bb:	data_out=16'h8a00;
17'h102bc:	data_out=16'h8a00;
17'h102bd:	data_out=16'h93d;
17'h102be:	data_out=16'h89fc;
17'h102bf:	data_out=16'h89fe;
17'h102c0:	data_out=16'h2c6;
17'h102c1:	data_out=16'h8a00;
17'h102c2:	data_out=16'h97d;
17'h102c3:	data_out=16'h8a00;
17'h102c4:	data_out=16'h8a00;
17'h102c5:	data_out=16'h5bc;
17'h102c6:	data_out=16'h8a00;
17'h102c7:	data_out=16'h9ac;
17'h102c8:	data_out=16'h9f8;
17'h102c9:	data_out=16'h509;
17'h102ca:	data_out=16'h8a00;
17'h102cb:	data_out=16'h9e9;
17'h102cc:	data_out=16'ha00;
17'h102cd:	data_out=16'ha00;
17'h102ce:	data_out=16'h64b;
17'h102cf:	data_out=16'ha00;
17'h102d0:	data_out=16'h9ef;
17'h102d1:	data_out=16'h8a00;
17'h102d2:	data_out=16'h8a00;
17'h102d3:	data_out=16'h8a00;
17'h102d4:	data_out=16'h642;
17'h102d5:	data_out=16'h8a00;
17'h102d6:	data_out=16'h8a00;
17'h102d7:	data_out=16'h89f9;
17'h102d8:	data_out=16'h8a00;
17'h102d9:	data_out=16'ha00;
17'h102da:	data_out=16'h8a00;
17'h102db:	data_out=16'h8a00;
17'h102dc:	data_out=16'h8a00;
17'h102dd:	data_out=16'h9e3;
17'h102de:	data_out=16'h827;
17'h102df:	data_out=16'h9f4;
17'h102e0:	data_out=16'h8a00;
17'h102e1:	data_out=16'h8a00;
17'h102e2:	data_out=16'h8a00;
17'h102e3:	data_out=16'h8a00;
17'h102e4:	data_out=16'h4bd;
17'h102e5:	data_out=16'h972;
17'h102e6:	data_out=16'h8a00;
17'h102e7:	data_out=16'h683;
17'h102e8:	data_out=16'h89f6;
17'h102e9:	data_out=16'h8a00;
17'h102ea:	data_out=16'h89f8;
17'h102eb:	data_out=16'h81a;
17'h102ec:	data_out=16'h90f;
17'h102ed:	data_out=16'h8a00;
17'h102ee:	data_out=16'h89f8;
17'h102ef:	data_out=16'h189;
17'h102f0:	data_out=16'h89f8;
17'h102f1:	data_out=16'h8a00;
17'h102f2:	data_out=16'ha00;
17'h102f3:	data_out=16'h74d;
17'h102f4:	data_out=16'h8a00;
17'h102f5:	data_out=16'h8a00;
17'h102f6:	data_out=16'h8a00;
17'h102f7:	data_out=16'h956;
17'h102f8:	data_out=16'h89db;
17'h102f9:	data_out=16'hc0;
17'h102fa:	data_out=16'h8a00;
17'h102fb:	data_out=16'h89fc;
17'h102fc:	data_out=16'h8a00;
17'h102fd:	data_out=16'h89ac;
17'h102fe:	data_out=16'ha00;
17'h102ff:	data_out=16'ha00;
17'h10300:	data_out=16'h1f3;
17'h10301:	data_out=16'h8a00;
17'h10302:	data_out=16'h8a00;
17'h10303:	data_out=16'h8e2;
17'h10304:	data_out=16'h8a00;
17'h10305:	data_out=16'h8a00;
17'h10306:	data_out=16'h9ec;
17'h10307:	data_out=16'h8a00;
17'h10308:	data_out=16'h8a00;
17'h10309:	data_out=16'h9ef;
17'h1030a:	data_out=16'h8a00;
17'h1030b:	data_out=16'h8a00;
17'h1030c:	data_out=16'h8a00;
17'h1030d:	data_out=16'h9be;
17'h1030e:	data_out=16'h89fa;
17'h1030f:	data_out=16'h89f7;
17'h10310:	data_out=16'h9ca;
17'h10311:	data_out=16'h8a00;
17'h10312:	data_out=16'h921;
17'h10313:	data_out=16'h9f9;
17'h10314:	data_out=16'h4eb;
17'h10315:	data_out=16'h949;
17'h10316:	data_out=16'h930;
17'h10317:	data_out=16'h8256;
17'h10318:	data_out=16'h8a00;
17'h10319:	data_out=16'h8a00;
17'h1031a:	data_out=16'h8a00;
17'h1031b:	data_out=16'h8a00;
17'h1031c:	data_out=16'h89ff;
17'h1031d:	data_out=16'h8a00;
17'h1031e:	data_out=16'h948;
17'h1031f:	data_out=16'h575;
17'h10320:	data_out=16'h6b3;
17'h10321:	data_out=16'h89f3;
17'h10322:	data_out=16'h9d0;
17'h10323:	data_out=16'h8a00;
17'h10324:	data_out=16'h8a00;
17'h10325:	data_out=16'h56f;
17'h10326:	data_out=16'h8a00;
17'h10327:	data_out=16'h8a00;
17'h10328:	data_out=16'h89ef;
17'h10329:	data_out=16'h8a00;
17'h1032a:	data_out=16'h8a00;
17'h1032b:	data_out=16'h8a00;
17'h1032c:	data_out=16'h98b;
17'h1032d:	data_out=16'h89ff;
17'h1032e:	data_out=16'h89fc;
17'h1032f:	data_out=16'h6f3;
17'h10330:	data_out=16'h89f3;
17'h10331:	data_out=16'h8a00;
17'h10332:	data_out=16'h8a00;
17'h10333:	data_out=16'h9b4;
17'h10334:	data_out=16'h8a00;
17'h10335:	data_out=16'h8a00;
17'h10336:	data_out=16'h8a00;
17'h10337:	data_out=16'h8a00;
17'h10338:	data_out=16'ha00;
17'h10339:	data_out=16'h9d5;
17'h1033a:	data_out=16'h9fa;
17'h1033b:	data_out=16'h8a00;
17'h1033c:	data_out=16'h8a00;
17'h1033d:	data_out=16'h8fa;
17'h1033e:	data_out=16'h89f0;
17'h1033f:	data_out=16'h8a00;
17'h10340:	data_out=16'h8502;
17'h10341:	data_out=16'h8a00;
17'h10342:	data_out=16'h82e0;
17'h10343:	data_out=16'h8a00;
17'h10344:	data_out=16'h8a00;
17'h10345:	data_out=16'h956;
17'h10346:	data_out=16'h8a00;
17'h10347:	data_out=16'h9ff;
17'h10348:	data_out=16'h9f9;
17'h10349:	data_out=16'h83c5;
17'h1034a:	data_out=16'h8a00;
17'h1034b:	data_out=16'h966;
17'h1034c:	data_out=16'h9d6;
17'h1034d:	data_out=16'h9ca;
17'h1034e:	data_out=16'h85f;
17'h1034f:	data_out=16'h532;
17'h10350:	data_out=16'h9d1;
17'h10351:	data_out=16'h89f1;
17'h10352:	data_out=16'h8a00;
17'h10353:	data_out=16'h8a00;
17'h10354:	data_out=16'h67d;
17'h10355:	data_out=16'h89f8;
17'h10356:	data_out=16'h8a00;
17'h10357:	data_out=16'h89f6;
17'h10358:	data_out=16'h8a00;
17'h10359:	data_out=16'h562;
17'h1035a:	data_out=16'h8a00;
17'h1035b:	data_out=16'h8a00;
17'h1035c:	data_out=16'h8a00;
17'h1035d:	data_out=16'h94b;
17'h1035e:	data_out=16'h9d5;
17'h1035f:	data_out=16'h9f4;
17'h10360:	data_out=16'h8a00;
17'h10361:	data_out=16'h8a00;
17'h10362:	data_out=16'h8a00;
17'h10363:	data_out=16'h8c8;
17'h10364:	data_out=16'h48d;
17'h10365:	data_out=16'h849f;
17'h10366:	data_out=16'h8a00;
17'h10367:	data_out=16'h8a00;
17'h10368:	data_out=16'h89e4;
17'h10369:	data_out=16'h8a00;
17'h1036a:	data_out=16'h89fb;
17'h1036b:	data_out=16'h731;
17'h1036c:	data_out=16'h513;
17'h1036d:	data_out=16'h915;
17'h1036e:	data_out=16'h89fb;
17'h1036f:	data_out=16'h8a00;
17'h10370:	data_out=16'h89fb;
17'h10371:	data_out=16'h89fb;
17'h10372:	data_out=16'h997;
17'h10373:	data_out=16'h8a00;
17'h10374:	data_out=16'h89f9;
17'h10375:	data_out=16'h8a00;
17'h10376:	data_out=16'h8a00;
17'h10377:	data_out=16'h9ce;
17'h10378:	data_out=16'h89f9;
17'h10379:	data_out=16'h369;
17'h1037a:	data_out=16'h44d;
17'h1037b:	data_out=16'h89f1;
17'h1037c:	data_out=16'h879d;
17'h1037d:	data_out=16'h9a8;
17'h1037e:	data_out=16'h9f4;
17'h1037f:	data_out=16'ha00;
17'h10380:	data_out=16'h89ff;
17'h10381:	data_out=16'h8a00;
17'h10382:	data_out=16'h8a00;
17'h10383:	data_out=16'h8821;
17'h10384:	data_out=16'h89f9;
17'h10385:	data_out=16'h8a00;
17'h10386:	data_out=16'h9da;
17'h10387:	data_out=16'h852f;
17'h10388:	data_out=16'h8a00;
17'h10389:	data_out=16'h9ce;
17'h1038a:	data_out=16'h8a00;
17'h1038b:	data_out=16'h89fb;
17'h1038c:	data_out=16'h89ff;
17'h1038d:	data_out=16'h73f;
17'h1038e:	data_out=16'h16c;
17'h1038f:	data_out=16'h89f2;
17'h10390:	data_out=16'h97b;
17'h10391:	data_out=16'h8a00;
17'h10392:	data_out=16'h949;
17'h10393:	data_out=16'h9f8;
17'h10394:	data_out=16'h3e;
17'h10395:	data_out=16'h8638;
17'h10396:	data_out=16'h89f9;
17'h10397:	data_out=16'h88f1;
17'h10398:	data_out=16'h9b5;
17'h10399:	data_out=16'h89fc;
17'h1039a:	data_out=16'h8a00;
17'h1039b:	data_out=16'h8a00;
17'h1039c:	data_out=16'h89fd;
17'h1039d:	data_out=16'h8a00;
17'h1039e:	data_out=16'h8cf;
17'h1039f:	data_out=16'h36a;
17'h103a0:	data_out=16'h6fd;
17'h103a1:	data_out=16'h39d;
17'h103a2:	data_out=16'h2b6;
17'h103a3:	data_out=16'h8a00;
17'h103a4:	data_out=16'h8a00;
17'h103a5:	data_out=16'h1ab;
17'h103a6:	data_out=16'h8a00;
17'h103a7:	data_out=16'h8a00;
17'h103a8:	data_out=16'h616;
17'h103a9:	data_out=16'h8a00;
17'h103aa:	data_out=16'h8a00;
17'h103ab:	data_out=16'h8a00;
17'h103ac:	data_out=16'h89d8;
17'h103ad:	data_out=16'h89f9;
17'h103ae:	data_out=16'h89ff;
17'h103af:	data_out=16'h88a;
17'h103b0:	data_out=16'h9b2;
17'h103b1:	data_out=16'h8a00;
17'h103b2:	data_out=16'h8a00;
17'h103b3:	data_out=16'h9e3;
17'h103b4:	data_out=16'h8a00;
17'h103b5:	data_out=16'h8a00;
17'h103b6:	data_out=16'h8a00;
17'h103b7:	data_out=16'h8a00;
17'h103b8:	data_out=16'h9fa;
17'h103b9:	data_out=16'h9f0;
17'h103ba:	data_out=16'h9e8;
17'h103bb:	data_out=16'h8a00;
17'h103bc:	data_out=16'h8a00;
17'h103bd:	data_out=16'h741;
17'h103be:	data_out=16'h61e;
17'h103bf:	data_out=16'h8a00;
17'h103c0:	data_out=16'h307;
17'h103c1:	data_out=16'h89b8;
17'h103c2:	data_out=16'h89fd;
17'h103c3:	data_out=16'h89f4;
17'h103c4:	data_out=16'h8a00;
17'h103c5:	data_out=16'h85e6;
17'h103c6:	data_out=16'h8a00;
17'h103c7:	data_out=16'h9ee;
17'h103c8:	data_out=16'h9d8;
17'h103c9:	data_out=16'h81c3;
17'h103ca:	data_out=16'h9bb;
17'h103cb:	data_out=16'h31a;
17'h103cc:	data_out=16'h39f;
17'h103cd:	data_out=16'h5c4;
17'h103ce:	data_out=16'h81ea;
17'h103cf:	data_out=16'h254;
17'h103d0:	data_out=16'h9af;
17'h103d1:	data_out=16'h89b7;
17'h103d2:	data_out=16'h8a00;
17'h103d3:	data_out=16'h8a00;
17'h103d4:	data_out=16'h58a;
17'h103d5:	data_out=16'h89d8;
17'h103d6:	data_out=16'h8a00;
17'h103d7:	data_out=16'h89f2;
17'h103d8:	data_out=16'h89fd;
17'h103d9:	data_out=16'h18d;
17'h103da:	data_out=16'h89bd;
17'h103db:	data_out=16'h8a00;
17'h103dc:	data_out=16'h8a00;
17'h103dd:	data_out=16'h4f7;
17'h103de:	data_out=16'ha00;
17'h103df:	data_out=16'h9d6;
17'h103e0:	data_out=16'h8a00;
17'h103e1:	data_out=16'h8a00;
17'h103e2:	data_out=16'h8a00;
17'h103e3:	data_out=16'h948;
17'h103e4:	data_out=16'h453;
17'h103e5:	data_out=16'h8358;
17'h103e6:	data_out=16'h9f9;
17'h103e7:	data_out=16'h8a00;
17'h103e8:	data_out=16'h4f1;
17'h103e9:	data_out=16'h884d;
17'h103ea:	data_out=16'h801f;
17'h103eb:	data_out=16'h85d;
17'h103ec:	data_out=16'h8a00;
17'h103ed:	data_out=16'h95d;
17'h103ee:	data_out=16'h8019;
17'h103ef:	data_out=16'h8a00;
17'h103f0:	data_out=16'hb4;
17'h103f1:	data_out=16'h8220;
17'h103f2:	data_out=16'h2e1;
17'h103f3:	data_out=16'h8a00;
17'h103f4:	data_out=16'h87c;
17'h103f5:	data_out=16'h8a00;
17'h103f6:	data_out=16'h8a00;
17'h103f7:	data_out=16'h8a0;
17'h103f8:	data_out=16'h8a00;
17'h103f9:	data_out=16'h848b;
17'h103fa:	data_out=16'h2fb;
17'h103fb:	data_out=16'h61f;
17'h103fc:	data_out=16'h9bc;
17'h103fd:	data_out=16'h9f1;
17'h103fe:	data_out=16'h9e1;
17'h103ff:	data_out=16'h9be;
17'h10400:	data_out=16'h89d7;
17'h10401:	data_out=16'h8a00;
17'h10402:	data_out=16'h8a00;
17'h10403:	data_out=16'h89b4;
17'h10404:	data_out=16'h79f;
17'h10405:	data_out=16'h84fb;
17'h10406:	data_out=16'h9a4;
17'h10407:	data_out=16'h9f0;
17'h10408:	data_out=16'h792;
17'h10409:	data_out=16'hdf;
17'h1040a:	data_out=16'h89ff;
17'h1040b:	data_out=16'h89d8;
17'h1040c:	data_out=16'h6d4;
17'h1040d:	data_out=16'h89c3;
17'h1040e:	data_out=16'h92b;
17'h1040f:	data_out=16'h8a00;
17'h10410:	data_out=16'h64c;
17'h10411:	data_out=16'h8a00;
17'h10412:	data_out=16'h1b4;
17'h10413:	data_out=16'h9eb;
17'h10414:	data_out=16'h89de;
17'h10415:	data_out=16'h89d7;
17'h10416:	data_out=16'h89b8;
17'h10417:	data_out=16'h89ed;
17'h10418:	data_out=16'h9c2;
17'h10419:	data_out=16'ha00;
17'h1041a:	data_out=16'hb8;
17'h1041b:	data_out=16'h89fd;
17'h1041c:	data_out=16'h89f7;
17'h1041d:	data_out=16'h89fd;
17'h1041e:	data_out=16'h89d6;
17'h1041f:	data_out=16'h8886;
17'h10420:	data_out=16'h893;
17'h10421:	data_out=16'h964;
17'h10422:	data_out=16'h8a00;
17'h10423:	data_out=16'h89ea;
17'h10424:	data_out=16'h89ea;
17'h10425:	data_out=16'h8241;
17'h10426:	data_out=16'h8a00;
17'h10427:	data_out=16'h1cc;
17'h10428:	data_out=16'h9b2;
17'h10429:	data_out=16'h8a00;
17'h1042a:	data_out=16'h8a00;
17'h1042b:	data_out=16'h89c7;
17'h1042c:	data_out=16'h89a4;
17'h1042d:	data_out=16'h89fb;
17'h1042e:	data_out=16'h8a00;
17'h1042f:	data_out=16'h7f6;
17'h10430:	data_out=16'ha00;
17'h10431:	data_out=16'h8997;
17'h10432:	data_out=16'h83ac;
17'h10433:	data_out=16'h5fb;
17'h10434:	data_out=16'h89fe;
17'h10435:	data_out=16'h3c0;
17'h10436:	data_out=16'h286;
17'h10437:	data_out=16'h8a00;
17'h10438:	data_out=16'h38f;
17'h10439:	data_out=16'h809e;
17'h1043a:	data_out=16'h904;
17'h1043b:	data_out=16'h9e5;
17'h1043c:	data_out=16'h8a00;
17'h1043d:	data_out=16'h281;
17'h1043e:	data_out=16'h9b3;
17'h1043f:	data_out=16'h8572;
17'h10440:	data_out=16'h42e;
17'h10441:	data_out=16'h5f8;
17'h10442:	data_out=16'h89fd;
17'h10443:	data_out=16'h840b;
17'h10444:	data_out=16'h810d;
17'h10445:	data_out=16'h89d7;
17'h10446:	data_out=16'h8a00;
17'h10447:	data_out=16'h5cc;
17'h10448:	data_out=16'h8c7;
17'h10449:	data_out=16'h263;
17'h1044a:	data_out=16'h9ef;
17'h1044b:	data_out=16'h89fb;
17'h1044c:	data_out=16'h89ff;
17'h1044d:	data_out=16'h8a00;
17'h1044e:	data_out=16'h2e3;
17'h1044f:	data_out=16'h81e2;
17'h10450:	data_out=16'h184;
17'h10451:	data_out=16'h89fd;
17'h10452:	data_out=16'h89fa;
17'h10453:	data_out=16'h83d6;
17'h10454:	data_out=16'ha2;
17'h10455:	data_out=16'h89ff;
17'h10456:	data_out=16'h89fe;
17'h10457:	data_out=16'h8a00;
17'h10458:	data_out=16'h89fe;
17'h10459:	data_out=16'h81d0;
17'h1045a:	data_out=16'h8997;
17'h1045b:	data_out=16'h8a00;
17'h1045c:	data_out=16'h8a00;
17'h1045d:	data_out=16'h896e;
17'h1045e:	data_out=16'ha00;
17'h1045f:	data_out=16'h85f2;
17'h10460:	data_out=16'h8a00;
17'h10461:	data_out=16'h8a00;
17'h10462:	data_out=16'h89ff;
17'h10463:	data_out=16'h357;
17'h10464:	data_out=16'h8047;
17'h10465:	data_out=16'hee;
17'h10466:	data_out=16'ha00;
17'h10467:	data_out=16'h8a00;
17'h10468:	data_out=16'h992;
17'h10469:	data_out=16'h1de;
17'h1046a:	data_out=16'h8f5;
17'h1046b:	data_out=16'h992;
17'h1046c:	data_out=16'h89ff;
17'h1046d:	data_out=16'h3d1;
17'h1046e:	data_out=16'h8f7;
17'h1046f:	data_out=16'h37e;
17'h10470:	data_out=16'h917;
17'h10471:	data_out=16'h89f9;
17'h10472:	data_out=16'h86b8;
17'h10473:	data_out=16'h8a00;
17'h10474:	data_out=16'ha00;
17'h10475:	data_out=16'h8a00;
17'h10476:	data_out=16'h8a00;
17'h10477:	data_out=16'h1ab;
17'h10478:	data_out=16'h8a00;
17'h10479:	data_out=16'h8800;
17'h1047a:	data_out=16'h8464;
17'h1047b:	data_out=16'h9b3;
17'h1047c:	data_out=16'h9da;
17'h1047d:	data_out=16'h9d0;
17'h1047e:	data_out=16'h9b9;
17'h1047f:	data_out=16'h197;
17'h10480:	data_out=16'h897b;
17'h10481:	data_out=16'h89e6;
17'h10482:	data_out=16'h89f2;
17'h10483:	data_out=16'h8986;
17'h10484:	data_out=16'h9eb;
17'h10485:	data_out=16'h89c2;
17'h10486:	data_out=16'h2d8;
17'h10487:	data_out=16'ha00;
17'h10488:	data_out=16'h9fc;
17'h10489:	data_out=16'h743;
17'h1048a:	data_out=16'h89ee;
17'h1048b:	data_out=16'h9f0;
17'h1048c:	data_out=16'h9cf;
17'h1048d:	data_out=16'h89ff;
17'h1048e:	data_out=16'h9ac;
17'h1048f:	data_out=16'h8721;
17'h10490:	data_out=16'h980;
17'h10491:	data_out=16'h89c8;
17'h10492:	data_out=16'h89f9;
17'h10493:	data_out=16'h9f6;
17'h10494:	data_out=16'h82fa;
17'h10495:	data_out=16'h8872;
17'h10496:	data_out=16'h89ad;
17'h10497:	data_out=16'h896e;
17'h10498:	data_out=16'h2f2;
17'h10499:	data_out=16'ha00;
17'h1049a:	data_out=16'h413;
17'h1049b:	data_out=16'h9d8;
17'h1049c:	data_out=16'h89fc;
17'h1049d:	data_out=16'h86e6;
17'h1049e:	data_out=16'h85d2;
17'h1049f:	data_out=16'h89d7;
17'h104a0:	data_out=16'h92c;
17'h104a1:	data_out=16'h9ca;
17'h104a2:	data_out=16'h8a00;
17'h104a3:	data_out=16'h9f4;
17'h104a4:	data_out=16'h9f4;
17'h104a5:	data_out=16'h556;
17'h104a6:	data_out=16'h89d4;
17'h104a7:	data_out=16'h9f3;
17'h104a8:	data_out=16'h9ed;
17'h104a9:	data_out=16'h8a00;
17'h104aa:	data_out=16'h88b2;
17'h104ab:	data_out=16'h9dc;
17'h104ac:	data_out=16'h89af;
17'h104ad:	data_out=16'h795;
17'h104ae:	data_out=16'h89e7;
17'h104af:	data_out=16'h9e4;
17'h104b0:	data_out=16'ha00;
17'h104b1:	data_out=16'h888c;
17'h104b2:	data_out=16'h78f;
17'h104b3:	data_out=16'h277;
17'h104b4:	data_out=16'h89a3;
17'h104b5:	data_out=16'h9e4;
17'h104b6:	data_out=16'h9f2;
17'h104b7:	data_out=16'h89f7;
17'h104b8:	data_out=16'h89b8;
17'h104b9:	data_out=16'h87c1;
17'h104ba:	data_out=16'h9d3;
17'h104bb:	data_out=16'ha00;
17'h104bc:	data_out=16'h8a00;
17'h104bd:	data_out=16'h82e1;
17'h104be:	data_out=16'h9ed;
17'h104bf:	data_out=16'h89c3;
17'h104c0:	data_out=16'h9e6;
17'h104c1:	data_out=16'h7dd;
17'h104c2:	data_out=16'h89d4;
17'h104c3:	data_out=16'h997;
17'h104c4:	data_out=16'h9c8;
17'h104c5:	data_out=16'h8873;
17'h104c6:	data_out=16'h89c7;
17'h104c7:	data_out=16'h2cd;
17'h104c8:	data_out=16'h50;
17'h104c9:	data_out=16'h7b5;
17'h104ca:	data_out=16'ha00;
17'h104cb:	data_out=16'h89c6;
17'h104cc:	data_out=16'h89fe;
17'h104cd:	data_out=16'h89d4;
17'h104ce:	data_out=16'h9ff;
17'h104cf:	data_out=16'h835f;
17'h104d0:	data_out=16'h2c2;
17'h104d1:	data_out=16'h8a00;
17'h104d2:	data_out=16'h9df;
17'h104d3:	data_out=16'h9c1;
17'h104d4:	data_out=16'h662;
17'h104d5:	data_out=16'h8233;
17'h104d6:	data_out=16'h8446;
17'h104d7:	data_out=16'h89fe;
17'h104d8:	data_out=16'h2e2;
17'h104d9:	data_out=16'h561;
17'h104da:	data_out=16'h8990;
17'h104db:	data_out=16'h8a1;
17'h104dc:	data_out=16'h8a00;
17'h104dd:	data_out=16'h8169;
17'h104de:	data_out=16'ha00;
17'h104df:	data_out=16'h8994;
17'h104e0:	data_out=16'h89e0;
17'h104e1:	data_out=16'h89f9;
17'h104e2:	data_out=16'h8898;
17'h104e3:	data_out=16'h6f8;
17'h104e4:	data_out=16'h8982;
17'h104e5:	data_out=16'h8c7;
17'h104e6:	data_out=16'ha00;
17'h104e7:	data_out=16'h89df;
17'h104e8:	data_out=16'h9ed;
17'h104e9:	data_out=16'h308;
17'h104ea:	data_out=16'h990;
17'h104eb:	data_out=16'h716;
17'h104ec:	data_out=16'h8988;
17'h104ed:	data_out=16'h703;
17'h104ee:	data_out=16'h990;
17'h104ef:	data_out=16'h642;
17'h104f0:	data_out=16'h9a1;
17'h104f1:	data_out=16'h89aa;
17'h104f2:	data_out=16'h8963;
17'h104f3:	data_out=16'h89fd;
17'h104f4:	data_out=16'ha00;
17'h104f5:	data_out=16'h8a00;
17'h104f6:	data_out=16'h89fb;
17'h104f7:	data_out=16'h985;
17'h104f8:	data_out=16'h8a00;
17'h104f9:	data_out=16'h9e9;
17'h104fa:	data_out=16'h869;
17'h104fb:	data_out=16'h9ed;
17'h104fc:	data_out=16'h80c0;
17'h104fd:	data_out=16'h9cf;
17'h104fe:	data_out=16'h9ee;
17'h104ff:	data_out=16'h89ec;
17'h10500:	data_out=16'h89fc;
17'h10501:	data_out=16'h89fc;
17'h10502:	data_out=16'h8244;
17'h10503:	data_out=16'h855b;
17'h10504:	data_out=16'h9fc;
17'h10505:	data_out=16'h58f;
17'h10506:	data_out=16'h89c5;
17'h10507:	data_out=16'ha00;
17'h10508:	data_out=16'h8892;
17'h10509:	data_out=16'h9f7;
17'h1050a:	data_out=16'h89fb;
17'h1050b:	data_out=16'h9ff;
17'h1050c:	data_out=16'h9c9;
17'h1050d:	data_out=16'h89f0;
17'h1050e:	data_out=16'h9e2;
17'h1050f:	data_out=16'h326;
17'h10510:	data_out=16'h9f9;
17'h10511:	data_out=16'h89fa;
17'h10512:	data_out=16'h8a00;
17'h10513:	data_out=16'h9f3;
17'h10514:	data_out=16'h82d1;
17'h10515:	data_out=16'h89c8;
17'h10516:	data_out=16'h884e;
17'h10517:	data_out=16'h82e4;
17'h10518:	data_out=16'h8a00;
17'h10519:	data_out=16'ha00;
17'h1051a:	data_out=16'h9be;
17'h1051b:	data_out=16'h9fa;
17'h1051c:	data_out=16'h89ec;
17'h1051d:	data_out=16'h89c7;
17'h1051e:	data_out=16'h85b7;
17'h1051f:	data_out=16'h403;
17'h10520:	data_out=16'h8402;
17'h10521:	data_out=16'h9eb;
17'h10522:	data_out=16'h85de;
17'h10523:	data_out=16'h9f9;
17'h10524:	data_out=16'h9fa;
17'h10525:	data_out=16'h685;
17'h10526:	data_out=16'h8963;
17'h10527:	data_out=16'h973;
17'h10528:	data_out=16'h9ee;
17'h10529:	data_out=16'h89f1;
17'h1052a:	data_out=16'h80d1;
17'h1052b:	data_out=16'h9fe;
17'h1052c:	data_out=16'h89b2;
17'h1052d:	data_out=16'h8475;
17'h1052e:	data_out=16'h8312;
17'h1052f:	data_out=16'h9ec;
17'h10530:	data_out=16'ha00;
17'h10531:	data_out=16'h89be;
17'h10532:	data_out=16'h9fe;
17'h10533:	data_out=16'h894d;
17'h10534:	data_out=16'h89e4;
17'h10535:	data_out=16'h989;
17'h10536:	data_out=16'h9f3;
17'h10537:	data_out=16'h3d3;
17'h10538:	data_out=16'h8a00;
17'h10539:	data_out=16'h89b0;
17'h1053a:	data_out=16'h9fb;
17'h1053b:	data_out=16'ha00;
17'h1053c:	data_out=16'h110;
17'h1053d:	data_out=16'h897b;
17'h1053e:	data_out=16'h9ee;
17'h1053f:	data_out=16'h4d8;
17'h10540:	data_out=16'h9f4;
17'h10541:	data_out=16'h5de;
17'h10542:	data_out=16'h89db;
17'h10543:	data_out=16'h9f9;
17'h10544:	data_out=16'h89f;
17'h10545:	data_out=16'h89b9;
17'h10546:	data_out=16'h89f3;
17'h10547:	data_out=16'h854e;
17'h10548:	data_out=16'h570;
17'h10549:	data_out=16'h9ea;
17'h1054a:	data_out=16'ha00;
17'h1054b:	data_out=16'h89d6;
17'h1054c:	data_out=16'h8834;
17'h1054d:	data_out=16'h85b4;
17'h1054e:	data_out=16'h9fc;
17'h1054f:	data_out=16'hd1;
17'h10550:	data_out=16'h9f0;
17'h10551:	data_out=16'h89c8;
17'h10552:	data_out=16'h9e8;
17'h10553:	data_out=16'h9fc;
17'h10554:	data_out=16'h8470;
17'h10555:	data_out=16'h9e6;
17'h10556:	data_out=16'h87e1;
17'h10557:	data_out=16'h89ff;
17'h10558:	data_out=16'h8906;
17'h10559:	data_out=16'h991;
17'h1055a:	data_out=16'h87a2;
17'h1055b:	data_out=16'h80e8;
17'h1055c:	data_out=16'h89fa;
17'h1055d:	data_out=16'h23c;
17'h1055e:	data_out=16'h9fd;
17'h1055f:	data_out=16'h89dc;
17'h10560:	data_out=16'h8992;
17'h10561:	data_out=16'h89f3;
17'h10562:	data_out=16'h959;
17'h10563:	data_out=16'h867d;
17'h10564:	data_out=16'h89bf;
17'h10565:	data_out=16'ha00;
17'h10566:	data_out=16'ha00;
17'h10567:	data_out=16'ha00;
17'h10568:	data_out=16'h9ed;
17'h10569:	data_out=16'h89df;
17'h1056a:	data_out=16'h9cb;
17'h1056b:	data_out=16'h9a0;
17'h1056c:	data_out=16'h89e5;
17'h1056d:	data_out=16'h8705;
17'h1056e:	data_out=16'h9cc;
17'h1056f:	data_out=16'h9ea;
17'h10570:	data_out=16'h9da;
17'h10571:	data_out=16'h861c;
17'h10572:	data_out=16'h89a4;
17'h10573:	data_out=16'h89ff;
17'h10574:	data_out=16'ha00;
17'h10575:	data_out=16'h8a00;
17'h10576:	data_out=16'ha00;
17'h10577:	data_out=16'h9f6;
17'h10578:	data_out=16'h8151;
17'h10579:	data_out=16'h897;
17'h1057a:	data_out=16'h82b5;
17'h1057b:	data_out=16'h9ee;
17'h1057c:	data_out=16'h89f8;
17'h1057d:	data_out=16'h9f0;
17'h1057e:	data_out=16'h24;
17'h1057f:	data_out=16'h89f8;
17'h10580:	data_out=16'h8a00;
17'h10581:	data_out=16'h8a00;
17'h10582:	data_out=16'h3ea;
17'h10583:	data_out=16'h8350;
17'h10584:	data_out=16'ha00;
17'h10585:	data_out=16'h984;
17'h10586:	data_out=16'h89cc;
17'h10587:	data_out=16'ha00;
17'h10588:	data_out=16'h8eb;
17'h10589:	data_out=16'h48e;
17'h1058a:	data_out=16'h8a00;
17'h1058b:	data_out=16'h9ff;
17'h1058c:	data_out=16'h9ee;
17'h1058d:	data_out=16'h89ef;
17'h1058e:	data_out=16'h9ef;
17'h1058f:	data_out=16'h6b4;
17'h10590:	data_out=16'h912;
17'h10591:	data_out=16'h89f0;
17'h10592:	data_out=16'h8a00;
17'h10593:	data_out=16'h8544;
17'h10594:	data_out=16'h845f;
17'h10595:	data_out=16'h872b;
17'h10596:	data_out=16'h8510;
17'h10597:	data_out=16'h84e2;
17'h10598:	data_out=16'h89ff;
17'h10599:	data_out=16'ha00;
17'h1059a:	data_out=16'h9cb;
17'h1059b:	data_out=16'h9dd;
17'h1059c:	data_out=16'h89f4;
17'h1059d:	data_out=16'h89fa;
17'h1059e:	data_out=16'h84fb;
17'h1059f:	data_out=16'h4f;
17'h105a0:	data_out=16'h8995;
17'h105a1:	data_out=16'h9f1;
17'h105a2:	data_out=16'h81e2;
17'h105a3:	data_out=16'h9fe;
17'h105a4:	data_out=16'h9fe;
17'h105a5:	data_out=16'h61b;
17'h105a6:	data_out=16'h8351;
17'h105a7:	data_out=16'h739;
17'h105a8:	data_out=16'h9f3;
17'h105a9:	data_out=16'h9da;
17'h105aa:	data_out=16'h577;
17'h105ab:	data_out=16'h9ff;
17'h105ac:	data_out=16'h86d1;
17'h105ad:	data_out=16'h89e4;
17'h105ae:	data_out=16'h167;
17'h105af:	data_out=16'h308;
17'h105b0:	data_out=16'ha00;
17'h105b1:	data_out=16'h89fa;
17'h105b2:	data_out=16'ha00;
17'h105b3:	data_out=16'h89c6;
17'h105b4:	data_out=16'h8a00;
17'h105b5:	data_out=16'h9c4;
17'h105b6:	data_out=16'h9fd;
17'h105b7:	data_out=16'h9b2;
17'h105b8:	data_out=16'h8a00;
17'h105b9:	data_out=16'h89d3;
17'h105ba:	data_out=16'h595;
17'h105bb:	data_out=16'ha00;
17'h105bc:	data_out=16'h828d;
17'h105bd:	data_out=16'h8610;
17'h105be:	data_out=16'h9f3;
17'h105bf:	data_out=16'h963;
17'h105c0:	data_out=16'ha00;
17'h105c1:	data_out=16'h959;
17'h105c2:	data_out=16'h89fb;
17'h105c3:	data_out=16'ha00;
17'h105c4:	data_out=16'h9c2;
17'h105c5:	data_out=16'h86e2;
17'h105c6:	data_out=16'h8a00;
17'h105c7:	data_out=16'h84c7;
17'h105c8:	data_out=16'h82db;
17'h105c9:	data_out=16'h971;
17'h105ca:	data_out=16'ha00;
17'h105cb:	data_out=16'h89f1;
17'h105cc:	data_out=16'h8578;
17'h105cd:	data_out=16'h837d;
17'h105ce:	data_out=16'h9fa;
17'h105cf:	data_out=16'h8162;
17'h105d0:	data_out=16'ha00;
17'h105d1:	data_out=16'h89e9;
17'h105d2:	data_out=16'ha00;
17'h105d3:	data_out=16'h9b5;
17'h105d4:	data_out=16'h8790;
17'h105d5:	data_out=16'h9f9;
17'h105d6:	data_out=16'h99c;
17'h105d7:	data_out=16'h84bd;
17'h105d8:	data_out=16'h821a;
17'h105d9:	data_out=16'h9ce;
17'h105da:	data_out=16'h89df;
17'h105db:	data_out=16'h9b1;
17'h105dc:	data_out=16'h89fd;
17'h105dd:	data_out=16'h274;
17'h105de:	data_out=16'h735;
17'h105df:	data_out=16'h89b6;
17'h105e0:	data_out=16'h8857;
17'h105e1:	data_out=16'h84b5;
17'h105e2:	data_out=16'ha00;
17'h105e3:	data_out=16'h88d3;
17'h105e4:	data_out=16'h8a00;
17'h105e5:	data_out=16'ha00;
17'h105e6:	data_out=16'ha00;
17'h105e7:	data_out=16'ha00;
17'h105e8:	data_out=16'h9f3;
17'h105e9:	data_out=16'h37;
17'h105ea:	data_out=16'h9ed;
17'h105eb:	data_out=16'h870;
17'h105ec:	data_out=16'h89f9;
17'h105ed:	data_out=16'h892e;
17'h105ee:	data_out=16'h9ed;
17'h105ef:	data_out=16'h9f0;
17'h105f0:	data_out=16'h9ee;
17'h105f1:	data_out=16'h815f;
17'h105f2:	data_out=16'h89d4;
17'h105f3:	data_out=16'h89fd;
17'h105f4:	data_out=16'ha00;
17'h105f5:	data_out=16'h8a00;
17'h105f6:	data_out=16'ha00;
17'h105f7:	data_out=16'ha00;
17'h105f8:	data_out=16'h663;
17'h105f9:	data_out=16'h9b6;
17'h105fa:	data_out=16'h84b0;
17'h105fb:	data_out=16'h9f3;
17'h105fc:	data_out=16'h89fc;
17'h105fd:	data_out=16'h4d4;
17'h105fe:	data_out=16'h89d8;
17'h105ff:	data_out=16'h89fe;
17'h10600:	data_out=16'h8a00;
17'h10601:	data_out=16'h8a00;
17'h10602:	data_out=16'h8062;
17'h10603:	data_out=16'h859e;
17'h10604:	data_out=16'ha00;
17'h10605:	data_out=16'h984;
17'h10606:	data_out=16'h89be;
17'h10607:	data_out=16'h9ff;
17'h10608:	data_out=16'h943;
17'h10609:	data_out=16'h8304;
17'h1060a:	data_out=16'h8999;
17'h1060b:	data_out=16'h862a;
17'h1060c:	data_out=16'h9fa;
17'h1060d:	data_out=16'h89eb;
17'h1060e:	data_out=16'h9f6;
17'h1060f:	data_out=16'h731;
17'h10610:	data_out=16'h8219;
17'h10611:	data_out=16'h286;
17'h10612:	data_out=16'h89f8;
17'h10613:	data_out=16'h8953;
17'h10614:	data_out=16'h882d;
17'h10615:	data_out=16'h8389;
17'h10616:	data_out=16'h810d;
17'h10617:	data_out=16'h8845;
17'h10618:	data_out=16'h89fc;
17'h10619:	data_out=16'ha00;
17'h1061a:	data_out=16'h9c5;
17'h1061b:	data_out=16'h81de;
17'h1061c:	data_out=16'h89fa;
17'h1061d:	data_out=16'h8a00;
17'h1061e:	data_out=16'h8653;
17'h1061f:	data_out=16'h838c;
17'h10620:	data_out=16'h87f5;
17'h10621:	data_out=16'h9f8;
17'h10622:	data_out=16'h855e;
17'h10623:	data_out=16'h9f8;
17'h10624:	data_out=16'h9f8;
17'h10625:	data_out=16'hd0;
17'h10626:	data_out=16'h8801;
17'h10627:	data_out=16'h974;
17'h10628:	data_out=16'h9f8;
17'h10629:	data_out=16'h9d9;
17'h1062a:	data_out=16'h572;
17'h1062b:	data_out=16'ha00;
17'h1062c:	data_out=16'h82fd;
17'h1062d:	data_out=16'h8a00;
17'h1062e:	data_out=16'h80e7;
17'h1062f:	data_out=16'h805c;
17'h10630:	data_out=16'ha00;
17'h10631:	data_out=16'h89f3;
17'h10632:	data_out=16'h9ff;
17'h10633:	data_out=16'h89a8;
17'h10634:	data_out=16'h8a00;
17'h10635:	data_out=16'h99e;
17'h10636:	data_out=16'h9fc;
17'h10637:	data_out=16'h166;
17'h10638:	data_out=16'h8a00;
17'h10639:	data_out=16'h89e4;
17'h1063a:	data_out=16'h8192;
17'h1063b:	data_out=16'ha00;
17'h1063c:	data_out=16'h8967;
17'h1063d:	data_out=16'h83b0;
17'h1063e:	data_out=16'h9f8;
17'h1063f:	data_out=16'h981;
17'h10640:	data_out=16'ha00;
17'h10641:	data_out=16'h98e;
17'h10642:	data_out=16'h89d8;
17'h10643:	data_out=16'h9fb;
17'h10644:	data_out=16'h9d3;
17'h10645:	data_out=16'h8338;
17'h10646:	data_out=16'h8a00;
17'h10647:	data_out=16'h848a;
17'h10648:	data_out=16'h88e1;
17'h10649:	data_out=16'h29a;
17'h1064a:	data_out=16'ha00;
17'h1064b:	data_out=16'h89d2;
17'h1064c:	data_out=16'h852e;
17'h1064d:	data_out=16'h8598;
17'h1064e:	data_out=16'h692;
17'h1064f:	data_out=16'h83ea;
17'h10650:	data_out=16'h5b5;
17'h10651:	data_out=16'h88c9;
17'h10652:	data_out=16'h9fd;
17'h10653:	data_out=16'h9b3;
17'h10654:	data_out=16'h86f6;
17'h10655:	data_out=16'h238;
17'h10656:	data_out=16'h9f0;
17'h10657:	data_out=16'h8478;
17'h10658:	data_out=16'h44;
17'h10659:	data_out=16'h6ae;
17'h1065a:	data_out=16'h89e8;
17'h1065b:	data_out=16'h9d7;
17'h1065c:	data_out=16'h89fe;
17'h1065d:	data_out=16'h533;
17'h1065e:	data_out=16'h15a;
17'h1065f:	data_out=16'h8920;
17'h10660:	data_out=16'h89da;
17'h10661:	data_out=16'h99f;
17'h10662:	data_out=16'h22a;
17'h10663:	data_out=16'h8973;
17'h10664:	data_out=16'h8a00;
17'h10665:	data_out=16'ha00;
17'h10666:	data_out=16'ha00;
17'h10667:	data_out=16'ha00;
17'h10668:	data_out=16'h9f8;
17'h10669:	data_out=16'h29b;
17'h1066a:	data_out=16'h9f3;
17'h1066b:	data_out=16'h8e8;
17'h1066c:	data_out=16'h89cc;
17'h1066d:	data_out=16'h897b;
17'h1066e:	data_out=16'h9f3;
17'h1066f:	data_out=16'h9e8;
17'h10670:	data_out=16'h9f5;
17'h10671:	data_out=16'h8131;
17'h10672:	data_out=16'h891a;
17'h10673:	data_out=16'h873f;
17'h10674:	data_out=16'h9fb;
17'h10675:	data_out=16'h8a00;
17'h10676:	data_out=16'ha00;
17'h10677:	data_out=16'ha00;
17'h10678:	data_out=16'h614;
17'h10679:	data_out=16'h9e1;
17'h1067a:	data_out=16'h88ad;
17'h1067b:	data_out=16'h9f8;
17'h1067c:	data_out=16'h89fe;
17'h1067d:	data_out=16'h839d;
17'h1067e:	data_out=16'h89f3;
17'h1067f:	data_out=16'h8997;
17'h10680:	data_out=16'h8791;
17'h10681:	data_out=16'h8a00;
17'h10682:	data_out=16'h8786;
17'h10683:	data_out=16'h89ed;
17'h10684:	data_out=16'ha00;
17'h10685:	data_out=16'h9d3;
17'h10686:	data_out=16'h89ec;
17'h10687:	data_out=16'h9fc;
17'h10688:	data_out=16'h750;
17'h10689:	data_out=16'h8824;
17'h1068a:	data_out=16'h961;
17'h1068b:	data_out=16'h871c;
17'h1068c:	data_out=16'h9e8;
17'h1068d:	data_out=16'h89ec;
17'h1068e:	data_out=16'h4ba;
17'h1068f:	data_out=16'h8306;
17'h10690:	data_out=16'h89f2;
17'h10691:	data_out=16'h985;
17'h10692:	data_out=16'h89f7;
17'h10693:	data_out=16'h89e2;
17'h10694:	data_out=16'h89b1;
17'h10695:	data_out=16'h8499;
17'h10696:	data_out=16'h833a;
17'h10697:	data_out=16'h89cd;
17'h10698:	data_out=16'h89e0;
17'h10699:	data_out=16'ha00;
17'h1069a:	data_out=16'ha00;
17'h1069b:	data_out=16'h898b;
17'h1069c:	data_out=16'h89fd;
17'h1069d:	data_out=16'h81af;
17'h1069e:	data_out=16'h8990;
17'h1069f:	data_out=16'h85d8;
17'h106a0:	data_out=16'h8328;
17'h106a1:	data_out=16'h513;
17'h106a2:	data_out=16'h8959;
17'h106a3:	data_out=16'h32f;
17'h106a4:	data_out=16'h358;
17'h106a5:	data_out=16'h85b8;
17'h106a6:	data_out=16'h899d;
17'h106a7:	data_out=16'h9bc;
17'h106a8:	data_out=16'h5dd;
17'h106a9:	data_out=16'h71e;
17'h106aa:	data_out=16'h8271;
17'h106ab:	data_out=16'ha00;
17'h106ac:	data_out=16'h8411;
17'h106ad:	data_out=16'h8a00;
17'h106ae:	data_out=16'h872b;
17'h106af:	data_out=16'h84f0;
17'h106b0:	data_out=16'h9fb;
17'h106b1:	data_out=16'h7c2;
17'h106b2:	data_out=16'h9fa;
17'h106b3:	data_out=16'h89e7;
17'h106b4:	data_out=16'h8a00;
17'h106b5:	data_out=16'h9cd;
17'h106b6:	data_out=16'h8046;
17'h106b7:	data_out=16'h86e7;
17'h106b8:	data_out=16'h8a00;
17'h106b9:	data_out=16'h89ef;
17'h106ba:	data_out=16'h873f;
17'h106bb:	data_out=16'ha00;
17'h106bc:	data_out=16'h89f7;
17'h106bd:	data_out=16'h8431;
17'h106be:	data_out=16'h5e4;
17'h106bf:	data_out=16'h9d0;
17'h106c0:	data_out=16'ha00;
17'h106c1:	data_out=16'h6c9;
17'h106c2:	data_out=16'h89c4;
17'h106c3:	data_out=16'ha00;
17'h106c4:	data_out=16'ha00;
17'h106c5:	data_out=16'h846b;
17'h106c6:	data_out=16'h8a00;
17'h106c7:	data_out=16'h8766;
17'h106c8:	data_out=16'h89d5;
17'h106c9:	data_out=16'h849a;
17'h106ca:	data_out=16'ha00;
17'h106cb:	data_out=16'h8274;
17'h106cc:	data_out=16'h8886;
17'h106cd:	data_out=16'h89b9;
17'h106ce:	data_out=16'h32f;
17'h106cf:	data_out=16'h87df;
17'h106d0:	data_out=16'h83c6;
17'h106d1:	data_out=16'h89d1;
17'h106d2:	data_out=16'h324;
17'h106d3:	data_out=16'ha00;
17'h106d4:	data_out=16'h88c1;
17'h106d5:	data_out=16'h877c;
17'h106d6:	data_out=16'h9ed;
17'h106d7:	data_out=16'h87fa;
17'h106d8:	data_out=16'h89ea;
17'h106d9:	data_out=16'h969;
17'h106da:	data_out=16'h89eb;
17'h106db:	data_out=16'ha00;
17'h106dc:	data_out=16'h8092;
17'h106dd:	data_out=16'he9;
17'h106de:	data_out=16'h84a1;
17'h106df:	data_out=16'h89bb;
17'h106e0:	data_out=16'h89de;
17'h106e1:	data_out=16'h9de;
17'h106e2:	data_out=16'h8823;
17'h106e3:	data_out=16'h89d1;
17'h106e4:	data_out=16'h89fe;
17'h106e5:	data_out=16'h9f0;
17'h106e6:	data_out=16'ha00;
17'h106e7:	data_out=16'ha00;
17'h106e8:	data_out=16'h55c;
17'h106e9:	data_out=16'haa;
17'h106ea:	data_out=16'h44a;
17'h106eb:	data_out=16'h99e;
17'h106ec:	data_out=16'h86b7;
17'h106ed:	data_out=16'h89d8;
17'h106ee:	data_out=16'h44d;
17'h106ef:	data_out=16'ha00;
17'h106f0:	data_out=16'h492;
17'h106f1:	data_out=16'h8448;
17'h106f2:	data_out=16'h89f8;
17'h106f3:	data_out=16'h8095;
17'h106f4:	data_out=16'h9ab;
17'h106f5:	data_out=16'h89e8;
17'h106f6:	data_out=16'ha00;
17'h106f7:	data_out=16'h8410;
17'h106f8:	data_out=16'h7b2;
17'h106f9:	data_out=16'h9f3;
17'h106fa:	data_out=16'h89b2;
17'h106fb:	data_out=16'h5e5;
17'h106fc:	data_out=16'h89b0;
17'h106fd:	data_out=16'h810b;
17'h106fe:	data_out=16'h8a00;
17'h106ff:	data_out=16'h873f;
17'h10700:	data_out=16'h8643;
17'h10701:	data_out=16'h840;
17'h10702:	data_out=16'h89e2;
17'h10703:	data_out=16'h89fb;
17'h10704:	data_out=16'ha00;
17'h10705:	data_out=16'h9ff;
17'h10706:	data_out=16'h89ff;
17'h10707:	data_out=16'h9c4;
17'h10708:	data_out=16'h89f9;
17'h10709:	data_out=16'h89fd;
17'h1070a:	data_out=16'h9fd;
17'h1070b:	data_out=16'h411;
17'h1070c:	data_out=16'h9a3;
17'h1070d:	data_out=16'h89ff;
17'h1070e:	data_out=16'h46;
17'h1070f:	data_out=16'h89f4;
17'h10710:	data_out=16'h89fb;
17'h10711:	data_out=16'h9ea;
17'h10712:	data_out=16'h89fe;
17'h10713:	data_out=16'h89fa;
17'h10714:	data_out=16'h89fa;
17'h10715:	data_out=16'h817d;
17'h10716:	data_out=16'h893c;
17'h10717:	data_out=16'h89fd;
17'h10718:	data_out=16'h89fa;
17'h10719:	data_out=16'ha00;
17'h1071a:	data_out=16'ha00;
17'h1071b:	data_out=16'h89fc;
17'h1071c:	data_out=16'h89fe;
17'h1071d:	data_out=16'h7da;
17'h1071e:	data_out=16'h89f9;
17'h1071f:	data_out=16'h893d;
17'h10720:	data_out=16'h8014;
17'h10721:	data_out=16'h25;
17'h10722:	data_out=16'h2f1;
17'h10723:	data_out=16'h11e;
17'h10724:	data_out=16'h140;
17'h10725:	data_out=16'h89dd;
17'h10726:	data_out=16'h89ed;
17'h10727:	data_out=16'h9cc;
17'h10728:	data_out=16'h1a;
17'h10729:	data_out=16'h8663;
17'h1072a:	data_out=16'h89f3;
17'h1072b:	data_out=16'ha00;
17'h1072c:	data_out=16'h8887;
17'h1072d:	data_out=16'h8a00;
17'h1072e:	data_out=16'h89db;
17'h1072f:	data_out=16'h8968;
17'h10730:	data_out=16'h9f7;
17'h10731:	data_out=16'h9d7;
17'h10732:	data_out=16'h9f5;
17'h10733:	data_out=16'h89f9;
17'h10734:	data_out=16'h8a00;
17'h10735:	data_out=16'h9ee;
17'h10736:	data_out=16'h89f4;
17'h10737:	data_out=16'h89e0;
17'h10738:	data_out=16'h856f;
17'h10739:	data_out=16'h89f8;
17'h1073a:	data_out=16'h89fb;
17'h1073b:	data_out=16'h9ff;
17'h1073c:	data_out=16'h89ef;
17'h1073d:	data_out=16'h80af;
17'h1073e:	data_out=16'h16;
17'h1073f:	data_out=16'h9ff;
17'h10740:	data_out=16'ha00;
17'h10741:	data_out=16'h884c;
17'h10742:	data_out=16'h8a00;
17'h10743:	data_out=16'h8177;
17'h10744:	data_out=16'ha00;
17'h10745:	data_out=16'h8242;
17'h10746:	data_out=16'h8a00;
17'h10747:	data_out=16'h89dd;
17'h10748:	data_out=16'h89fd;
17'h10749:	data_out=16'h8919;
17'h1074a:	data_out=16'h9e1;
17'h1074b:	data_out=16'h947;
17'h1074c:	data_out=16'h89de;
17'h1074d:	data_out=16'h6c8;
17'h1074e:	data_out=16'h27a;
17'h1074f:	data_out=16'h89ff;
17'h10750:	data_out=16'h8743;
17'h10751:	data_out=16'h89ec;
17'h10752:	data_out=16'h9fa;
17'h10753:	data_out=16'h9fa;
17'h10754:	data_out=16'h873e;
17'h10755:	data_out=16'h89e0;
17'h10756:	data_out=16'h11c;
17'h10757:	data_out=16'h88f8;
17'h10758:	data_out=16'h89f7;
17'h10759:	data_out=16'h9e4;
17'h1075a:	data_out=16'h8a00;
17'h1075b:	data_out=16'ha00;
17'h1075c:	data_out=16'h5f8;
17'h1075d:	data_out=16'h85e8;
17'h1075e:	data_out=16'h89ac;
17'h1075f:	data_out=16'h89f8;
17'h10760:	data_out=16'h89fe;
17'h10761:	data_out=16'ha00;
17'h10762:	data_out=16'h89fa;
17'h10763:	data_out=16'h89f9;
17'h10764:	data_out=16'h8743;
17'h10765:	data_out=16'h9d3;
17'h10766:	data_out=16'ha00;
17'h10767:	data_out=16'ha00;
17'h10768:	data_out=16'h27;
17'h10769:	data_out=16'h89fe;
17'h1076a:	data_out=16'h3d;
17'h1076b:	data_out=16'h998;
17'h1076c:	data_out=16'h8685;
17'h1076d:	data_out=16'h89f9;
17'h1076e:	data_out=16'h3d;
17'h1076f:	data_out=16'h9f7;
17'h10770:	data_out=16'h43;
17'h10771:	data_out=16'h89f1;
17'h10772:	data_out=16'h892;
17'h10773:	data_out=16'ha00;
17'h10774:	data_out=16'h993;
17'h10775:	data_out=16'h89c5;
17'h10776:	data_out=16'ha00;
17'h10777:	data_out=16'h89fa;
17'h10778:	data_out=16'h8066;
17'h10779:	data_out=16'h23;
17'h1077a:	data_out=16'h89fa;
17'h1077b:	data_out=16'h12;
17'h1077c:	data_out=16'h89f3;
17'h1077d:	data_out=16'h8204;
17'h1077e:	data_out=16'h8a00;
17'h1077f:	data_out=16'h89e7;
17'h10780:	data_out=16'h9ce;
17'h10781:	data_out=16'h8ec;
17'h10782:	data_out=16'h89fd;
17'h10783:	data_out=16'h8a00;
17'h10784:	data_out=16'ha00;
17'h10785:	data_out=16'h9f8;
17'h10786:	data_out=16'h8a00;
17'h10787:	data_out=16'h3a;
17'h10788:	data_out=16'h89fe;
17'h10789:	data_out=16'h8386;
17'h1078a:	data_out=16'ha00;
17'h1078b:	data_out=16'h88be;
17'h1078c:	data_out=16'h88cb;
17'h1078d:	data_out=16'h8a00;
17'h1078e:	data_out=16'h168;
17'h1078f:	data_out=16'h89ff;
17'h10790:	data_out=16'h82d2;
17'h10791:	data_out=16'ha00;
17'h10792:	data_out=16'h89ff;
17'h10793:	data_out=16'h89ef;
17'h10794:	data_out=16'h8a00;
17'h10795:	data_out=16'h9fe;
17'h10796:	data_out=16'h87a9;
17'h10797:	data_out=16'h8a00;
17'h10798:	data_out=16'h89f4;
17'h10799:	data_out=16'ha00;
17'h1079a:	data_out=16'ha00;
17'h1079b:	data_out=16'h8a00;
17'h1079c:	data_out=16'h82a0;
17'h1079d:	data_out=16'h9d0;
17'h1079e:	data_out=16'h89f8;
17'h1079f:	data_out=16'h85f2;
17'h107a0:	data_out=16'ha00;
17'h107a1:	data_out=16'hf7;
17'h107a2:	data_out=16'h9ff;
17'h107a3:	data_out=16'h8a1;
17'h107a4:	data_out=16'h8b1;
17'h107a5:	data_out=16'hba;
17'h107a6:	data_out=16'h89fe;
17'h107a7:	data_out=16'h9fa;
17'h107a8:	data_out=16'h3e;
17'h107a9:	data_out=16'h88bb;
17'h107aa:	data_out=16'h89fe;
17'h107ab:	data_out=16'ha00;
17'h107ac:	data_out=16'h69f;
17'h107ad:	data_out=16'h8a00;
17'h107ae:	data_out=16'h89fc;
17'h107af:	data_out=16'h88d6;
17'h107b0:	data_out=16'h9dd;
17'h107b1:	data_out=16'h9f3;
17'h107b2:	data_out=16'h9eb;
17'h107b3:	data_out=16'h89fc;
17'h107b4:	data_out=16'h4b3;
17'h107b5:	data_out=16'ha00;
17'h107b6:	data_out=16'h89fd;
17'h107b7:	data_out=16'h89fb;
17'h107b8:	data_out=16'h8e6;
17'h107b9:	data_out=16'h89f8;
17'h107ba:	data_out=16'h88a;
17'h107bb:	data_out=16'h9cf;
17'h107bc:	data_out=16'h89f8;
17'h107bd:	data_out=16'h9ff;
17'h107be:	data_out=16'h34;
17'h107bf:	data_out=16'h9f8;
17'h107c0:	data_out=16'ha00;
17'h107c1:	data_out=16'h89fd;
17'h107c2:	data_out=16'h8a00;
17'h107c3:	data_out=16'h86b0;
17'h107c4:	data_out=16'ha00;
17'h107c5:	data_out=16'h9fd;
17'h107c6:	data_out=16'h8a00;
17'h107c7:	data_out=16'he1;
17'h107c8:	data_out=16'h8a00;
17'h107c9:	data_out=16'h4df;
17'h107ca:	data_out=16'h39;
17'h107cb:	data_out=16'h844a;
17'h107cc:	data_out=16'h8632;
17'h107cd:	data_out=16'h9ff;
17'h107ce:	data_out=16'h818c;
17'h107cf:	data_out=16'h16d;
17'h107d0:	data_out=16'h8f2;
17'h107d1:	data_out=16'h89f6;
17'h107d2:	data_out=16'h9ec;
17'h107d3:	data_out=16'h824a;
17'h107d4:	data_out=16'h9d7;
17'h107d5:	data_out=16'h89fd;
17'h107d6:	data_out=16'h688;
17'h107d7:	data_out=16'ha00;
17'h107d8:	data_out=16'h8a00;
17'h107d9:	data_out=16'ha00;
17'h107da:	data_out=16'h8a00;
17'h107db:	data_out=16'ha00;
17'h107dc:	data_out=16'h402;
17'h107dd:	data_out=16'h82c0;
17'h107de:	data_out=16'h88b7;
17'h107df:	data_out=16'h878f;
17'h107e0:	data_out=16'h89ff;
17'h107e1:	data_out=16'h9fd;
17'h107e2:	data_out=16'h8a00;
17'h107e3:	data_out=16'h8a00;
17'h107e4:	data_out=16'h9da;
17'h107e5:	data_out=16'h9e8;
17'h107e6:	data_out=16'ha00;
17'h107e7:	data_out=16'ha00;
17'h107e8:	data_out=16'hc5;
17'h107e9:	data_out=16'h89ff;
17'h107ea:	data_out=16'h1b7;
17'h107eb:	data_out=16'h9fa;
17'h107ec:	data_out=16'h6b2;
17'h107ed:	data_out=16'h8a00;
17'h107ee:	data_out=16'h1b4;
17'h107ef:	data_out=16'h45d;
17'h107f0:	data_out=16'h182;
17'h107f1:	data_out=16'h89fe;
17'h107f2:	data_out=16'ha00;
17'h107f3:	data_out=16'ha00;
17'h107f4:	data_out=16'h8ec;
17'h107f5:	data_out=16'h89d6;
17'h107f6:	data_out=16'ha00;
17'h107f7:	data_out=16'h8646;
17'h107f8:	data_out=16'h8503;
17'h107f9:	data_out=16'h8867;
17'h107fa:	data_out=16'h8a00;
17'h107fb:	data_out=16'h2e;
17'h107fc:	data_out=16'h8757;
17'h107fd:	data_out=16'h3e7;
17'h107fe:	data_out=16'h8a00;
17'h107ff:	data_out=16'ha00;
17'h10800:	data_out=16'ha00;
17'h10801:	data_out=16'h9ff;
17'h10802:	data_out=16'h8a00;
17'h10803:	data_out=16'h8016;
17'h10804:	data_out=16'ha00;
17'h10805:	data_out=16'h9f8;
17'h10806:	data_out=16'h8a00;
17'h10807:	data_out=16'h8a00;
17'h10808:	data_out=16'h89ff;
17'h10809:	data_out=16'h9ab;
17'h1080a:	data_out=16'ha00;
17'h1080b:	data_out=16'h89fe;
17'h1080c:	data_out=16'h8a00;
17'h1080d:	data_out=16'h8a00;
17'h1080e:	data_out=16'h299;
17'h1080f:	data_out=16'h8a00;
17'h10810:	data_out=16'ha00;
17'h10811:	data_out=16'ha00;
17'h10812:	data_out=16'h89ff;
17'h10813:	data_out=16'h8335;
17'h10814:	data_out=16'h8a00;
17'h10815:	data_out=16'ha00;
17'h10816:	data_out=16'h9d6;
17'h10817:	data_out=16'h8a00;
17'h10818:	data_out=16'h25d;
17'h10819:	data_out=16'ha00;
17'h1081a:	data_out=16'ha00;
17'h1081b:	data_out=16'h8a00;
17'h1081c:	data_out=16'h6a2;
17'h1081d:	data_out=16'ha00;
17'h1081e:	data_out=16'h820e;
17'h1081f:	data_out=16'h115;
17'h10820:	data_out=16'ha00;
17'h10821:	data_out=16'h1fd;
17'h10822:	data_out=16'h9fe;
17'h10823:	data_out=16'h814c;
17'h10824:	data_out=16'h8134;
17'h10825:	data_out=16'ha00;
17'h10826:	data_out=16'h89ff;
17'h10827:	data_out=16'ha00;
17'h10828:	data_out=16'h104;
17'h10829:	data_out=16'h8a00;
17'h1082a:	data_out=16'h89fe;
17'h1082b:	data_out=16'ha00;
17'h1082c:	data_out=16'ha00;
17'h1082d:	data_out=16'h83a9;
17'h1082e:	data_out=16'h8a00;
17'h1082f:	data_out=16'h9f3;
17'h10830:	data_out=16'h970;
17'h10831:	data_out=16'ha00;
17'h10832:	data_out=16'h9ac;
17'h10833:	data_out=16'h8475;
17'h10834:	data_out=16'h98c;
17'h10835:	data_out=16'ha00;
17'h10836:	data_out=16'h89ee;
17'h10837:	data_out=16'h8a00;
17'h10838:	data_out=16'ha00;
17'h10839:	data_out=16'had;
17'h1083a:	data_out=16'ha00;
17'h1083b:	data_out=16'h702;
17'h1083c:	data_out=16'h8a00;
17'h1083d:	data_out=16'ha00;
17'h1083e:	data_out=16'hf9;
17'h1083f:	data_out=16'h9fc;
17'h10840:	data_out=16'ha00;
17'h10841:	data_out=16'h89ff;
17'h10842:	data_out=16'h8946;
17'h10843:	data_out=16'h89f5;
17'h10844:	data_out=16'ha00;
17'h10845:	data_out=16'ha00;
17'h10846:	data_out=16'h8a00;
17'h10847:	data_out=16'h9f8;
17'h10848:	data_out=16'h8833;
17'h10849:	data_out=16'ha00;
17'h1084a:	data_out=16'h8a00;
17'h1084b:	data_out=16'h8a00;
17'h1084c:	data_out=16'h8059;
17'h1084d:	data_out=16'ha00;
17'h1084e:	data_out=16'h87a8;
17'h1084f:	data_out=16'h9f9;
17'h10850:	data_out=16'h9ff;
17'h10851:	data_out=16'h8a00;
17'h10852:	data_out=16'h9fd;
17'h10853:	data_out=16'h892b;
17'h10854:	data_out=16'ha00;
17'h10855:	data_out=16'h8a00;
17'h10856:	data_out=16'h9e5;
17'h10857:	data_out=16'ha00;
17'h10858:	data_out=16'h8a00;
17'h10859:	data_out=16'ha00;
17'h1085a:	data_out=16'h8a00;
17'h1085b:	data_out=16'ha00;
17'h1085c:	data_out=16'h2fd;
17'h1085d:	data_out=16'ha00;
17'h1085e:	data_out=16'h9be;
17'h1085f:	data_out=16'ha00;
17'h10860:	data_out=16'h8a00;
17'h10861:	data_out=16'ha00;
17'h10862:	data_out=16'h8a00;
17'h10863:	data_out=16'h897e;
17'h10864:	data_out=16'ha00;
17'h10865:	data_out=16'ha00;
17'h10866:	data_out=16'ha00;
17'h10867:	data_out=16'ha00;
17'h10868:	data_out=16'h1aa;
17'h10869:	data_out=16'h8a00;
17'h1086a:	data_out=16'h305;
17'h1086b:	data_out=16'ha00;
17'h1086c:	data_out=16'ha00;
17'h1086d:	data_out=16'h870f;
17'h1086e:	data_out=16'h302;
17'h1086f:	data_out=16'h78f;
17'h10870:	data_out=16'h2be;
17'h10871:	data_out=16'h8a00;
17'h10872:	data_out=16'ha00;
17'h10873:	data_out=16'ha00;
17'h10874:	data_out=16'h7c5;
17'h10875:	data_out=16'h8a00;
17'h10876:	data_out=16'ha00;
17'h10877:	data_out=16'h973;
17'h10878:	data_out=16'h868d;
17'h10879:	data_out=16'h8886;
17'h1087a:	data_out=16'h8a00;
17'h1087b:	data_out=16'hf2;
17'h1087c:	data_out=16'h720;
17'h1087d:	data_out=16'h5f7;
17'h1087e:	data_out=16'h81e;
17'h1087f:	data_out=16'ha00;
17'h10880:	data_out=16'ha00;
17'h10881:	data_out=16'ha00;
17'h10882:	data_out=16'h8a00;
17'h10883:	data_out=16'h9fd;
17'h10884:	data_out=16'ha00;
17'h10885:	data_out=16'h9da;
17'h10886:	data_out=16'h9fe;
17'h10887:	data_out=16'h8125;
17'h10888:	data_out=16'h8a00;
17'h10889:	data_out=16'ha00;
17'h1088a:	data_out=16'ha00;
17'h1088b:	data_out=16'h8387;
17'h1088c:	data_out=16'h8a00;
17'h1088d:	data_out=16'h8a00;
17'h1088e:	data_out=16'h8168;
17'h1088f:	data_out=16'h89ff;
17'h10890:	data_out=16'ha00;
17'h10891:	data_out=16'ha00;
17'h10892:	data_out=16'h824c;
17'h10893:	data_out=16'ha00;
17'h10894:	data_out=16'h973;
17'h10895:	data_out=16'ha00;
17'h10896:	data_out=16'ha00;
17'h10897:	data_out=16'h8401;
17'h10898:	data_out=16'h81b3;
17'h10899:	data_out=16'ha00;
17'h1089a:	data_out=16'ha00;
17'h1089b:	data_out=16'h88f7;
17'h1089c:	data_out=16'h9e9;
17'h1089d:	data_out=16'ha00;
17'h1089e:	data_out=16'ha00;
17'h1089f:	data_out=16'ha00;
17'h108a0:	data_out=16'ha00;
17'h108a1:	data_out=16'h8178;
17'h108a2:	data_out=16'h9ff;
17'h108a3:	data_out=16'h8a00;
17'h108a4:	data_out=16'h8a00;
17'h108a5:	data_out=16'ha00;
17'h108a6:	data_out=16'h8681;
17'h108a7:	data_out=16'ha00;
17'h108a8:	data_out=16'h817f;
17'h108a9:	data_out=16'h75c;
17'h108aa:	data_out=16'h882f;
17'h108ab:	data_out=16'ha00;
17'h108ac:	data_out=16'ha00;
17'h108ad:	data_out=16'h9fd;
17'h108ae:	data_out=16'h89ff;
17'h108af:	data_out=16'ha00;
17'h108b0:	data_out=16'h81b5;
17'h108b1:	data_out=16'ha00;
17'h108b2:	data_out=16'h304;
17'h108b3:	data_out=16'ha00;
17'h108b4:	data_out=16'ha00;
17'h108b5:	data_out=16'h580;
17'h108b6:	data_out=16'h864a;
17'h108b7:	data_out=16'h8a00;
17'h108b8:	data_out=16'ha00;
17'h108b9:	data_out=16'ha00;
17'h108ba:	data_out=16'ha00;
17'h108bb:	data_out=16'h36a;
17'h108bc:	data_out=16'h8a00;
17'h108bd:	data_out=16'ha00;
17'h108be:	data_out=16'h8181;
17'h108bf:	data_out=16'h9de;
17'h108c0:	data_out=16'ha00;
17'h108c1:	data_out=16'h8a00;
17'h108c2:	data_out=16'h827a;
17'h108c3:	data_out=16'ha00;
17'h108c4:	data_out=16'ha00;
17'h108c5:	data_out=16'ha00;
17'h108c6:	data_out=16'h8a00;
17'h108c7:	data_out=16'ha00;
17'h108c8:	data_out=16'ha00;
17'h108c9:	data_out=16'ha00;
17'h108ca:	data_out=16'h80d5;
17'h108cb:	data_out=16'h8909;
17'h108cc:	data_out=16'h9fa;
17'h108cd:	data_out=16'ha00;
17'h108ce:	data_out=16'h88e5;
17'h108cf:	data_out=16'h9fd;
17'h108d0:	data_out=16'ha00;
17'h108d1:	data_out=16'h8a00;
17'h108d2:	data_out=16'h8617;
17'h108d3:	data_out=16'h9fd;
17'h108d4:	data_out=16'ha00;
17'h108d5:	data_out=16'h8a00;
17'h108d6:	data_out=16'h9e4;
17'h108d7:	data_out=16'ha00;
17'h108d8:	data_out=16'h8a00;
17'h108d9:	data_out=16'ha00;
17'h108da:	data_out=16'h8a00;
17'h108db:	data_out=16'ha00;
17'h108dc:	data_out=16'h744;
17'h108dd:	data_out=16'ha00;
17'h108de:	data_out=16'ha00;
17'h108df:	data_out=16'h8d1;
17'h108e0:	data_out=16'h8a00;
17'h108e1:	data_out=16'ha00;
17'h108e2:	data_out=16'h896c;
17'h108e3:	data_out=16'ha00;
17'h108e4:	data_out=16'ha00;
17'h108e5:	data_out=16'ha00;
17'h108e6:	data_out=16'ha00;
17'h108e7:	data_out=16'ha00;
17'h108e8:	data_out=16'h8175;
17'h108e9:	data_out=16'h8a00;
17'h108ea:	data_out=16'h8177;
17'h108eb:	data_out=16'ha00;
17'h108ec:	data_out=16'ha00;
17'h108ed:	data_out=16'ha00;
17'h108ee:	data_out=16'h818d;
17'h108ef:	data_out=16'h93e;
17'h108f0:	data_out=16'h8169;
17'h108f1:	data_out=16'h8a00;
17'h108f2:	data_out=16'ha00;
17'h108f3:	data_out=16'ha00;
17'h108f4:	data_out=16'h83a5;
17'h108f5:	data_out=16'h8a00;
17'h108f6:	data_out=16'ha00;
17'h108f7:	data_out=16'h9fb;
17'h108f8:	data_out=16'h9fe;
17'h108f9:	data_out=16'h877d;
17'h108fa:	data_out=16'h9ff;
17'h108fb:	data_out=16'h8184;
17'h108fc:	data_out=16'h8027;
17'h108fd:	data_out=16'ha00;
17'h108fe:	data_out=16'ha00;
17'h108ff:	data_out=16'ha00;
17'h10900:	data_out=16'h7cc;
17'h10901:	data_out=16'h3e8;
17'h10902:	data_out=16'h10d;
17'h10903:	data_out=16'h574;
17'h10904:	data_out=16'h27a;
17'h10905:	data_out=16'h1eb;
17'h10906:	data_out=16'h9c;
17'h10907:	data_out=16'h314;
17'h10908:	data_out=16'h109;
17'h10909:	data_out=16'h7f0;
17'h1090a:	data_out=16'h2d9;
17'h1090b:	data_out=16'h257;
17'h1090c:	data_out=16'h831b;
17'h1090d:	data_out=16'h2d5;
17'h1090e:	data_out=16'h9c;
17'h1090f:	data_out=16'h222;
17'h10910:	data_out=16'h772;
17'h10911:	data_out=16'h2c0;
17'h10912:	data_out=16'h646;
17'h10913:	data_out=16'h5f2;
17'h10914:	data_out=16'h37a;
17'h10915:	data_out=16'h2b3;
17'h10916:	data_out=16'h2b8;
17'h10917:	data_out=16'h2e9;
17'h10918:	data_out=16'h11f;
17'h10919:	data_out=16'h2b;
17'h1091a:	data_out=16'h289;
17'h1091b:	data_out=16'h476;
17'h1091c:	data_out=16'h3fb;
17'h1091d:	data_out=16'h529;
17'h1091e:	data_out=16'h4dd;
17'h1091f:	data_out=16'h248;
17'h10920:	data_out=16'ha00;
17'h10921:	data_out=16'h9e;
17'h10922:	data_out=16'h944;
17'h10923:	data_out=16'h8369;
17'h10924:	data_out=16'h836a;
17'h10925:	data_out=16'h515;
17'h10926:	data_out=16'h46a;
17'h10927:	data_out=16'h4e0;
17'h10928:	data_out=16'hc1;
17'h10929:	data_out=16'h703;
17'h1092a:	data_out=16'h504;
17'h1092b:	data_out=16'h589;
17'h1092c:	data_out=16'h2d5;
17'h1092d:	data_out=16'h629;
17'h1092e:	data_out=16'h48d;
17'h1092f:	data_out=16'h6b4;
17'h10930:	data_out=16'h4f;
17'h10931:	data_out=16'h46a;
17'h10932:	data_out=16'h9c;
17'h10933:	data_out=16'h48e;
17'h10934:	data_out=16'h455;
17'h10935:	data_out=16'h823c;
17'h10936:	data_out=16'h1cc;
17'h10937:	data_out=16'h11e;
17'h10938:	data_out=16'h6ce;
17'h10939:	data_out=16'h4af;
17'h1093a:	data_out=16'h8c3;
17'h1093b:	data_out=16'h145;
17'h1093c:	data_out=16'h54;
17'h1093d:	data_out=16'h9dc;
17'h1093e:	data_out=16'hce;
17'h1093f:	data_out=16'h16b;
17'h10940:	data_out=16'h57c;
17'h10941:	data_out=16'h80ac;
17'h10942:	data_out=16'h3e6;
17'h10943:	data_out=16'h104;
17'h10944:	data_out=16'h2b9;
17'h10945:	data_out=16'h2be;
17'h10946:	data_out=16'h399;
17'h10947:	data_out=16'h710;
17'h10948:	data_out=16'h643;
17'h10949:	data_out=16'h550;
17'h1094a:	data_out=16'h2d8;
17'h1094b:	data_out=16'h80c9;
17'h1094c:	data_out=16'h4a2;
17'h1094d:	data_out=16'h973;
17'h1094e:	data_out=16'h50e;
17'h1094f:	data_out=16'h470;
17'h10950:	data_out=16'h5a6;
17'h10951:	data_out=16'h8206;
17'h10952:	data_out=16'h81d9;
17'h10953:	data_out=16'h544;
17'h10954:	data_out=16'h7b1;
17'h10955:	data_out=16'h833f;
17'h10956:	data_out=16'h590;
17'h10957:	data_out=16'h6b4;
17'h10958:	data_out=16'h82d9;
17'h10959:	data_out=16'h60b;
17'h1095a:	data_out=16'he0;
17'h1095b:	data_out=16'h80b2;
17'h1095c:	data_out=16'h176;
17'h1095d:	data_out=16'h5d0;
17'h1095e:	data_out=16'h6e6;
17'h1095f:	data_out=16'h2d0;
17'h10960:	data_out=16'h3a3;
17'h10961:	data_out=16'h21a;
17'h10962:	data_out=16'h24;
17'h10963:	data_out=16'h44c;
17'h10964:	data_out=16'h614;
17'h10965:	data_out=16'h278;
17'h10966:	data_out=16'h16;
17'h10967:	data_out=16'h628;
17'h10968:	data_out=16'hb9;
17'h10969:	data_out=16'hb3;
17'h1096a:	data_out=16'h7d;
17'h1096b:	data_out=16'h47a;
17'h1096c:	data_out=16'h69e;
17'h1096d:	data_out=16'h477;
17'h1096e:	data_out=16'h7b;
17'h1096f:	data_out=16'h42b;
17'h10970:	data_out=16'h9b;
17'h10971:	data_out=16'h71;
17'h10972:	data_out=16'h502;
17'h10973:	data_out=16'h534;
17'h10974:	data_out=16'h2b;
17'h10975:	data_out=16'h84f6;
17'h10976:	data_out=16'h3f1;
17'h10977:	data_out=16'h5f7;
17'h10978:	data_out=16'h20d;
17'h10979:	data_out=16'h41b;
17'h1097a:	data_out=16'h3ca;
17'h1097b:	data_out=16'hcc;
17'h1097c:	data_out=16'ha1;
17'h1097d:	data_out=16'hf;
17'h1097e:	data_out=16'h876;
17'h1097f:	data_out=16'h41c;
17'h10980:	data_out=16'h1a5;
17'h10981:	data_out=16'h9b;
17'h10982:	data_out=16'h824d;
17'h10983:	data_out=16'hc4;
17'h10984:	data_out=16'h8047;
17'h10985:	data_out=16'he0;
17'h10986:	data_out=16'h8015;
17'h10987:	data_out=16'h80bc;
17'h10988:	data_out=16'h81ae;
17'h10989:	data_out=16'h804e;
17'h1098a:	data_out=16'hb;
17'h1098b:	data_out=16'h8113;
17'h1098c:	data_out=16'h82a7;
17'h1098d:	data_out=16'hcb;
17'h1098e:	data_out=16'h8041;
17'h1098f:	data_out=16'h80d0;
17'h10990:	data_out=16'h8090;
17'h10991:	data_out=16'h8038;
17'h10992:	data_out=16'h810b;
17'h10993:	data_out=16'he8;
17'h10994:	data_out=16'hdf;
17'h10995:	data_out=16'h178;
17'h10996:	data_out=16'h1ba;
17'h10997:	data_out=16'h67;
17'h10998:	data_out=16'h807e;
17'h10999:	data_out=16'h80f1;
17'h1099a:	data_out=16'h28;
17'h1099b:	data_out=16'h8048;
17'h1099c:	data_out=16'h1de;
17'h1099d:	data_out=16'h8057;
17'h1099e:	data_out=16'hb2;
17'h1099f:	data_out=16'h800f;
17'h109a0:	data_out=16'h1c6;
17'h109a1:	data_out=16'h803d;
17'h109a2:	data_out=16'h8060;
17'h109a3:	data_out=16'h823e;
17'h109a4:	data_out=16'h823c;
17'h109a5:	data_out=16'h8107;
17'h109a6:	data_out=16'h818d;
17'h109a7:	data_out=16'h808b;
17'h109a8:	data_out=16'h8044;
17'h109a9:	data_out=16'hde;
17'h109aa:	data_out=16'h81e4;
17'h109ab:	data_out=16'h8032;
17'h109ac:	data_out=16'h105;
17'h109ad:	data_out=16'h8164;
17'h109ae:	data_out=16'h81d1;
17'h109af:	data_out=16'he8;
17'h109b0:	data_out=16'h4c;
17'h109b1:	data_out=16'h195;
17'h109b2:	data_out=16'h66;
17'h109b3:	data_out=16'h115;
17'h109b4:	data_out=16'ha7;
17'h109b5:	data_out=16'h8181;
17'h109b6:	data_out=16'h817b;
17'h109b7:	data_out=16'h8205;
17'h109b8:	data_out=16'h16b;
17'h109b9:	data_out=16'h140;
17'h109ba:	data_out=16'h80bf;
17'h109bb:	data_out=16'h8010;
17'h109bc:	data_out=16'h81ad;
17'h109bd:	data_out=16'h1e3;
17'h109be:	data_out=16'h804b;
17'h109bf:	data_out=16'hbf;
17'h109c0:	data_out=16'h80bc;
17'h109c1:	data_out=16'h8152;
17'h109c2:	data_out=16'h81b6;
17'h109c3:	data_out=16'h8005;
17'h109c4:	data_out=16'h8c;
17'h109c5:	data_out=16'h17a;
17'h109c6:	data_out=16'h8224;
17'h109c7:	data_out=16'h8103;
17'h109c8:	data_out=16'h8141;
17'h109c9:	data_out=16'h80eb;
17'h109ca:	data_out=16'h8190;
17'h109cb:	data_out=16'h827f;
17'h109cc:	data_out=16'h819d;
17'h109cd:	data_out=16'h24;
17'h109ce:	data_out=16'h8175;
17'h109cf:	data_out=16'h8162;
17'h109d0:	data_out=16'h1b;
17'h109d1:	data_out=16'hd7;
17'h109d2:	data_out=16'h8189;
17'h109d3:	data_out=16'h806c;
17'h109d4:	data_out=16'hc2;
17'h109d5:	data_out=16'h8106;
17'h109d6:	data_out=16'h807e;
17'h109d7:	data_out=16'h80e2;
17'h109d8:	data_out=16'h81ca;
17'h109d9:	data_out=16'h808c;
17'h109da:	data_out=16'h81a7;
17'h109db:	data_out=16'hd2;
17'h109dc:	data_out=16'h73;
17'h109dd:	data_out=16'h8036;
17'h109de:	data_out=16'hb2;
17'h109df:	data_out=16'h8006;
17'h109e0:	data_out=16'h81bd;
17'h109e1:	data_out=16'hff;
17'h109e2:	data_out=16'h807c;
17'h109e3:	data_out=16'heb;
17'h109e4:	data_out=16'hed;
17'h109e5:	data_out=16'h80ba;
17'h109e6:	data_out=16'h80d5;
17'h109e7:	data_out=16'h80df;
17'h109e8:	data_out=16'h8046;
17'h109e9:	data_out=16'h81fd;
17'h109ea:	data_out=16'h8050;
17'h109eb:	data_out=16'h16b;
17'h109ec:	data_out=16'h67;
17'h109ed:	data_out=16'h118;
17'h109ee:	data_out=16'h8041;
17'h109ef:	data_out=16'h13c;
17'h109f0:	data_out=16'h8049;
17'h109f1:	data_out=16'h816d;
17'h109f2:	data_out=16'h1c6;
17'h109f3:	data_out=16'h1a7;
17'h109f4:	data_out=16'h42;
17'h109f5:	data_out=16'h809b;
17'h109f6:	data_out=16'h8051;
17'h109f7:	data_out=16'h8102;
17'h109f8:	data_out=16'had;
17'h109f9:	data_out=16'h8204;
17'h109fa:	data_out=16'hdb;
17'h109fb:	data_out=16'h804a;
17'h109fc:	data_out=16'h8039;
17'h109fd:	data_out=16'h87;
17'h109fe:	data_out=16'h8046;
17'h109ff:	data_out=16'h800c;
17'h10a00:	data_out=16'h8003;
17'h10a01:	data_out=16'h5;
17'h10a02:	data_out=16'h1;
17'h10a03:	data_out=16'h5;
17'h10a04:	data_out=16'h7;
17'h10a05:	data_out=16'h9;
17'h10a06:	data_out=16'h4;
17'h10a07:	data_out=16'h8003;
17'h10a08:	data_out=16'h0;
17'h10a09:	data_out=16'h6;
17'h10a0a:	data_out=16'h8003;
17'h10a0b:	data_out=16'hc;
17'h10a0c:	data_out=16'h8004;
17'h10a0d:	data_out=16'h8005;
17'h10a0e:	data_out=16'h1;
17'h10a0f:	data_out=16'h2;
17'h10a10:	data_out=16'h8;
17'h10a11:	data_out=16'h9;
17'h10a12:	data_out=16'h8002;
17'h10a13:	data_out=16'h8003;
17'h10a14:	data_out=16'hc;
17'h10a15:	data_out=16'ha;
17'h10a16:	data_out=16'ha;
17'h10a17:	data_out=16'h6;
17'h10a18:	data_out=16'h8;
17'h10a19:	data_out=16'h6;
17'h10a1a:	data_out=16'h7;
17'h10a1b:	data_out=16'h8005;
17'h10a1c:	data_out=16'h5;
17'h10a1d:	data_out=16'hc;
17'h10a1e:	data_out=16'h8005;
17'h10a1f:	data_out=16'hb;
17'h10a20:	data_out=16'h6;
17'h10a21:	data_out=16'h8001;
17'h10a22:	data_out=16'h3;
17'h10a23:	data_out=16'h0;
17'h10a24:	data_out=16'h8003;
17'h10a25:	data_out=16'h8004;
17'h10a26:	data_out=16'h5;
17'h10a27:	data_out=16'h6;
17'h10a28:	data_out=16'h7;
17'h10a29:	data_out=16'h9;
17'h10a2a:	data_out=16'h7;
17'h10a2b:	data_out=16'h8;
17'h10a2c:	data_out=16'ha;
17'h10a2d:	data_out=16'h8004;
17'h10a2e:	data_out=16'h2;
17'h10a2f:	data_out=16'h5;
17'h10a30:	data_out=16'h8007;
17'h10a31:	data_out=16'h2;
17'h10a32:	data_out=16'h8;
17'h10a33:	data_out=16'hc;
17'h10a34:	data_out=16'h1;
17'h10a35:	data_out=16'h8;
17'h10a36:	data_out=16'h5;
17'h10a37:	data_out=16'h0;
17'h10a38:	data_out=16'h1;
17'h10a39:	data_out=16'h8001;
17'h10a3a:	data_out=16'h1;
17'h10a3b:	data_out=16'h8002;
17'h10a3c:	data_out=16'h8001;
17'h10a3d:	data_out=16'h0;
17'h10a3e:	data_out=16'h8004;
17'h10a3f:	data_out=16'hb;
17'h10a40:	data_out=16'h9;
17'h10a41:	data_out=16'h7;
17'h10a42:	data_out=16'h2;
17'h10a43:	data_out=16'h8005;
17'h10a44:	data_out=16'h9;
17'h10a45:	data_out=16'h8007;
17'h10a46:	data_out=16'h7;
17'h10a47:	data_out=16'h7;
17'h10a48:	data_out=16'ha;
17'h10a49:	data_out=16'h1;
17'h10a4a:	data_out=16'h5;
17'h10a4b:	data_out=16'h7;
17'h10a4c:	data_out=16'h5;
17'h10a4d:	data_out=16'ha;
17'h10a4e:	data_out=16'h1;
17'h10a4f:	data_out=16'h5;
17'h10a50:	data_out=16'h2;
17'h10a51:	data_out=16'h8004;
17'h10a52:	data_out=16'h1;
17'h10a53:	data_out=16'hb;
17'h10a54:	data_out=16'ha;
17'h10a55:	data_out=16'h8004;
17'h10a56:	data_out=16'h8001;
17'h10a57:	data_out=16'h2;
17'h10a58:	data_out=16'h1;
17'h10a59:	data_out=16'h5;
17'h10a5a:	data_out=16'h7;
17'h10a5b:	data_out=16'h4;
17'h10a5c:	data_out=16'h8007;
17'h10a5d:	data_out=16'hb;
17'h10a5e:	data_out=16'h5;
17'h10a5f:	data_out=16'h8;
17'h10a60:	data_out=16'h5;
17'h10a61:	data_out=16'h8006;
17'h10a62:	data_out=16'ha;
17'h10a63:	data_out=16'h3;
17'h10a64:	data_out=16'h8006;
17'h10a65:	data_out=16'h6;
17'h10a66:	data_out=16'h8007;
17'h10a67:	data_out=16'ha;
17'h10a68:	data_out=16'h8007;
17'h10a69:	data_out=16'h6;
17'h10a6a:	data_out=16'h1;
17'h10a6b:	data_out=16'h4;
17'h10a6c:	data_out=16'h4;
17'h10a6d:	data_out=16'ha;
17'h10a6e:	data_out=16'h8005;
17'h10a6f:	data_out=16'hb;
17'h10a70:	data_out=16'h9;
17'h10a71:	data_out=16'h8;
17'h10a72:	data_out=16'h9;
17'h10a73:	data_out=16'h8;
17'h10a74:	data_out=16'h7;
17'h10a75:	data_out=16'h8006;
17'h10a76:	data_out=16'h8002;
17'h10a77:	data_out=16'h8002;
17'h10a78:	data_out=16'h5;
17'h10a79:	data_out=16'he;
17'h10a7a:	data_out=16'h9;
17'h10a7b:	data_out=16'h5;
17'h10a7c:	data_out=16'h9;
17'h10a7d:	data_out=16'h0;
17'h10a7e:	data_out=16'h3;
17'h10a7f:	data_out=16'h4;
17'h10a80:	data_out=16'h116;
17'h10a81:	data_out=16'h12d;
17'h10a82:	data_out=16'ha2;
17'h10a83:	data_out=16'h8035;
17'h10a84:	data_out=16'h80a7;
17'h10a85:	data_out=16'h80eb;
17'h10a86:	data_out=16'h8156;
17'h10a87:	data_out=16'h802c;
17'h10a88:	data_out=16'hdd;
17'h10a89:	data_out=16'ha;
17'h10a8a:	data_out=16'h1a3;
17'h10a8b:	data_out=16'h24;
17'h10a8c:	data_out=16'hec;
17'h10a8d:	data_out=16'h806f;
17'h10a8e:	data_out=16'h8047;
17'h10a8f:	data_out=16'h8061;
17'h10a90:	data_out=16'h79;
17'h10a91:	data_out=16'h8023;
17'h10a92:	data_out=16'h89;
17'h10a93:	data_out=16'h805d;
17'h10a94:	data_out=16'h62;
17'h10a95:	data_out=16'h8085;
17'h10a96:	data_out=16'h8066;
17'h10a97:	data_out=16'ha4;
17'h10a98:	data_out=16'h803b;
17'h10a99:	data_out=16'h24;
17'h10a9a:	data_out=16'h80b8;
17'h10a9b:	data_out=16'hb9;
17'h10a9c:	data_out=16'h80dc;
17'h10a9d:	data_out=16'h1d2;
17'h10a9e:	data_out=16'h6e;
17'h10a9f:	data_out=16'h8164;
17'h10aa0:	data_out=16'hf8;
17'h10aa1:	data_out=16'h8036;
17'h10aa2:	data_out=16'hab;
17'h10aa3:	data_out=16'h12;
17'h10aa4:	data_out=16'h13;
17'h10aa5:	data_out=16'haf;
17'h10aa6:	data_out=16'ha4;
17'h10aa7:	data_out=16'h19c;
17'h10aa8:	data_out=16'h8038;
17'h10aa9:	data_out=16'h5c;
17'h10aaa:	data_out=16'hb2;
17'h10aab:	data_out=16'h137;
17'h10aac:	data_out=16'h802f;
17'h10aad:	data_out=16'h1a8;
17'h10aae:	data_out=16'h64;
17'h10aaf:	data_out=16'hcf;
17'h10ab0:	data_out=16'h8097;
17'h10ab1:	data_out=16'h162;
17'h10ab2:	data_out=16'h809e;
17'h10ab3:	data_out=16'h65;
17'h10ab4:	data_out=16'h9b;
17'h10ab5:	data_out=16'h25;
17'h10ab6:	data_out=16'hd7;
17'h10ab7:	data_out=16'h93;
17'h10ab8:	data_out=16'h8115;
17'h10ab9:	data_out=16'h8035;
17'h10aba:	data_out=16'h12d;
17'h10abb:	data_out=16'h5a;
17'h10abc:	data_out=16'h12e;
17'h10abd:	data_out=16'h8092;
17'h10abe:	data_out=16'h8044;
17'h10abf:	data_out=16'h811a;
17'h10ac0:	data_out=16'h80eb;
17'h10ac1:	data_out=16'h4e;
17'h10ac2:	data_out=16'h1a7;
17'h10ac3:	data_out=16'h8190;
17'h10ac4:	data_out=16'h8028;
17'h10ac5:	data_out=16'h8099;
17'h10ac6:	data_out=16'h17c;
17'h10ac7:	data_out=16'h22;
17'h10ac8:	data_out=16'h33;
17'h10ac9:	data_out=16'h81;
17'h10aca:	data_out=16'h8043;
17'h10acb:	data_out=16'h1fa;
17'h10acc:	data_out=16'h83;
17'h10acd:	data_out=16'hb7;
17'h10ace:	data_out=16'hb7;
17'h10acf:	data_out=16'h60;
17'h10ad0:	data_out=16'h8107;
17'h10ad1:	data_out=16'h8168;
17'h10ad2:	data_out=16'h802f;
17'h10ad3:	data_out=16'h1ea;
17'h10ad4:	data_out=16'hc7;
17'h10ad5:	data_out=16'h8023;
17'h10ad6:	data_out=16'h802b;
17'h10ad7:	data_out=16'h806b;
17'h10ad8:	data_out=16'h6b;
17'h10ad9:	data_out=16'h80d4;
17'h10ada:	data_out=16'hf0;
17'h10adb:	data_out=16'h815e;
17'h10adc:	data_out=16'h9d;
17'h10add:	data_out=16'h8c;
17'h10ade:	data_out=16'hdb;
17'h10adf:	data_out=16'h7c;
17'h10ae0:	data_out=16'he2;
17'h10ae1:	data_out=16'h8107;
17'h10ae2:	data_out=16'h8017;
17'h10ae3:	data_out=16'h5c;
17'h10ae4:	data_out=16'h4e;
17'h10ae5:	data_out=16'h6c;
17'h10ae6:	data_out=16'h1e;
17'h10ae7:	data_out=16'h8001;
17'h10ae8:	data_out=16'h8036;
17'h10ae9:	data_out=16'hf7;
17'h10aea:	data_out=16'h8043;
17'h10aeb:	data_out=16'h8106;
17'h10aec:	data_out=16'h348;
17'h10aed:	data_out=16'h6d;
17'h10aee:	data_out=16'h8041;
17'h10aef:	data_out=16'h8056;
17'h10af0:	data_out=16'h8046;
17'h10af1:	data_out=16'h807c;
17'h10af2:	data_out=16'h8138;
17'h10af3:	data_out=16'h8122;
17'h10af4:	data_out=16'h8099;
17'h10af5:	data_out=16'h8131;
17'h10af6:	data_out=16'h83;
17'h10af7:	data_out=16'h8143;
17'h10af8:	data_out=16'h8158;
17'h10af9:	data_out=16'h44;
17'h10afa:	data_out=16'h69;
17'h10afb:	data_out=16'h803c;
17'h10afc:	data_out=16'h8030;
17'h10afd:	data_out=16'h81ad;
17'h10afe:	data_out=16'h802f;
17'h10aff:	data_out=16'h812f;
17'h10b00:	data_out=16'h8579;
17'h10b01:	data_out=16'h1eb;
17'h10b02:	data_out=16'h77e;
17'h10b03:	data_out=16'h8038;
17'h10b04:	data_out=16'h81b9;
17'h10b05:	data_out=16'h45e;
17'h10b06:	data_out=16'h1b2;
17'h10b07:	data_out=16'h365;
17'h10b08:	data_out=16'h957;
17'h10b09:	data_out=16'h8115;
17'h10b0a:	data_out=16'h830a;
17'h10b0b:	data_out=16'h42c;
17'h10b0c:	data_out=16'h76b;
17'h10b0d:	data_out=16'h258;
17'h10b0e:	data_out=16'h18d;
17'h10b0f:	data_out=16'h966;
17'h10b10:	data_out=16'h8014;
17'h10b11:	data_out=16'hd7;
17'h10b12:	data_out=16'h540;
17'h10b13:	data_out=16'h806d;
17'h10b14:	data_out=16'h30d;
17'h10b15:	data_out=16'h8095;
17'h10b16:	data_out=16'hfa;
17'h10b17:	data_out=16'h223;
17'h10b18:	data_out=16'h220;
17'h10b19:	data_out=16'h8055;
17'h10b1a:	data_out=16'h8172;
17'h10b1b:	data_out=16'h4ed;
17'h10b1c:	data_out=16'h346;
17'h10b1d:	data_out=16'h2c1;
17'h10b1e:	data_out=16'h585;
17'h10b1f:	data_out=16'h657;
17'h10b20:	data_out=16'h431;
17'h10b21:	data_out=16'h19f;
17'h10b22:	data_out=16'h8312;
17'h10b23:	data_out=16'h1c4;
17'h10b24:	data_out=16'h1c6;
17'h10b25:	data_out=16'h81e7;
17'h10b26:	data_out=16'h211;
17'h10b27:	data_out=16'h467;
17'h10b28:	data_out=16'h1ed;
17'h10b29:	data_out=16'h801f;
17'h10b2a:	data_out=16'h6d1;
17'h10b2b:	data_out=16'h3e0;
17'h10b2c:	data_out=16'h33;
17'h10b2d:	data_out=16'h8891;
17'h10b2e:	data_out=16'h7f3;
17'h10b2f:	data_out=16'h41d;
17'h10b30:	data_out=16'h8105;
17'h10b31:	data_out=16'h9;
17'h10b32:	data_out=16'h8157;
17'h10b33:	data_out=16'h454;
17'h10b34:	data_out=16'h13b;
17'h10b35:	data_out=16'h68c;
17'h10b36:	data_out=16'h97d;
17'h10b37:	data_out=16'h6f2;
17'h10b38:	data_out=16'h5d;
17'h10b39:	data_out=16'h548;
17'h10b3a:	data_out=16'h8054;
17'h10b3b:	data_out=16'h9f;
17'h10b3c:	data_out=16'h463;
17'h10b3d:	data_out=16'h8286;
17'h10b3e:	data_out=16'h1fc;
17'h10b3f:	data_out=16'h45b;
17'h10b40:	data_out=16'hb7;
17'h10b41:	data_out=16'h960;
17'h10b42:	data_out=16'h8496;
17'h10b43:	data_out=16'h1d9;
17'h10b44:	data_out=16'h803e;
17'h10b45:	data_out=16'h8088;
17'h10b46:	data_out=16'h1f7;
17'h10b47:	data_out=16'hdc;
17'h10b48:	data_out=16'h451;
17'h10b49:	data_out=16'h8227;
17'h10b4a:	data_out=16'h725;
17'h10b4b:	data_out=16'h2bc;
17'h10b4c:	data_out=16'hff;
17'h10b4d:	data_out=16'h831f;
17'h10b4e:	data_out=16'h834;
17'h10b4f:	data_out=16'h117;
17'h10b50:	data_out=16'h27f;
17'h10b51:	data_out=16'h612;
17'h10b52:	data_out=16'h6b;
17'h10b53:	data_out=16'h6d3;
17'h10b54:	data_out=16'h3a8;
17'h10b55:	data_out=16'h7e0;
17'h10b56:	data_out=16'h2cf;
17'h10b57:	data_out=16'h141;
17'h10b58:	data_out=16'h890;
17'h10b59:	data_out=16'hf8;
17'h10b5a:	data_out=16'h117;
17'h10b5b:	data_out=16'h53c;
17'h10b5c:	data_out=16'h444;
17'h10b5d:	data_out=16'h1ae;
17'h10b5e:	data_out=16'h39f;
17'h10b5f:	data_out=16'h1e4;
17'h10b60:	data_out=16'h8080;
17'h10b61:	data_out=16'h274;
17'h10b62:	data_out=16'h473;
17'h10b63:	data_out=16'h4a3;
17'h10b64:	data_out=16'h6f;
17'h10b65:	data_out=16'h8022;
17'h10b66:	data_out=16'h8014;
17'h10b67:	data_out=16'h33c;
17'h10b68:	data_out=16'h1b2;
17'h10b69:	data_out=16'h8f7;
17'h10b6a:	data_out=16'h162;
17'h10b6b:	data_out=16'h7b;
17'h10b6c:	data_out=16'h84f7;
17'h10b6d:	data_out=16'h48e;
17'h10b6e:	data_out=16'h16b;
17'h10b6f:	data_out=16'h8215;
17'h10b70:	data_out=16'h17b;
17'h10b71:	data_out=16'h99e;
17'h10b72:	data_out=16'h8357;
17'h10b73:	data_out=16'h80b6;
17'h10b74:	data_out=16'h80f5;
17'h10b75:	data_out=16'h3c5;
17'h10b76:	data_out=16'h276;
17'h10b77:	data_out=16'hd3;
17'h10b78:	data_out=16'h117;
17'h10b79:	data_out=16'ha00;
17'h10b7a:	data_out=16'h3c1;
17'h10b7b:	data_out=16'h1f5;
17'h10b7c:	data_out=16'h2fb;
17'h10b7d:	data_out=16'h4d1;
17'h10b7e:	data_out=16'h8119;
17'h10b7f:	data_out=16'h1ca;
17'h10b80:	data_out=16'h8a00;
17'h10b81:	data_out=16'h8416;
17'h10b82:	data_out=16'h9f6;
17'h10b83:	data_out=16'h1;
17'h10b84:	data_out=16'h9b0;
17'h10b85:	data_out=16'h9fa;
17'h10b86:	data_out=16'h9ff;
17'h10b87:	data_out=16'h89fb;
17'h10b88:	data_out=16'h826a;
17'h10b89:	data_out=16'h89fb;
17'h10b8a:	data_out=16'h8a00;
17'h10b8b:	data_out=16'h9b3;
17'h10b8c:	data_out=16'h8a00;
17'h10b8d:	data_out=16'h799;
17'h10b8e:	data_out=16'h353;
17'h10b8f:	data_out=16'h9f1;
17'h10b90:	data_out=16'h89f1;
17'h10b91:	data_out=16'ha00;
17'h10b92:	data_out=16'h9ff;
17'h10b93:	data_out=16'h207;
17'h10b94:	data_out=16'ha00;
17'h10b95:	data_out=16'h83dc;
17'h10b96:	data_out=16'h8a00;
17'h10b97:	data_out=16'h9ff;
17'h10b98:	data_out=16'h2cc;
17'h10b99:	data_out=16'ha00;
17'h10b9a:	data_out=16'ha00;
17'h10b9b:	data_out=16'ha00;
17'h10b9c:	data_out=16'h9fa;
17'h10b9d:	data_out=16'h884;
17'h10b9e:	data_out=16'h9fc;
17'h10b9f:	data_out=16'ha00;
17'h10ba0:	data_out=16'ha00;
17'h10ba1:	data_out=16'h3c5;
17'h10ba2:	data_out=16'h89f9;
17'h10ba3:	data_out=16'h8a00;
17'h10ba4:	data_out=16'h8a00;
17'h10ba5:	data_out=16'h89fb;
17'h10ba6:	data_out=16'h8a00;
17'h10ba7:	data_out=16'ha00;
17'h10ba8:	data_out=16'h4f1;
17'h10ba9:	data_out=16'h89ff;
17'h10baa:	data_out=16'h89fd;
17'h10bab:	data_out=16'ha00;
17'h10bac:	data_out=16'h8a00;
17'h10bad:	data_out=16'h8a00;
17'h10bae:	data_out=16'ha00;
17'h10baf:	data_out=16'ha00;
17'h10bb0:	data_out=16'h8a00;
17'h10bb1:	data_out=16'h652;
17'h10bb2:	data_out=16'h89e8;
17'h10bb3:	data_out=16'ha00;
17'h10bb4:	data_out=16'h8a00;
17'h10bb5:	data_out=16'h9d0;
17'h10bb6:	data_out=16'h64c;
17'h10bb7:	data_out=16'h9f7;
17'h10bb8:	data_out=16'ha00;
17'h10bb9:	data_out=16'ha00;
17'h10bba:	data_out=16'h89f9;
17'h10bbb:	data_out=16'h8454;
17'h10bbc:	data_out=16'h9ff;
17'h10bbd:	data_out=16'h622;
17'h10bbe:	data_out=16'h52a;
17'h10bbf:	data_out=16'h9fa;
17'h10bc0:	data_out=16'h87e0;
17'h10bc1:	data_out=16'h9fa;
17'h10bc2:	data_out=16'h8a00;
17'h10bc3:	data_out=16'h9fe;
17'h10bc4:	data_out=16'ha00;
17'h10bc5:	data_out=16'h847b;
17'h10bc6:	data_out=16'h8a00;
17'h10bc7:	data_out=16'h89ff;
17'h10bc8:	data_out=16'ha00;
17'h10bc9:	data_out=16'h89fe;
17'h10bca:	data_out=16'h551;
17'h10bcb:	data_out=16'h8a00;
17'h10bcc:	data_out=16'h8a00;
17'h10bcd:	data_out=16'h89fb;
17'h10bce:	data_out=16'h5b8;
17'h10bcf:	data_out=16'h8a00;
17'h10bd0:	data_out=16'h836c;
17'h10bd1:	data_out=16'h9f4;
17'h10bd2:	data_out=16'h8a00;
17'h10bd3:	data_out=16'ha00;
17'h10bd4:	data_out=16'ha00;
17'h10bd5:	data_out=16'h9f7;
17'h10bd6:	data_out=16'h89ed;
17'h10bd7:	data_out=16'h89e1;
17'h10bd8:	data_out=16'h9fd;
17'h10bd9:	data_out=16'h89f5;
17'h10bda:	data_out=16'ha00;
17'h10bdb:	data_out=16'ha00;
17'h10bdc:	data_out=16'ha00;
17'h10bdd:	data_out=16'h89fd;
17'h10bde:	data_out=16'ha00;
17'h10bdf:	data_out=16'h80cc;
17'h10be0:	data_out=16'h8a00;
17'h10be1:	data_out=16'h9f9;
17'h10be2:	data_out=16'h92c;
17'h10be3:	data_out=16'ha00;
17'h10be4:	data_out=16'h16e;
17'h10be5:	data_out=16'h9d8;
17'h10be6:	data_out=16'ha00;
17'h10be7:	data_out=16'h84f6;
17'h10be8:	data_out=16'h41f;
17'h10be9:	data_out=16'h8875;
17'h10bea:	data_out=16'h311;
17'h10beb:	data_out=16'h9ff;
17'h10bec:	data_out=16'h8a00;
17'h10bed:	data_out=16'ha00;
17'h10bee:	data_out=16'h312;
17'h10bef:	data_out=16'h8288;
17'h10bf0:	data_out=16'h337;
17'h10bf1:	data_out=16'h9fb;
17'h10bf2:	data_out=16'h84f2;
17'h10bf3:	data_out=16'h7cc;
17'h10bf4:	data_out=16'h8a00;
17'h10bf5:	data_out=16'h9f7;
17'h10bf6:	data_out=16'ha00;
17'h10bf7:	data_out=16'h89fc;
17'h10bf8:	data_out=16'h9fc;
17'h10bf9:	data_out=16'h7f0;
17'h10bfa:	data_out=16'ha00;
17'h10bfb:	data_out=16'h574;
17'h10bfc:	data_out=16'h811;
17'h10bfd:	data_out=16'ha00;
17'h10bfe:	data_out=16'h89e5;
17'h10bff:	data_out=16'h8867;
17'h10c00:	data_out=16'h89c2;
17'h10c01:	data_out=16'h9ed;
17'h10c02:	data_out=16'h9d3;
17'h10c03:	data_out=16'h8a00;
17'h10c04:	data_out=16'ha00;
17'h10c05:	data_out=16'h9e0;
17'h10c06:	data_out=16'h5ef;
17'h10c07:	data_out=16'h876b;
17'h10c08:	data_out=16'h9f9;
17'h10c09:	data_out=16'h89fb;
17'h10c0a:	data_out=16'h657;
17'h10c0b:	data_out=16'h6ce;
17'h10c0c:	data_out=16'h89fe;
17'h10c0d:	data_out=16'h8a00;
17'h10c0e:	data_out=16'h569;
17'h10c0f:	data_out=16'h3f6;
17'h10c10:	data_out=16'h89f8;
17'h10c11:	data_out=16'ha00;
17'h10c12:	data_out=16'h9eb;
17'h10c13:	data_out=16'h83eb;
17'h10c14:	data_out=16'h9dc;
17'h10c15:	data_out=16'h93d;
17'h10c16:	data_out=16'h8a00;
17'h10c17:	data_out=16'h41b;
17'h10c18:	data_out=16'h9ff;
17'h10c19:	data_out=16'ha00;
17'h10c1a:	data_out=16'h9e9;
17'h10c1b:	data_out=16'h9dd;
17'h10c1c:	data_out=16'h858;
17'h10c1d:	data_out=16'h9fe;
17'h10c1e:	data_out=16'h7de;
17'h10c1f:	data_out=16'h9f9;
17'h10c20:	data_out=16'h9fc;
17'h10c21:	data_out=16'h5d7;
17'h10c22:	data_out=16'h89fb;
17'h10c23:	data_out=16'h8546;
17'h10c24:	data_out=16'h852d;
17'h10c25:	data_out=16'h89fa;
17'h10c26:	data_out=16'h8a00;
17'h10c27:	data_out=16'ha00;
17'h10c28:	data_out=16'h913;
17'h10c29:	data_out=16'h8a00;
17'h10c2a:	data_out=16'h89fa;
17'h10c2b:	data_out=16'ha00;
17'h10c2c:	data_out=16'h89ff;
17'h10c2d:	data_out=16'h89fe;
17'h10c2e:	data_out=16'h614;
17'h10c2f:	data_out=16'h9e1;
17'h10c30:	data_out=16'h8a00;
17'h10c31:	data_out=16'h9fd;
17'h10c32:	data_out=16'h89fc;
17'h10c33:	data_out=16'h9f1;
17'h10c34:	data_out=16'h620;
17'h10c35:	data_out=16'h9fe;
17'h10c36:	data_out=16'h9ec;
17'h10c37:	data_out=16'h9d7;
17'h10c38:	data_out=16'h9f8;
17'h10c39:	data_out=16'h9ef;
17'h10c3a:	data_out=16'h89fa;
17'h10c3b:	data_out=16'h9fe;
17'h10c3c:	data_out=16'h7b8;
17'h10c3d:	data_out=16'h9d8;
17'h10c3e:	data_out=16'h921;
17'h10c3f:	data_out=16'h9e0;
17'h10c40:	data_out=16'h9e3;
17'h10c41:	data_out=16'h9ca;
17'h10c42:	data_out=16'h8a00;
17'h10c43:	data_out=16'h23;
17'h10c44:	data_out=16'ha00;
17'h10c45:	data_out=16'h8d0;
17'h10c46:	data_out=16'h8844;
17'h10c47:	data_out=16'h89f9;
17'h10c48:	data_out=16'h9ee;
17'h10c49:	data_out=16'h89fb;
17'h10c4a:	data_out=16'ha00;
17'h10c4b:	data_out=16'h8a00;
17'h10c4c:	data_out=16'h89fd;
17'h10c4d:	data_out=16'h89fa;
17'h10c4e:	data_out=16'h6e1;
17'h10c4f:	data_out=16'h89ff;
17'h10c50:	data_out=16'h89fd;
17'h10c51:	data_out=16'h6aa;
17'h10c52:	data_out=16'h8a00;
17'h10c53:	data_out=16'ha00;
17'h10c54:	data_out=16'h9ef;
17'h10c55:	data_out=16'hb0;
17'h10c56:	data_out=16'h6d8;
17'h10c57:	data_out=16'h8138;
17'h10c58:	data_out=16'h9d7;
17'h10c59:	data_out=16'h81fc;
17'h10c5a:	data_out=16'ha00;
17'h10c5b:	data_out=16'ha00;
17'h10c5c:	data_out=16'h9f0;
17'h10c5d:	data_out=16'h89fa;
17'h10c5e:	data_out=16'h9d8;
17'h10c5f:	data_out=16'h7e4;
17'h10c60:	data_out=16'h8a00;
17'h10c61:	data_out=16'h9e5;
17'h10c62:	data_out=16'h875c;
17'h10c63:	data_out=16'h9f1;
17'h10c64:	data_out=16'h9ff;
17'h10c65:	data_out=16'h9ff;
17'h10c66:	data_out=16'ha00;
17'h10c67:	data_out=16'h89d8;
17'h10c68:	data_out=16'h7ed;
17'h10c69:	data_out=16'h14;
17'h10c6a:	data_out=16'h511;
17'h10c6b:	data_out=16'h9de;
17'h10c6c:	data_out=16'h89fa;
17'h10c6d:	data_out=16'h9f1;
17'h10c6e:	data_out=16'h50f;
17'h10c6f:	data_out=16'h8a00;
17'h10c70:	data_out=16'h545;
17'h10c71:	data_out=16'h9d8;
17'h10c72:	data_out=16'h8055;
17'h10c73:	data_out=16'h4bf;
17'h10c74:	data_out=16'h8a00;
17'h10c75:	data_out=16'h9ce;
17'h10c76:	data_out=16'h9ff;
17'h10c77:	data_out=16'h89fb;
17'h10c78:	data_out=16'h8a00;
17'h10c79:	data_out=16'h7a;
17'h10c7a:	data_out=16'h9e8;
17'h10c7b:	data_out=16'h922;
17'h10c7c:	data_out=16'ha00;
17'h10c7d:	data_out=16'ha00;
17'h10c7e:	data_out=16'h89f4;
17'h10c7f:	data_out=16'h4a6;
17'h10c80:	data_out=16'h89f0;
17'h10c81:	data_out=16'h9f8;
17'h10c82:	data_out=16'h926;
17'h10c83:	data_out=16'h8a00;
17'h10c84:	data_out=16'h9e0;
17'h10c85:	data_out=16'h295;
17'h10c86:	data_out=16'h996;
17'h10c87:	data_out=16'h887;
17'h10c88:	data_out=16'ha00;
17'h10c89:	data_out=16'h89f9;
17'h10c8a:	data_out=16'h9ff;
17'h10c8b:	data_out=16'h9e0;
17'h10c8c:	data_out=16'h89f6;
17'h10c8d:	data_out=16'h8a00;
17'h10c8e:	data_out=16'h9fa;
17'h10c8f:	data_out=16'h89dc;
17'h10c90:	data_out=16'h89fd;
17'h10c91:	data_out=16'ha00;
17'h10c92:	data_out=16'h8d9;
17'h10c93:	data_out=16'h211;
17'h10c94:	data_out=16'h2d1;
17'h10c95:	data_out=16'hc5;
17'h10c96:	data_out=16'h8a00;
17'h10c97:	data_out=16'h8734;
17'h10c98:	data_out=16'h762;
17'h10c99:	data_out=16'ha00;
17'h10c9a:	data_out=16'h9b1;
17'h10c9b:	data_out=16'h96e;
17'h10c9c:	data_out=16'h863e;
17'h10c9d:	data_out=16'h9ff;
17'h10c9e:	data_out=16'h891c;
17'h10c9f:	data_out=16'ha00;
17'h10ca0:	data_out=16'h9c2;
17'h10ca1:	data_out=16'h9fa;
17'h10ca2:	data_out=16'h89ff;
17'h10ca3:	data_out=16'ha00;
17'h10ca4:	data_out=16'ha00;
17'h10ca5:	data_out=16'h89f7;
17'h10ca6:	data_out=16'h89e6;
17'h10ca7:	data_out=16'ha00;
17'h10ca8:	data_out=16'h9fa;
17'h10ca9:	data_out=16'h8a00;
17'h10caa:	data_out=16'h89fb;
17'h10cab:	data_out=16'ha00;
17'h10cac:	data_out=16'h8a00;
17'h10cad:	data_out=16'h89e3;
17'h10cae:	data_out=16'h488;
17'h10caf:	data_out=16'h8310;
17'h10cb0:	data_out=16'h81e;
17'h10cb1:	data_out=16'ha00;
17'h10cb2:	data_out=16'h9d1;
17'h10cb3:	data_out=16'h9e9;
17'h10cb4:	data_out=16'h93f;
17'h10cb5:	data_out=16'h9ff;
17'h10cb6:	data_out=16'h595;
17'h10cb7:	data_out=16'h9f0;
17'h10cb8:	data_out=16'h9df;
17'h10cb9:	data_out=16'h8aa;
17'h10cba:	data_out=16'h89f9;
17'h10cbb:	data_out=16'ha00;
17'h10cbc:	data_out=16'h9c2;
17'h10cbd:	data_out=16'h8746;
17'h10cbe:	data_out=16'h9fa;
17'h10cbf:	data_out=16'h235;
17'h10cc0:	data_out=16'h9b3;
17'h10cc1:	data_out=16'h80f7;
17'h10cc2:	data_out=16'h8a00;
17'h10cc3:	data_out=16'h89ff;
17'h10cc4:	data_out=16'ha00;
17'h10cc5:	data_out=16'h8020;
17'h10cc6:	data_out=16'h9bc;
17'h10cc7:	data_out=16'h89f7;
17'h10cc8:	data_out=16'h8e1;
17'h10cc9:	data_out=16'h89f7;
17'h10cca:	data_out=16'h9fd;
17'h10ccb:	data_out=16'h8a00;
17'h10ccc:	data_out=16'h89fd;
17'h10ccd:	data_out=16'h89ff;
17'h10cce:	data_out=16'ha00;
17'h10ccf:	data_out=16'h89fe;
17'h10cd0:	data_out=16'h8a00;
17'h10cd1:	data_out=16'h8686;
17'h10cd2:	data_out=16'h248;
17'h10cd3:	data_out=16'ha00;
17'h10cd4:	data_out=16'h9b8;
17'h10cd5:	data_out=16'h8733;
17'h10cd6:	data_out=16'h9e0;
17'h10cd7:	data_out=16'h9b8;
17'h10cd8:	data_out=16'h921;
17'h10cd9:	data_out=16'h65d;
17'h10cda:	data_out=16'ha00;
17'h10cdb:	data_out=16'ha00;
17'h10cdc:	data_out=16'h9f9;
17'h10cdd:	data_out=16'h89ff;
17'h10cde:	data_out=16'h89fa;
17'h10cdf:	data_out=16'h85fe;
17'h10ce0:	data_out=16'h89cc;
17'h10ce1:	data_out=16'h9d2;
17'h10ce2:	data_out=16'h89d3;
17'h10ce3:	data_out=16'h9ef;
17'h10ce4:	data_out=16'h9f9;
17'h10ce5:	data_out=16'h9ff;
17'h10ce6:	data_out=16'ha00;
17'h10ce7:	data_out=16'h89f5;
17'h10ce8:	data_out=16'h9fa;
17'h10ce9:	data_out=16'h744;
17'h10cea:	data_out=16'h9fa;
17'h10ceb:	data_out=16'h10a;
17'h10cec:	data_out=16'h89fa;
17'h10ced:	data_out=16'h9ee;
17'h10cee:	data_out=16'h9fa;
17'h10cef:	data_out=16'h8a00;
17'h10cf0:	data_out=16'h9fa;
17'h10cf1:	data_out=16'h830;
17'h10cf2:	data_out=16'h808a;
17'h10cf3:	data_out=16'h9c4;
17'h10cf4:	data_out=16'h7d1;
17'h10cf5:	data_out=16'h9ae;
17'h10cf6:	data_out=16'h9ec;
17'h10cf7:	data_out=16'h89fe;
17'h10cf8:	data_out=16'h8a00;
17'h10cf9:	data_out=16'h89d0;
17'h10cfa:	data_out=16'h8aa;
17'h10cfb:	data_out=16'h9fa;
17'h10cfc:	data_out=16'h9fd;
17'h10cfd:	data_out=16'h9e9;
17'h10cfe:	data_out=16'h8323;
17'h10cff:	data_out=16'h8a00;
17'h10d00:	data_out=16'h89ce;
17'h10d01:	data_out=16'h9fc;
17'h10d02:	data_out=16'h4eb;
17'h10d03:	data_out=16'h89f7;
17'h10d04:	data_out=16'h9ed;
17'h10d05:	data_out=16'h47d;
17'h10d06:	data_out=16'h9ec;
17'h10d07:	data_out=16'h8066;
17'h10d08:	data_out=16'h82f7;
17'h10d09:	data_out=16'h89f2;
17'h10d0a:	data_out=16'ha00;
17'h10d0b:	data_out=16'h9ff;
17'h10d0c:	data_out=16'h89e5;
17'h10d0d:	data_out=16'h8a00;
17'h10d0e:	data_out=16'h9f6;
17'h10d0f:	data_out=16'h89a4;
17'h10d10:	data_out=16'h89fa;
17'h10d11:	data_out=16'ha00;
17'h10d12:	data_out=16'h821f;
17'h10d13:	data_out=16'ha00;
17'h10d14:	data_out=16'h89ba;
17'h10d15:	data_out=16'hef;
17'h10d16:	data_out=16'h89fb;
17'h10d17:	data_out=16'h89e0;
17'h10d18:	data_out=16'h89eb;
17'h10d19:	data_out=16'h9fb;
17'h10d1a:	data_out=16'h9a3;
17'h10d1b:	data_out=16'h8969;
17'h10d1c:	data_out=16'h89fa;
17'h10d1d:	data_out=16'ha00;
17'h10d1e:	data_out=16'h89c6;
17'h10d1f:	data_out=16'ha00;
17'h10d20:	data_out=16'h9c2;
17'h10d21:	data_out=16'h9f6;
17'h10d22:	data_out=16'h89fb;
17'h10d23:	data_out=16'h9ff;
17'h10d24:	data_out=16'h9ff;
17'h10d25:	data_out=16'h89d9;
17'h10d26:	data_out=16'h8990;
17'h10d27:	data_out=16'ha00;
17'h10d28:	data_out=16'h9f6;
17'h10d29:	data_out=16'h8a00;
17'h10d2a:	data_out=16'h899f;
17'h10d2b:	data_out=16'h9fe;
17'h10d2c:	data_out=16'h89fb;
17'h10d2d:	data_out=16'h8656;
17'h10d2e:	data_out=16'h83ea;
17'h10d2f:	data_out=16'h89d2;
17'h10d30:	data_out=16'h9da;
17'h10d31:	data_out=16'ha00;
17'h10d32:	data_out=16'h9d4;
17'h10d33:	data_out=16'h89c5;
17'h10d34:	data_out=16'ha00;
17'h10d35:	data_out=16'ha00;
17'h10d36:	data_out=16'h8936;
17'h10d37:	data_out=16'h9e5;
17'h10d38:	data_out=16'h9e9;
17'h10d39:	data_out=16'h89e1;
17'h10d3a:	data_out=16'h89f7;
17'h10d3b:	data_out=16'ha00;
17'h10d3c:	data_out=16'h9d1;
17'h10d3d:	data_out=16'h848d;
17'h10d3e:	data_out=16'h9f6;
17'h10d3f:	data_out=16'h436;
17'h10d40:	data_out=16'h9b5;
17'h10d41:	data_out=16'h89fe;
17'h10d42:	data_out=16'h8a00;
17'h10d43:	data_out=16'h89f9;
17'h10d44:	data_out=16'ha00;
17'h10d45:	data_out=16'h37;
17'h10d46:	data_out=16'h9c0;
17'h10d47:	data_out=16'h89d0;
17'h10d48:	data_out=16'h826d;
17'h10d49:	data_out=16'h89ee;
17'h10d4a:	data_out=16'h9d0;
17'h10d4b:	data_out=16'h89f0;
17'h10d4c:	data_out=16'h89fc;
17'h10d4d:	data_out=16'h89fe;
17'h10d4e:	data_out=16'h9f6;
17'h10d4f:	data_out=16'h89fd;
17'h10d50:	data_out=16'h89fc;
17'h10d51:	data_out=16'h89f7;
17'h10d52:	data_out=16'h945;
17'h10d53:	data_out=16'h9ff;
17'h10d54:	data_out=16'h6b2;
17'h10d55:	data_out=16'h8979;
17'h10d56:	data_out=16'h9d8;
17'h10d57:	data_out=16'h9a4;
17'h10d58:	data_out=16'h89fb;
17'h10d59:	data_out=16'h995;
17'h10d5a:	data_out=16'h9fa;
17'h10d5b:	data_out=16'ha00;
17'h10d5c:	data_out=16'h9e1;
17'h10d5d:	data_out=16'h89f8;
17'h10d5e:	data_out=16'h89d0;
17'h10d5f:	data_out=16'h89f1;
17'h10d60:	data_out=16'h89bc;
17'h10d61:	data_out=16'h9c9;
17'h10d62:	data_out=16'h8927;
17'h10d63:	data_out=16'h89a4;
17'h10d64:	data_out=16'ha00;
17'h10d65:	data_out=16'ha00;
17'h10d66:	data_out=16'h9ff;
17'h10d67:	data_out=16'h89f4;
17'h10d68:	data_out=16'h9f6;
17'h10d69:	data_out=16'h89be;
17'h10d6a:	data_out=16'h9f6;
17'h10d6b:	data_out=16'h3a5;
17'h10d6c:	data_out=16'h89f5;
17'h10d6d:	data_out=16'h89ad;
17'h10d6e:	data_out=16'h9f6;
17'h10d6f:	data_out=16'h8ac;
17'h10d70:	data_out=16'h9f6;
17'h10d71:	data_out=16'h8958;
17'h10d72:	data_out=16'h98a;
17'h10d73:	data_out=16'h9c9;
17'h10d74:	data_out=16'h9ca;
17'h10d75:	data_out=16'h941;
17'h10d76:	data_out=16'h330;
17'h10d77:	data_out=16'h89f9;
17'h10d78:	data_out=16'h8a00;
17'h10d79:	data_out=16'h89ff;
17'h10d7a:	data_out=16'h89a5;
17'h10d7b:	data_out=16'h9f6;
17'h10d7c:	data_out=16'h81bb;
17'h10d7d:	data_out=16'h9ee;
17'h10d7e:	data_out=16'h9f3;
17'h10d7f:	data_out=16'h8a00;
17'h10d80:	data_out=16'h89c3;
17'h10d81:	data_out=16'h9f6;
17'h10d82:	data_out=16'h8a00;
17'h10d83:	data_out=16'h89f7;
17'h10d84:	data_out=16'h9ec;
17'h10d85:	data_out=16'h59f;
17'h10d86:	data_out=16'h9f8;
17'h10d87:	data_out=16'h89fc;
17'h10d88:	data_out=16'h8a00;
17'h10d89:	data_out=16'h89d8;
17'h10d8a:	data_out=16'ha00;
17'h10d8b:	data_out=16'h860a;
17'h10d8c:	data_out=16'h8a00;
17'h10d8d:	data_out=16'h8a00;
17'h10d8e:	data_out=16'h9f9;
17'h10d8f:	data_out=16'h8a00;
17'h10d90:	data_out=16'h89f8;
17'h10d91:	data_out=16'ha00;
17'h10d92:	data_out=16'h8a00;
17'h10d93:	data_out=16'ha00;
17'h10d94:	data_out=16'h89d9;
17'h10d95:	data_out=16'h89fc;
17'h10d96:	data_out=16'h89fa;
17'h10d97:	data_out=16'h89d0;
17'h10d98:	data_out=16'h8a00;
17'h10d99:	data_out=16'h9eb;
17'h10d9a:	data_out=16'h9b1;
17'h10d9b:	data_out=16'h89e8;
17'h10d9c:	data_out=16'h89fd;
17'h10d9d:	data_out=16'ha00;
17'h10d9e:	data_out=16'h89f9;
17'h10d9f:	data_out=16'h8889;
17'h10da0:	data_out=16'h89b9;
17'h10da1:	data_out=16'h9f8;
17'h10da2:	data_out=16'h89f9;
17'h10da3:	data_out=16'h9f2;
17'h10da4:	data_out=16'h9f2;
17'h10da5:	data_out=16'h899c;
17'h10da6:	data_out=16'h89cc;
17'h10da7:	data_out=16'ha00;
17'h10da8:	data_out=16'h9f8;
17'h10da9:	data_out=16'h8a00;
17'h10daa:	data_out=16'h89fe;
17'h10dab:	data_out=16'h9fb;
17'h10dac:	data_out=16'h89fa;
17'h10dad:	data_out=16'ha00;
17'h10dae:	data_out=16'h8918;
17'h10daf:	data_out=16'h89f6;
17'h10db0:	data_out=16'h9db;
17'h10db1:	data_out=16'ha00;
17'h10db2:	data_out=16'h9cf;
17'h10db3:	data_out=16'h89e1;
17'h10db4:	data_out=16'ha00;
17'h10db5:	data_out=16'h9f0;
17'h10db6:	data_out=16'h89ff;
17'h10db7:	data_out=16'h89d2;
17'h10db8:	data_out=16'h9e9;
17'h10db9:	data_out=16'h89f4;
17'h10dba:	data_out=16'h89f5;
17'h10dbb:	data_out=16'h9f7;
17'h10dbc:	data_out=16'h679;
17'h10dbd:	data_out=16'h89c8;
17'h10dbe:	data_out=16'h9f8;
17'h10dbf:	data_out=16'h564;
17'h10dc0:	data_out=16'h9d1;
17'h10dc1:	data_out=16'h8a00;
17'h10dc2:	data_out=16'h89ff;
17'h10dc3:	data_out=16'h89f7;
17'h10dc4:	data_out=16'ha00;
17'h10dc5:	data_out=16'h89fc;
17'h10dc6:	data_out=16'h8771;
17'h10dc7:	data_out=16'h89f7;
17'h10dc8:	data_out=16'h897e;
17'h10dc9:	data_out=16'h8937;
17'h10dca:	data_out=16'h89e8;
17'h10dcb:	data_out=16'h89e9;
17'h10dcc:	data_out=16'h89fb;
17'h10dcd:	data_out=16'h89f9;
17'h10dce:	data_out=16'h89e9;
17'h10dcf:	data_out=16'h89eb;
17'h10dd0:	data_out=16'h89f7;
17'h10dd1:	data_out=16'h89ff;
17'h10dd2:	data_out=16'h9b5;
17'h10dd3:	data_out=16'h1e4;
17'h10dd4:	data_out=16'h89f5;
17'h10dd5:	data_out=16'h89f0;
17'h10dd6:	data_out=16'h9cd;
17'h10dd7:	data_out=16'h51e;
17'h10dd8:	data_out=16'h8a00;
17'h10dd9:	data_out=16'h9ba;
17'h10dda:	data_out=16'h85f4;
17'h10ddb:	data_out=16'ha00;
17'h10ddc:	data_out=16'h8135;
17'h10ddd:	data_out=16'h89f8;
17'h10dde:	data_out=16'h89f4;
17'h10ddf:	data_out=16'h89ff;
17'h10de0:	data_out=16'h89d8;
17'h10de1:	data_out=16'h9bf;
17'h10de2:	data_out=16'h8956;
17'h10de3:	data_out=16'h89d6;
17'h10de4:	data_out=16'ha00;
17'h10de5:	data_out=16'ha00;
17'h10de6:	data_out=16'h72d;
17'h10de7:	data_out=16'h89e1;
17'h10de8:	data_out=16'h9f8;
17'h10de9:	data_out=16'h8a00;
17'h10dea:	data_out=16'h9f9;
17'h10deb:	data_out=16'h8063;
17'h10dec:	data_out=16'h89d5;
17'h10ded:	data_out=16'h89da;
17'h10dee:	data_out=16'h9f9;
17'h10def:	data_out=16'h9c0;
17'h10df0:	data_out=16'h9f9;
17'h10df1:	data_out=16'h89f8;
17'h10df2:	data_out=16'h9b0;
17'h10df3:	data_out=16'h9e2;
17'h10df4:	data_out=16'h9b8;
17'h10df5:	data_out=16'h4f4;
17'h10df6:	data_out=16'h88ad;
17'h10df7:	data_out=16'h89ff;
17'h10df8:	data_out=16'h8a00;
17'h10df9:	data_out=16'h8a00;
17'h10dfa:	data_out=16'h89d9;
17'h10dfb:	data_out=16'h9f8;
17'h10dfc:	data_out=16'h8a00;
17'h10dfd:	data_out=16'h89e1;
17'h10dfe:	data_out=16'h97d;
17'h10dff:	data_out=16'h8a00;
17'h10e00:	data_out=16'h8936;
17'h10e01:	data_out=16'h9fb;
17'h10e02:	data_out=16'h8a00;
17'h10e03:	data_out=16'h89f6;
17'h10e04:	data_out=16'ha00;
17'h10e05:	data_out=16'h961;
17'h10e06:	data_out=16'h9fe;
17'h10e07:	data_out=16'h8a00;
17'h10e08:	data_out=16'h8a00;
17'h10e09:	data_out=16'h89aa;
17'h10e0a:	data_out=16'ha00;
17'h10e0b:	data_out=16'h8999;
17'h10e0c:	data_out=16'h8a00;
17'h10e0d:	data_out=16'h8a00;
17'h10e0e:	data_out=16'h979;
17'h10e0f:	data_out=16'h8a00;
17'h10e10:	data_out=16'h89d8;
17'h10e11:	data_out=16'ha00;
17'h10e12:	data_out=16'h8a00;
17'h10e13:	data_out=16'ha00;
17'h10e14:	data_out=16'h89da;
17'h10e15:	data_out=16'h89f4;
17'h10e16:	data_out=16'h89f7;
17'h10e17:	data_out=16'h89d5;
17'h10e18:	data_out=16'h8a00;
17'h10e19:	data_out=16'h9c5;
17'h10e1a:	data_out=16'h9df;
17'h10e1b:	data_out=16'h89e9;
17'h10e1c:	data_out=16'h89fa;
17'h10e1d:	data_out=16'ha00;
17'h10e1e:	data_out=16'h89fb;
17'h10e1f:	data_out=16'h8996;
17'h10e20:	data_out=16'h8956;
17'h10e21:	data_out=16'h6c6;
17'h10e22:	data_out=16'h89a9;
17'h10e23:	data_out=16'h9f7;
17'h10e24:	data_out=16'h9f7;
17'h10e25:	data_out=16'h85ba;
17'h10e26:	data_out=16'h89ce;
17'h10e27:	data_out=16'h9fe;
17'h10e28:	data_out=16'h2b5;
17'h10e29:	data_out=16'h8a00;
17'h10e2a:	data_out=16'h89c0;
17'h10e2b:	data_out=16'h231;
17'h10e2c:	data_out=16'h89f6;
17'h10e2d:	data_out=16'ha00;
17'h10e2e:	data_out=16'h891c;
17'h10e2f:	data_out=16'h89c4;
17'h10e30:	data_out=16'h9d8;
17'h10e31:	data_out=16'ha00;
17'h10e32:	data_out=16'h9e2;
17'h10e33:	data_out=16'h89e4;
17'h10e34:	data_out=16'ha00;
17'h10e35:	data_out=16'h9f7;
17'h10e36:	data_out=16'h89ec;
17'h10e37:	data_out=16'h89fb;
17'h10e38:	data_out=16'h9fa;
17'h10e39:	data_out=16'h89f2;
17'h10e3a:	data_out=16'h89e9;
17'h10e3b:	data_out=16'h9ec;
17'h10e3c:	data_out=16'h87b9;
17'h10e3d:	data_out=16'h88d7;
17'h10e3e:	data_out=16'h298;
17'h10e3f:	data_out=16'h950;
17'h10e40:	data_out=16'h9fb;
17'h10e41:	data_out=16'h8a00;
17'h10e42:	data_out=16'h8273;
17'h10e43:	data_out=16'h89fc;
17'h10e44:	data_out=16'ha00;
17'h10e45:	data_out=16'h89f7;
17'h10e46:	data_out=16'h87f5;
17'h10e47:	data_out=16'h89ff;
17'h10e48:	data_out=16'h880d;
17'h10e49:	data_out=16'h8325;
17'h10e4a:	data_out=16'h89fd;
17'h10e4b:	data_out=16'h89cd;
17'h10e4c:	data_out=16'h8203;
17'h10e4d:	data_out=16'h8968;
17'h10e4e:	data_out=16'h8a00;
17'h10e4f:	data_out=16'h8573;
17'h10e50:	data_out=16'h89d4;
17'h10e51:	data_out=16'h8a00;
17'h10e52:	data_out=16'h9c6;
17'h10e53:	data_out=16'h898d;
17'h10e54:	data_out=16'h899e;
17'h10e55:	data_out=16'h89ff;
17'h10e56:	data_out=16'h88ec;
17'h10e57:	data_out=16'h899e;
17'h10e58:	data_out=16'h8a00;
17'h10e59:	data_out=16'h9f5;
17'h10e5a:	data_out=16'h89ea;
17'h10e5b:	data_out=16'ha00;
17'h10e5c:	data_out=16'h89c6;
17'h10e5d:	data_out=16'h8964;
17'h10e5e:	data_out=16'h8926;
17'h10e5f:	data_out=16'h89eb;
17'h10e60:	data_out=16'h89ee;
17'h10e61:	data_out=16'h9e0;
17'h10e62:	data_out=16'h890f;
17'h10e63:	data_out=16'h89db;
17'h10e64:	data_out=16'ha00;
17'h10e65:	data_out=16'ha00;
17'h10e66:	data_out=16'h8965;
17'h10e67:	data_out=16'h89bb;
17'h10e68:	data_out=16'h513;
17'h10e69:	data_out=16'h8a00;
17'h10e6a:	data_out=16'h9ff;
17'h10e6b:	data_out=16'h81db;
17'h10e6c:	data_out=16'h88b6;
17'h10e6d:	data_out=16'h89dc;
17'h10e6e:	data_out=16'h9ff;
17'h10e6f:	data_out=16'h9ea;
17'h10e70:	data_out=16'h9ff;
17'h10e71:	data_out=16'h8a00;
17'h10e72:	data_out=16'h9f0;
17'h10e73:	data_out=16'ha00;
17'h10e74:	data_out=16'h9c3;
17'h10e75:	data_out=16'h8319;
17'h10e76:	data_out=16'h84f4;
17'h10e77:	data_out=16'h89fd;
17'h10e78:	data_out=16'h89fc;
17'h10e79:	data_out=16'h8a00;
17'h10e7a:	data_out=16'h89dc;
17'h10e7b:	data_out=16'h28c;
17'h10e7c:	data_out=16'h8a00;
17'h10e7d:	data_out=16'h89f1;
17'h10e7e:	data_out=16'h48e;
17'h10e7f:	data_out=16'h89f7;
17'h10e80:	data_out=16'h868c;
17'h10e81:	data_out=16'ha00;
17'h10e82:	data_out=16'h8a00;
17'h10e83:	data_out=16'h89db;
17'h10e84:	data_out=16'h9fe;
17'h10e85:	data_out=16'h9ec;
17'h10e86:	data_out=16'ha00;
17'h10e87:	data_out=16'h8a00;
17'h10e88:	data_out=16'h8a00;
17'h10e89:	data_out=16'h8714;
17'h10e8a:	data_out=16'ha00;
17'h10e8b:	data_out=16'h896e;
17'h10e8c:	data_out=16'h8a00;
17'h10e8d:	data_out=16'h8a00;
17'h10e8e:	data_out=16'h89e8;
17'h10e8f:	data_out=16'h8a00;
17'h10e90:	data_out=16'h8301;
17'h10e91:	data_out=16'ha00;
17'h10e92:	data_out=16'h8a00;
17'h10e93:	data_out=16'h54c;
17'h10e94:	data_out=16'h89ff;
17'h10e95:	data_out=16'h89d6;
17'h10e96:	data_out=16'h8989;
17'h10e97:	data_out=16'h89f8;
17'h10e98:	data_out=16'h8a00;
17'h10e99:	data_out=16'h9ed;
17'h10e9a:	data_out=16'h9f4;
17'h10e9b:	data_out=16'h8a00;
17'h10e9c:	data_out=16'h8a00;
17'h10e9d:	data_out=16'ha00;
17'h10e9e:	data_out=16'h89fd;
17'h10e9f:	data_out=16'h89c6;
17'h10ea0:	data_out=16'h870f;
17'h10ea1:	data_out=16'h89ea;
17'h10ea2:	data_out=16'h9ff;
17'h10ea3:	data_out=16'ha00;
17'h10ea4:	data_out=16'ha00;
17'h10ea5:	data_out=16'h9f9;
17'h10ea6:	data_out=16'h89e4;
17'h10ea7:	data_out=16'h385;
17'h10ea8:	data_out=16'h89ee;
17'h10ea9:	data_out=16'h8a00;
17'h10eaa:	data_out=16'h89ac;
17'h10eab:	data_out=16'h8722;
17'h10eac:	data_out=16'h895b;
17'h10ead:	data_out=16'ha00;
17'h10eae:	data_out=16'h88eb;
17'h10eaf:	data_out=16'h889f;
17'h10eb0:	data_out=16'h9ea;
17'h10eb1:	data_out=16'ha00;
17'h10eb2:	data_out=16'ha00;
17'h10eb3:	data_out=16'h8a00;
17'h10eb4:	data_out=16'ha00;
17'h10eb5:	data_out=16'h8303;
17'h10eb6:	data_out=16'h8a00;
17'h10eb7:	data_out=16'h8a00;
17'h10eb8:	data_out=16'h9fe;
17'h10eb9:	data_out=16'h8a00;
17'h10eba:	data_out=16'h87b5;
17'h10ebb:	data_out=16'h9d0;
17'h10ebc:	data_out=16'h8937;
17'h10ebd:	data_out=16'h84c5;
17'h10ebe:	data_out=16'h89ee;
17'h10ebf:	data_out=16'h9e9;
17'h10ec0:	data_out=16'ha00;
17'h10ec1:	data_out=16'h8a00;
17'h10ec2:	data_out=16'h9be;
17'h10ec3:	data_out=16'h8a00;
17'h10ec4:	data_out=16'h9f7;
17'h10ec5:	data_out=16'h89d3;
17'h10ec6:	data_out=16'h89f2;
17'h10ec7:	data_out=16'h89d9;
17'h10ec8:	data_out=16'h8088;
17'h10ec9:	data_out=16'h9e4;
17'h10eca:	data_out=16'h89ff;
17'h10ecb:	data_out=16'h9f1;
17'h10ecc:	data_out=16'h9ec;
17'h10ecd:	data_out=16'ha00;
17'h10ece:	data_out=16'h8a00;
17'h10ecf:	data_out=16'h9ff;
17'h10ed0:	data_out=16'h85c2;
17'h10ed1:	data_out=16'h8a00;
17'h10ed2:	data_out=16'h9de;
17'h10ed3:	data_out=16'h89ab;
17'h10ed4:	data_out=16'h8887;
17'h10ed5:	data_out=16'h8a00;
17'h10ed6:	data_out=16'h89ff;
17'h10ed7:	data_out=16'h89b7;
17'h10ed8:	data_out=16'h8a00;
17'h10ed9:	data_out=16'ha00;
17'h10eda:	data_out=16'h8a00;
17'h10edb:	data_out=16'ha00;
17'h10edc:	data_out=16'h89e6;
17'h10edd:	data_out=16'h8415;
17'h10ede:	data_out=16'h8611;
17'h10edf:	data_out=16'h89b3;
17'h10ee0:	data_out=16'h89c3;
17'h10ee1:	data_out=16'ha00;
17'h10ee2:	data_out=16'h88ac;
17'h10ee3:	data_out=16'h8a00;
17'h10ee4:	data_out=16'h9ef;
17'h10ee5:	data_out=16'ha00;
17'h10ee6:	data_out=16'h8a00;
17'h10ee7:	data_out=16'h8995;
17'h10ee8:	data_out=16'h89ec;
17'h10ee9:	data_out=16'h8a00;
17'h10eea:	data_out=16'h89e7;
17'h10eeb:	data_out=16'h9ef;
17'h10eec:	data_out=16'h9d2;
17'h10eed:	data_out=16'h8a00;
17'h10eee:	data_out=16'h89e7;
17'h10eef:	data_out=16'h9f9;
17'h10ef0:	data_out=16'h89e8;
17'h10ef1:	data_out=16'h8a00;
17'h10ef2:	data_out=16'ha00;
17'h10ef3:	data_out=16'ha00;
17'h10ef4:	data_out=16'h9b9;
17'h10ef5:	data_out=16'h881e;
17'h10ef6:	data_out=16'h8726;
17'h10ef7:	data_out=16'h8996;
17'h10ef8:	data_out=16'h8463;
17'h10ef9:	data_out=16'h8a00;
17'h10efa:	data_out=16'h8a00;
17'h10efb:	data_out=16'h89ee;
17'h10efc:	data_out=16'h8a00;
17'h10efd:	data_out=16'h89fe;
17'h10efe:	data_out=16'h9ff;
17'h10eff:	data_out=16'h89da;
17'h10f00:	data_out=16'h90f;
17'h10f01:	data_out=16'h9fd;
17'h10f02:	data_out=16'h8a00;
17'h10f03:	data_out=16'h89f0;
17'h10f04:	data_out=16'ha00;
17'h10f05:	data_out=16'h9d9;
17'h10f06:	data_out=16'ha00;
17'h10f07:	data_out=16'h8a00;
17'h10f08:	data_out=16'h8a00;
17'h10f09:	data_out=16'ha00;
17'h10f0a:	data_out=16'ha00;
17'h10f0b:	data_out=16'h8864;
17'h10f0c:	data_out=16'h86d1;
17'h10f0d:	data_out=16'h8a00;
17'h10f0e:	data_out=16'h8a00;
17'h10f0f:	data_out=16'h8a00;
17'h10f10:	data_out=16'ha00;
17'h10f11:	data_out=16'ha00;
17'h10f12:	data_out=16'h8a00;
17'h10f13:	data_out=16'h89f6;
17'h10f14:	data_out=16'h8a00;
17'h10f15:	data_out=16'h89f2;
17'h10f16:	data_out=16'h898b;
17'h10f17:	data_out=16'h8a00;
17'h10f18:	data_out=16'h8a00;
17'h10f19:	data_out=16'h9fb;
17'h10f1a:	data_out=16'h9ff;
17'h10f1b:	data_out=16'h8a00;
17'h10f1c:	data_out=16'h8a00;
17'h10f1d:	data_out=16'ha00;
17'h10f1e:	data_out=16'h8a00;
17'h10f1f:	data_out=16'h8a00;
17'h10f20:	data_out=16'h860c;
17'h10f21:	data_out=16'h8a00;
17'h10f22:	data_out=16'ha00;
17'h10f23:	data_out=16'ha00;
17'h10f24:	data_out=16'ha00;
17'h10f25:	data_out=16'ha00;
17'h10f26:	data_out=16'h89ff;
17'h10f27:	data_out=16'h85f4;
17'h10f28:	data_out=16'h8a00;
17'h10f29:	data_out=16'h8a00;
17'h10f2a:	data_out=16'h89f6;
17'h10f2b:	data_out=16'h895c;
17'h10f2c:	data_out=16'h88dd;
17'h10f2d:	data_out=16'h9fe;
17'h10f2e:	data_out=16'h897c;
17'h10f2f:	data_out=16'h883a;
17'h10f30:	data_out=16'h91c;
17'h10f31:	data_out=16'ha00;
17'h10f32:	data_out=16'ha00;
17'h10f33:	data_out=16'h8a00;
17'h10f34:	data_out=16'ha00;
17'h10f35:	data_out=16'h8612;
17'h10f36:	data_out=16'h8a00;
17'h10f37:	data_out=16'h8a00;
17'h10f38:	data_out=16'h9fd;
17'h10f39:	data_out=16'h8a00;
17'h10f3a:	data_out=16'h9fd;
17'h10f3b:	data_out=16'h9c0;
17'h10f3c:	data_out=16'h89e4;
17'h10f3d:	data_out=16'h9b1;
17'h10f3e:	data_out=16'h8a00;
17'h10f3f:	data_out=16'h9d7;
17'h10f40:	data_out=16'ha00;
17'h10f41:	data_out=16'h8a00;
17'h10f42:	data_out=16'h9ff;
17'h10f43:	data_out=16'h8a00;
17'h10f44:	data_out=16'h2cc;
17'h10f45:	data_out=16'h89ef;
17'h10f46:	data_out=16'h8a00;
17'h10f47:	data_out=16'h89c6;
17'h10f48:	data_out=16'ha00;
17'h10f49:	data_out=16'h9f7;
17'h10f4a:	data_out=16'h8932;
17'h10f4b:	data_out=16'h9ff;
17'h10f4c:	data_out=16'h9fb;
17'h10f4d:	data_out=16'ha00;
17'h10f4e:	data_out=16'h8a00;
17'h10f4f:	data_out=16'ha00;
17'h10f50:	data_out=16'h9fb;
17'h10f51:	data_out=16'h8a00;
17'h10f52:	data_out=16'ha00;
17'h10f53:	data_out=16'h8a00;
17'h10f54:	data_out=16'h88d5;
17'h10f55:	data_out=16'h8a00;
17'h10f56:	data_out=16'h8a00;
17'h10f57:	data_out=16'h89f9;
17'h10f58:	data_out=16'h8a00;
17'h10f59:	data_out=16'ha00;
17'h10f5a:	data_out=16'h8a00;
17'h10f5b:	data_out=16'h884d;
17'h10f5c:	data_out=16'h8a00;
17'h10f5d:	data_out=16'h82f;
17'h10f5e:	data_out=16'h81a4;
17'h10f5f:	data_out=16'h8977;
17'h10f60:	data_out=16'h89cc;
17'h10f61:	data_out=16'h9fa;
17'h10f62:	data_out=16'h898d;
17'h10f63:	data_out=16'h8a00;
17'h10f64:	data_out=16'h9d5;
17'h10f65:	data_out=16'ha00;
17'h10f66:	data_out=16'h8a00;
17'h10f67:	data_out=16'h89d4;
17'h10f68:	data_out=16'h8a00;
17'h10f69:	data_out=16'h8a00;
17'h10f6a:	data_out=16'h8a00;
17'h10f6b:	data_out=16'ha00;
17'h10f6c:	data_out=16'h9c5;
17'h10f6d:	data_out=16'h8a00;
17'h10f6e:	data_out=16'h8a00;
17'h10f6f:	data_out=16'h9ed;
17'h10f70:	data_out=16'h8a00;
17'h10f71:	data_out=16'h8a00;
17'h10f72:	data_out=16'ha00;
17'h10f73:	data_out=16'h9e2;
17'h10f74:	data_out=16'h85d;
17'h10f75:	data_out=16'h89e7;
17'h10f76:	data_out=16'h88e4;
17'h10f77:	data_out=16'h88c6;
17'h10f78:	data_out=16'h75f;
17'h10f79:	data_out=16'h8a00;
17'h10f7a:	data_out=16'h8a00;
17'h10f7b:	data_out=16'h8a00;
17'h10f7c:	data_out=16'h8a00;
17'h10f7d:	data_out=16'h8a00;
17'h10f7e:	data_out=16'ha00;
17'h10f7f:	data_out=16'h820c;
17'h10f80:	data_out=16'h99e;
17'h10f81:	data_out=16'h7b3;
17'h10f82:	data_out=16'h8a00;
17'h10f83:	data_out=16'h89f0;
17'h10f84:	data_out=16'ha00;
17'h10f85:	data_out=16'h61a;
17'h10f86:	data_out=16'ha00;
17'h10f87:	data_out=16'h89f8;
17'h10f88:	data_out=16'h8a00;
17'h10f89:	data_out=16'ha00;
17'h10f8a:	data_out=16'ha00;
17'h10f8b:	data_out=16'h89d1;
17'h10f8c:	data_out=16'h8014;
17'h10f8d:	data_out=16'h8a00;
17'h10f8e:	data_out=16'h8a00;
17'h10f8f:	data_out=16'h8a00;
17'h10f90:	data_out=16'ha00;
17'h10f91:	data_out=16'ha00;
17'h10f92:	data_out=16'h8a00;
17'h10f93:	data_out=16'h8a00;
17'h10f94:	data_out=16'h8a00;
17'h10f95:	data_out=16'h8862;
17'h10f96:	data_out=16'h2e;
17'h10f97:	data_out=16'h8a00;
17'h10f98:	data_out=16'h8a00;
17'h10f99:	data_out=16'h89fb;
17'h10f9a:	data_out=16'h9fa;
17'h10f9b:	data_out=16'h8a00;
17'h10f9c:	data_out=16'h8a00;
17'h10f9d:	data_out=16'h9fe;
17'h10f9e:	data_out=16'h8a00;
17'h10f9f:	data_out=16'h8a00;
17'h10fa0:	data_out=16'h95c;
17'h10fa1:	data_out=16'h8a00;
17'h10fa2:	data_out=16'ha00;
17'h10fa3:	data_out=16'h4a3;
17'h10fa4:	data_out=16'h47f;
17'h10fa5:	data_out=16'h9fc;
17'h10fa6:	data_out=16'h8a00;
17'h10fa7:	data_out=16'h89f9;
17'h10fa8:	data_out=16'h8a00;
17'h10fa9:	data_out=16'h8a00;
17'h10faa:	data_out=16'h8a00;
17'h10fab:	data_out=16'h8a00;
17'h10fac:	data_out=16'h9ea;
17'h10fad:	data_out=16'h9bf;
17'h10fae:	data_out=16'h8a00;
17'h10faf:	data_out=16'h9d8;
17'h10fb0:	data_out=16'h8033;
17'h10fb1:	data_out=16'h9f1;
17'h10fb2:	data_out=16'ha00;
17'h10fb3:	data_out=16'h8a00;
17'h10fb4:	data_out=16'h9cd;
17'h10fb5:	data_out=16'h89df;
17'h10fb6:	data_out=16'h8a00;
17'h10fb7:	data_out=16'h8a00;
17'h10fb8:	data_out=16'h96c;
17'h10fb9:	data_out=16'h8a00;
17'h10fba:	data_out=16'ha00;
17'h10fbb:	data_out=16'had;
17'h10fbc:	data_out=16'h8a00;
17'h10fbd:	data_out=16'h9bd;
17'h10fbe:	data_out=16'h8a00;
17'h10fbf:	data_out=16'h64b;
17'h10fc0:	data_out=16'ha00;
17'h10fc1:	data_out=16'h8a00;
17'h10fc2:	data_out=16'ha00;
17'h10fc3:	data_out=16'h8a00;
17'h10fc4:	data_out=16'h89ff;
17'h10fc5:	data_out=16'h8827;
17'h10fc6:	data_out=16'h8a00;
17'h10fc7:	data_out=16'h86aa;
17'h10fc8:	data_out=16'ha00;
17'h10fc9:	data_out=16'h9ff;
17'h10fca:	data_out=16'h821f;
17'h10fcb:	data_out=16'ha00;
17'h10fcc:	data_out=16'h9fd;
17'h10fcd:	data_out=16'ha00;
17'h10fce:	data_out=16'h8a00;
17'h10fcf:	data_out=16'ha00;
17'h10fd0:	data_out=16'ha00;
17'h10fd1:	data_out=16'h8a00;
17'h10fd2:	data_out=16'h9ff;
17'h10fd3:	data_out=16'h8a00;
17'h10fd4:	data_out=16'h845;
17'h10fd5:	data_out=16'h8a00;
17'h10fd6:	data_out=16'h8a00;
17'h10fd7:	data_out=16'h8a00;
17'h10fd8:	data_out=16'h8a00;
17'h10fd9:	data_out=16'ha00;
17'h10fda:	data_out=16'h8a00;
17'h10fdb:	data_out=16'h8a00;
17'h10fdc:	data_out=16'h8a00;
17'h10fdd:	data_out=16'ha00;
17'h10fde:	data_out=16'ha00;
17'h10fdf:	data_out=16'h8448;
17'h10fe0:	data_out=16'h8a00;
17'h10fe1:	data_out=16'h86ff;
17'h10fe2:	data_out=16'h89fc;
17'h10fe3:	data_out=16'h8a00;
17'h10fe4:	data_out=16'h9c6;
17'h10fe5:	data_out=16'ha00;
17'h10fe6:	data_out=16'h8a00;
17'h10fe7:	data_out=16'h8a00;
17'h10fe8:	data_out=16'h8a00;
17'h10fe9:	data_out=16'h8a00;
17'h10fea:	data_out=16'h8a00;
17'h10feb:	data_out=16'ha00;
17'h10fec:	data_out=16'h9d4;
17'h10fed:	data_out=16'h8a00;
17'h10fee:	data_out=16'h8a00;
17'h10fef:	data_out=16'h9d7;
17'h10ff0:	data_out=16'h8a00;
17'h10ff1:	data_out=16'h8a00;
17'h10ff2:	data_out=16'ha00;
17'h10ff3:	data_out=16'h9dc;
17'h10ff4:	data_out=16'h8142;
17'h10ff5:	data_out=16'h8a00;
17'h10ff6:	data_out=16'h8a00;
17'h10ff7:	data_out=16'h8287;
17'h10ff8:	data_out=16'h894f;
17'h10ff9:	data_out=16'h8a00;
17'h10ffa:	data_out=16'h8a00;
17'h10ffb:	data_out=16'h8a00;
17'h10ffc:	data_out=16'h8a00;
17'h10ffd:	data_out=16'h8a00;
17'h10ffe:	data_out=16'h9fe;
17'h10fff:	data_out=16'ha00;
17'h11000:	data_out=16'h977;
17'h11001:	data_out=16'h47f;
17'h11002:	data_out=16'h8a00;
17'h11003:	data_out=16'h89f4;
17'h11004:	data_out=16'h9fc;
17'h11005:	data_out=16'h89d0;
17'h11006:	data_out=16'h9fc;
17'h11007:	data_out=16'h8a00;
17'h11008:	data_out=16'h8a00;
17'h11009:	data_out=16'h9da;
17'h1100a:	data_out=16'ha00;
17'h1100b:	data_out=16'h8a00;
17'h1100c:	data_out=16'h88c9;
17'h1100d:	data_out=16'h8a00;
17'h1100e:	data_out=16'h8a00;
17'h1100f:	data_out=16'h8a00;
17'h11010:	data_out=16'ha00;
17'h11011:	data_out=16'ha00;
17'h11012:	data_out=16'h8a00;
17'h11013:	data_out=16'h881e;
17'h11014:	data_out=16'h8a00;
17'h11015:	data_out=16'h1fe;
17'h11016:	data_out=16'h989;
17'h11017:	data_out=16'h8a00;
17'h11018:	data_out=16'h8a00;
17'h11019:	data_out=16'h8a00;
17'h1101a:	data_out=16'h994;
17'h1101b:	data_out=16'h8a00;
17'h1101c:	data_out=16'h8a00;
17'h1101d:	data_out=16'h9fc;
17'h1101e:	data_out=16'h8a00;
17'h1101f:	data_out=16'h8a00;
17'h11020:	data_out=16'h57a;
17'h11021:	data_out=16'h8a00;
17'h11022:	data_out=16'h9fe;
17'h11023:	data_out=16'h89fd;
17'h11024:	data_out=16'h89fd;
17'h11025:	data_out=16'h805d;
17'h11026:	data_out=16'h8a00;
17'h11027:	data_out=16'h8a00;
17'h11028:	data_out=16'h8a00;
17'h11029:	data_out=16'h8a00;
17'h1102a:	data_out=16'h8a00;
17'h1102b:	data_out=16'h8a00;
17'h1102c:	data_out=16'h9ab;
17'h1102d:	data_out=16'h9b4;
17'h1102e:	data_out=16'h8a00;
17'h1102f:	data_out=16'h7d7;
17'h11030:	data_out=16'h8708;
17'h11031:	data_out=16'h0;
17'h11032:	data_out=16'h9ff;
17'h11033:	data_out=16'h8a00;
17'h11034:	data_out=16'h9dd;
17'h11035:	data_out=16'h8a00;
17'h11036:	data_out=16'h8a00;
17'h11037:	data_out=16'h8a00;
17'h11038:	data_out=16'h9e9;
17'h11039:	data_out=16'h8a00;
17'h1103a:	data_out=16'h9f0;
17'h1103b:	data_out=16'h8a00;
17'h1103c:	data_out=16'h8a00;
17'h1103d:	data_out=16'h854;
17'h1103e:	data_out=16'h8a00;
17'h1103f:	data_out=16'h89ca;
17'h11040:	data_out=16'h9ff;
17'h11041:	data_out=16'h8a00;
17'h11042:	data_out=16'ha00;
17'h11043:	data_out=16'h8a00;
17'h11044:	data_out=16'h8a00;
17'h11045:	data_out=16'h13b;
17'h11046:	data_out=16'h8a00;
17'h11047:	data_out=16'h89fd;
17'h11048:	data_out=16'ha00;
17'h11049:	data_out=16'h184;
17'h1104a:	data_out=16'h80b5;
17'h1104b:	data_out=16'h9ff;
17'h1104c:	data_out=16'h9f9;
17'h1104d:	data_out=16'ha00;
17'h1104e:	data_out=16'h8a00;
17'h1104f:	data_out=16'ha00;
17'h11050:	data_out=16'h9ff;
17'h11051:	data_out=16'h8a00;
17'h11052:	data_out=16'h899b;
17'h11053:	data_out=16'h8a00;
17'h11054:	data_out=16'h4d9;
17'h11055:	data_out=16'h8a00;
17'h11056:	data_out=16'h8a00;
17'h11057:	data_out=16'h8a00;
17'h11058:	data_out=16'h8a00;
17'h11059:	data_out=16'ha00;
17'h1105a:	data_out=16'h8a00;
17'h1105b:	data_out=16'h8a00;
17'h1105c:	data_out=16'h8a00;
17'h1105d:	data_out=16'h9ff;
17'h1105e:	data_out=16'ha00;
17'h1105f:	data_out=16'h9e4;
17'h11060:	data_out=16'h8a00;
17'h11061:	data_out=16'h899a;
17'h11062:	data_out=16'h8a00;
17'h11063:	data_out=16'h8a00;
17'h11064:	data_out=16'h993;
17'h11065:	data_out=16'ha00;
17'h11066:	data_out=16'h8a00;
17'h11067:	data_out=16'h8a00;
17'h11068:	data_out=16'h8a00;
17'h11069:	data_out=16'h8a00;
17'h1106a:	data_out=16'h8a00;
17'h1106b:	data_out=16'h942;
17'h1106c:	data_out=16'h9ce;
17'h1106d:	data_out=16'h8a00;
17'h1106e:	data_out=16'h8a00;
17'h1106f:	data_out=16'h642;
17'h11070:	data_out=16'h8a00;
17'h11071:	data_out=16'h8a00;
17'h11072:	data_out=16'h9fe;
17'h11073:	data_out=16'h9d8;
17'h11074:	data_out=16'h88ff;
17'h11075:	data_out=16'h8a00;
17'h11076:	data_out=16'h8a00;
17'h11077:	data_out=16'h84e3;
17'h11078:	data_out=16'h8935;
17'h11079:	data_out=16'h8529;
17'h1107a:	data_out=16'h8a00;
17'h1107b:	data_out=16'h8a00;
17'h1107c:	data_out=16'h8a00;
17'h1107d:	data_out=16'h8a00;
17'h1107e:	data_out=16'h4c5;
17'h1107f:	data_out=16'ha00;
17'h11080:	data_out=16'h8b3;
17'h11081:	data_out=16'h89ff;
17'h11082:	data_out=16'h8a00;
17'h11083:	data_out=16'h945;
17'h11084:	data_out=16'h872;
17'h11085:	data_out=16'h379;
17'h11086:	data_out=16'h9f5;
17'h11087:	data_out=16'h89f5;
17'h11088:	data_out=16'h8a00;
17'h11089:	data_out=16'h9f9;
17'h1108a:	data_out=16'ha00;
17'h1108b:	data_out=16'h8a00;
17'h1108c:	data_out=16'h8915;
17'h1108d:	data_out=16'h8176;
17'h1108e:	data_out=16'h89ff;
17'h1108f:	data_out=16'h8a00;
17'h11090:	data_out=16'ha00;
17'h11091:	data_out=16'h9ff;
17'h11092:	data_out=16'h8a00;
17'h11093:	data_out=16'h967;
17'h11094:	data_out=16'h8a00;
17'h11095:	data_out=16'h99d;
17'h11096:	data_out=16'h9c2;
17'h11097:	data_out=16'h89fe;
17'h11098:	data_out=16'h8a00;
17'h11099:	data_out=16'h8a00;
17'h1109a:	data_out=16'h8e6;
17'h1109b:	data_out=16'h8a00;
17'h1109c:	data_out=16'h8a00;
17'h1109d:	data_out=16'h107;
17'h1109e:	data_out=16'h31f;
17'h1109f:	data_out=16'h8a00;
17'h110a0:	data_out=16'h7a2;
17'h110a1:	data_out=16'h89ff;
17'h110a2:	data_out=16'h9f9;
17'h110a3:	data_out=16'h8a00;
17'h110a4:	data_out=16'h8a00;
17'h110a5:	data_out=16'h8221;
17'h110a6:	data_out=16'h8a00;
17'h110a7:	data_out=16'h8a00;
17'h110a8:	data_out=16'h89ff;
17'h110a9:	data_out=16'h8a00;
17'h110aa:	data_out=16'h89f9;
17'h110ab:	data_out=16'h8a00;
17'h110ac:	data_out=16'h9d8;
17'h110ad:	data_out=16'h89fc;
17'h110ae:	data_out=16'h8a00;
17'h110af:	data_out=16'h945;
17'h110b0:	data_out=16'h83d9;
17'h110b1:	data_out=16'h89ff;
17'h110b2:	data_out=16'h84d;
17'h110b3:	data_out=16'h8a00;
17'h110b4:	data_out=16'h8d3;
17'h110b5:	data_out=16'h89fd;
17'h110b6:	data_out=16'h8a00;
17'h110b7:	data_out=16'h8a00;
17'h110b8:	data_out=16'ha00;
17'h110b9:	data_out=16'h8a00;
17'h110ba:	data_out=16'h9fb;
17'h110bb:	data_out=16'h8a00;
17'h110bc:	data_out=16'h8a00;
17'h110bd:	data_out=16'h8da;
17'h110be:	data_out=16'h89ff;
17'h110bf:	data_out=16'h3d6;
17'h110c0:	data_out=16'h9ef;
17'h110c1:	data_out=16'h89e3;
17'h110c2:	data_out=16'h9f1;
17'h110c3:	data_out=16'h8a00;
17'h110c4:	data_out=16'h8a00;
17'h110c5:	data_out=16'h9ac;
17'h110c6:	data_out=16'h8a00;
17'h110c7:	data_out=16'h911;
17'h110c8:	data_out=16'h9ff;
17'h110c9:	data_out=16'h84a8;
17'h110ca:	data_out=16'h92a;
17'h110cb:	data_out=16'h9f7;
17'h110cc:	data_out=16'h5db;
17'h110cd:	data_out=16'ha00;
17'h110ce:	data_out=16'h96f;
17'h110cf:	data_out=16'h4e4;
17'h110d0:	data_out=16'ha00;
17'h110d1:	data_out=16'h8a00;
17'h110d2:	data_out=16'h89fb;
17'h110d3:	data_out=16'h8a00;
17'h110d4:	data_out=16'h836;
17'h110d5:	data_out=16'h8a00;
17'h110d6:	data_out=16'h8a00;
17'h110d7:	data_out=16'h8a00;
17'h110d8:	data_out=16'h8a00;
17'h110d9:	data_out=16'ha00;
17'h110da:	data_out=16'h8a00;
17'h110db:	data_out=16'h8a00;
17'h110dc:	data_out=16'h8a00;
17'h110dd:	data_out=16'h9fa;
17'h110de:	data_out=16'ha00;
17'h110df:	data_out=16'h9e6;
17'h110e0:	data_out=16'h8a00;
17'h110e1:	data_out=16'h89d1;
17'h110e2:	data_out=16'h8a00;
17'h110e3:	data_out=16'h8a00;
17'h110e4:	data_out=16'h8bf;
17'h110e5:	data_out=16'h9f6;
17'h110e6:	data_out=16'h89f9;
17'h110e7:	data_out=16'h8a00;
17'h110e8:	data_out=16'h89ff;
17'h110e9:	data_out=16'h8a00;
17'h110ea:	data_out=16'h89ff;
17'h110eb:	data_out=16'h9ac;
17'h110ec:	data_out=16'h93b;
17'h110ed:	data_out=16'h8a00;
17'h110ee:	data_out=16'h89ff;
17'h110ef:	data_out=16'h9cb;
17'h110f0:	data_out=16'h89ff;
17'h110f1:	data_out=16'h8a00;
17'h110f2:	data_out=16'h9fe;
17'h110f3:	data_out=16'h82cf;
17'h110f4:	data_out=16'h863c;
17'h110f5:	data_out=16'h8a00;
17'h110f6:	data_out=16'h8a00;
17'h110f7:	data_out=16'h9ea;
17'h110f8:	data_out=16'h8979;
17'h110f9:	data_out=16'h9fc;
17'h110fa:	data_out=16'h8a00;
17'h110fb:	data_out=16'h89ff;
17'h110fc:	data_out=16'h8a00;
17'h110fd:	data_out=16'h89fd;
17'h110fe:	data_out=16'h7b7;
17'h110ff:	data_out=16'ha00;
17'h11100:	data_out=16'he3;
17'h11101:	data_out=16'h8a00;
17'h11102:	data_out=16'h8a00;
17'h11103:	data_out=16'h5bc;
17'h11104:	data_out=16'h8a00;
17'h11105:	data_out=16'h8540;
17'h11106:	data_out=16'h9df;
17'h11107:	data_out=16'h81d;
17'h11108:	data_out=16'h8a00;
17'h11109:	data_out=16'h9fa;
17'h1110a:	data_out=16'h89f9;
17'h1110b:	data_out=16'h89ff;
17'h1110c:	data_out=16'h9c0;
17'h1110d:	data_out=16'h97c;
17'h1110e:	data_out=16'h8a00;
17'h1110f:	data_out=16'h89f5;
17'h11110:	data_out=16'h9d1;
17'h11111:	data_out=16'h8a00;
17'h11112:	data_out=16'h812c;
17'h11113:	data_out=16'ha00;
17'h11114:	data_out=16'h218;
17'h11115:	data_out=16'h86d;
17'h11116:	data_out=16'h945;
17'h11117:	data_out=16'h62b;
17'h11118:	data_out=16'h8a00;
17'h11119:	data_out=16'h8a00;
17'h1111a:	data_out=16'h311;
17'h1111b:	data_out=16'h8a00;
17'h1111c:	data_out=16'h89fe;
17'h1111d:	data_out=16'h8a00;
17'h1111e:	data_out=16'h91c;
17'h1111f:	data_out=16'h872a;
17'h11120:	data_out=16'h586;
17'h11121:	data_out=16'h8a00;
17'h11122:	data_out=16'h922;
17'h11123:	data_out=16'h8a00;
17'h11124:	data_out=16'h8a00;
17'h11125:	data_out=16'h8238;
17'h11126:	data_out=16'h8a00;
17'h11127:	data_out=16'h8a00;
17'h11128:	data_out=16'h89ff;
17'h11129:	data_out=16'h8a00;
17'h1112a:	data_out=16'h347;
17'h1112b:	data_out=16'h8a00;
17'h1112c:	data_out=16'h96b;
17'h1112d:	data_out=16'h89fe;
17'h1112e:	data_out=16'h89fc;
17'h1112f:	data_out=16'h964;
17'h11130:	data_out=16'h9ff;
17'h11131:	data_out=16'h8a00;
17'h11132:	data_out=16'h160;
17'h11133:	data_out=16'h9a7;
17'h11134:	data_out=16'h89fc;
17'h11135:	data_out=16'h8a00;
17'h11136:	data_out=16'h89ff;
17'h11137:	data_out=16'h8a00;
17'h11138:	data_out=16'ha00;
17'h11139:	data_out=16'h99b;
17'h1113a:	data_out=16'h9fc;
17'h1113b:	data_out=16'h8a00;
17'h1113c:	data_out=16'h8a00;
17'h1113d:	data_out=16'h562;
17'h1113e:	data_out=16'h89ff;
17'h1113f:	data_out=16'h857a;
17'h11140:	data_out=16'h6aa;
17'h11141:	data_out=16'h81f6;
17'h11142:	data_out=16'h7d2;
17'h11143:	data_out=16'h89f2;
17'h11144:	data_out=16'h8a00;
17'h11145:	data_out=16'h885;
17'h11146:	data_out=16'h8a00;
17'h11147:	data_out=16'h9f3;
17'h11148:	data_out=16'ha00;
17'h11149:	data_out=16'h85dc;
17'h1114a:	data_out=16'h9d0;
17'h1114b:	data_out=16'h9b5;
17'h1114c:	data_out=16'h80bc;
17'h1114d:	data_out=16'h9b4;
17'h1114e:	data_out=16'h91e;
17'h1114f:	data_out=16'h71;
17'h11150:	data_out=16'h9dc;
17'h11151:	data_out=16'h89fd;
17'h11152:	data_out=16'h8a00;
17'h11153:	data_out=16'h8a00;
17'h11154:	data_out=16'h6ba;
17'h11155:	data_out=16'h89fc;
17'h11156:	data_out=16'h8a00;
17'h11157:	data_out=16'h8a00;
17'h11158:	data_out=16'h8a00;
17'h11159:	data_out=16'h8569;
17'h1115a:	data_out=16'h89fe;
17'h1115b:	data_out=16'h8a00;
17'h1115c:	data_out=16'h8a00;
17'h1115d:	data_out=16'h9a1;
17'h1115e:	data_out=16'ha00;
17'h1115f:	data_out=16'h9ed;
17'h11160:	data_out=16'h8a00;
17'h11161:	data_out=16'h8a00;
17'h11162:	data_out=16'h89c6;
17'h11163:	data_out=16'h973;
17'h11164:	data_out=16'h76d;
17'h11165:	data_out=16'h883;
17'h11166:	data_out=16'h9d2;
17'h11167:	data_out=16'h8a00;
17'h11168:	data_out=16'h89ff;
17'h11169:	data_out=16'h8a00;
17'h1116a:	data_out=16'h8a00;
17'h1116b:	data_out=16'h80f;
17'h1116c:	data_out=16'hc6;
17'h1116d:	data_out=16'h979;
17'h1116e:	data_out=16'h8a00;
17'h1116f:	data_out=16'h834;
17'h11170:	data_out=16'h8a00;
17'h11171:	data_out=16'h1f5;
17'h11172:	data_out=16'h54e;
17'h11173:	data_out=16'h89fd;
17'h11174:	data_out=16'h9fe;
17'h11175:	data_out=16'h8a00;
17'h11176:	data_out=16'h8a00;
17'h11177:	data_out=16'h9df;
17'h11178:	data_out=16'h89e5;
17'h11179:	data_out=16'h9ff;
17'h1117a:	data_out=16'h6cb;
17'h1117b:	data_out=16'h89ff;
17'h1117c:	data_out=16'h89fd;
17'h1117d:	data_out=16'h9c0;
17'h1117e:	data_out=16'h9c8;
17'h1117f:	data_out=16'h9d0;
17'h11180:	data_out=16'h89fc;
17'h11181:	data_out=16'h8a00;
17'h11182:	data_out=16'h8a00;
17'h11183:	data_out=16'h8816;
17'h11184:	data_out=16'h688;
17'h11185:	data_out=16'h2ae;
17'h11186:	data_out=16'h9b0;
17'h11187:	data_out=16'h9f6;
17'h11188:	data_out=16'h89a5;
17'h11189:	data_out=16'h9d0;
17'h1118a:	data_out=16'h8a00;
17'h1118b:	data_out=16'h89f2;
17'h1118c:	data_out=16'h98d;
17'h1118d:	data_out=16'h223;
17'h1118e:	data_out=16'h5ac;
17'h1118f:	data_out=16'h88c4;
17'h11190:	data_out=16'h847;
17'h11191:	data_out=16'h8a00;
17'h11192:	data_out=16'h89c8;
17'h11193:	data_out=16'h9f5;
17'h11194:	data_out=16'h8462;
17'h11195:	data_out=16'h761;
17'h11196:	data_out=16'h86d;
17'h11197:	data_out=16'h83dc;
17'h11198:	data_out=16'h89f1;
17'h11199:	data_out=16'h97a;
17'h1119a:	data_out=16'h425;
17'h1119b:	data_out=16'h8a00;
17'h1119c:	data_out=16'h88a1;
17'h1119d:	data_out=16'h89ff;
17'h1119e:	data_out=16'h312;
17'h1119f:	data_out=16'h814d;
17'h111a0:	data_out=16'h5f6;
17'h111a1:	data_out=16'h7b7;
17'h111a2:	data_out=16'h8a00;
17'h111a3:	data_out=16'h8a00;
17'h111a4:	data_out=16'h8a00;
17'h111a5:	data_out=16'h82d6;
17'h111a6:	data_out=16'h8a00;
17'h111a7:	data_out=16'h8a00;
17'h111a8:	data_out=16'h950;
17'h111a9:	data_out=16'h8a00;
17'h111aa:	data_out=16'h89ff;
17'h111ab:	data_out=16'h89f8;
17'h111ac:	data_out=16'h94b;
17'h111ad:	data_out=16'h89fc;
17'h111ae:	data_out=16'h89ff;
17'h111af:	data_out=16'h92d;
17'h111b0:	data_out=16'ha00;
17'h111b1:	data_out=16'h8a00;
17'h111b2:	data_out=16'he8;
17'h111b3:	data_out=16'h4b3;
17'h111b4:	data_out=16'h89fd;
17'h111b5:	data_out=16'h803b;
17'h111b6:	data_out=16'h89c6;
17'h111b7:	data_out=16'h8a00;
17'h111b8:	data_out=16'h9ed;
17'h111b9:	data_out=16'h33d;
17'h111ba:	data_out=16'h9ec;
17'h111bb:	data_out=16'h869e;
17'h111bc:	data_out=16'h8a00;
17'h111bd:	data_out=16'h427;
17'h111be:	data_out=16'h952;
17'h111bf:	data_out=16'h28e;
17'h111c0:	data_out=16'h713;
17'h111c1:	data_out=16'h80ca;
17'h111c2:	data_out=16'h89fe;
17'h111c3:	data_out=16'h89c7;
17'h111c4:	data_out=16'h83af;
17'h111c5:	data_out=16'h8d9;
17'h111c6:	data_out=16'h8a00;
17'h111c7:	data_out=16'h8b8;
17'h111c8:	data_out=16'h9dc;
17'h111c9:	data_out=16'h81e0;
17'h111ca:	data_out=16'h9ed;
17'h111cb:	data_out=16'h36b;
17'h111cc:	data_out=16'h878e;
17'h111cd:	data_out=16'h8a00;
17'h111ce:	data_out=16'h4db;
17'h111cf:	data_out=16'h805a;
17'h111d0:	data_out=16'h9d0;
17'h111d1:	data_out=16'h89fa;
17'h111d2:	data_out=16'h8a00;
17'h111d3:	data_out=16'h83d7;
17'h111d4:	data_out=16'h2f3;
17'h111d5:	data_out=16'h89ec;
17'h111d6:	data_out=16'h8a00;
17'h111d7:	data_out=16'h8a00;
17'h111d8:	data_out=16'h89ff;
17'h111d9:	data_out=16'h37b;
17'h111da:	data_out=16'h89cb;
17'h111db:	data_out=16'h8a00;
17'h111dc:	data_out=16'h8a00;
17'h111dd:	data_out=16'h89d;
17'h111de:	data_out=16'ha00;
17'h111df:	data_out=16'h827a;
17'h111e0:	data_out=16'h8a00;
17'h111e1:	data_out=16'h8a00;
17'h111e2:	data_out=16'h89fd;
17'h111e3:	data_out=16'h3ce;
17'h111e4:	data_out=16'h655;
17'h111e5:	data_out=16'h4c9;
17'h111e6:	data_out=16'h9ff;
17'h111e7:	data_out=16'h8a00;
17'h111e8:	data_out=16'h8e1;
17'h111e9:	data_out=16'h89f4;
17'h111ea:	data_out=16'h438;
17'h111eb:	data_out=16'h9c6;
17'h111ec:	data_out=16'h89ff;
17'h111ed:	data_out=16'h405;
17'h111ee:	data_out=16'h440;
17'h111ef:	data_out=16'h988;
17'h111f0:	data_out=16'h50e;
17'h111f1:	data_out=16'h8389;
17'h111f2:	data_out=16'h8c2;
17'h111f3:	data_out=16'h835b;
17'h111f4:	data_out=16'ha00;
17'h111f5:	data_out=16'h8a00;
17'h111f6:	data_out=16'h8a00;
17'h111f7:	data_out=16'h4d7;
17'h111f8:	data_out=16'h89f9;
17'h111f9:	data_out=16'h835f;
17'h111fa:	data_out=16'hcd;
17'h111fb:	data_out=16'h954;
17'h111fc:	data_out=16'h89ec;
17'h111fd:	data_out=16'h9f0;
17'h111fe:	data_out=16'h9b3;
17'h111ff:	data_out=16'h7ed;
17'h11200:	data_out=16'h89b5;
17'h11201:	data_out=16'h89fc;
17'h11202:	data_out=16'h8a00;
17'h11203:	data_out=16'h578;
17'h11204:	data_out=16'h993;
17'h11205:	data_out=16'h71d;
17'h11206:	data_out=16'h722;
17'h11207:	data_out=16'h9fa;
17'h11208:	data_out=16'h89c9;
17'h11209:	data_out=16'h6b1;
17'h1120a:	data_out=16'h89fc;
17'h1120b:	data_out=16'h89bf;
17'h1120c:	data_out=16'h8e6;
17'h1120d:	data_out=16'h1b3;
17'h1120e:	data_out=16'h849;
17'h1120f:	data_out=16'h89ee;
17'h11210:	data_out=16'h612;
17'h11211:	data_out=16'h8a00;
17'h11212:	data_out=16'h89fb;
17'h11213:	data_out=16'h9d9;
17'h11214:	data_out=16'h31c;
17'h11215:	data_out=16'h250;
17'h11216:	data_out=16'h9e3;
17'h11217:	data_out=16'h80d;
17'h11218:	data_out=16'h89fa;
17'h11219:	data_out=16'ha00;
17'h1121a:	data_out=16'h7f4;
17'h1121b:	data_out=16'ha6;
17'h1121c:	data_out=16'h8a00;
17'h1121d:	data_out=16'h8580;
17'h1121e:	data_out=16'h4bf;
17'h1121f:	data_out=16'h41f;
17'h11220:	data_out=16'h6d8;
17'h11221:	data_out=16'h8c5;
17'h11222:	data_out=16'h8a00;
17'h11223:	data_out=16'h89e5;
17'h11224:	data_out=16'h89e5;
17'h11225:	data_out=16'h807e;
17'h11226:	data_out=16'h8a00;
17'h11227:	data_out=16'h5ab;
17'h11228:	data_out=16'h92a;
17'h11229:	data_out=16'h8a00;
17'h1122a:	data_out=16'h89bf;
17'h1122b:	data_out=16'h8808;
17'h1122c:	data_out=16'h9e8;
17'h1122d:	data_out=16'h89fd;
17'h1122e:	data_out=16'h8a00;
17'h1122f:	data_out=16'h9d6;
17'h11230:	data_out=16'ha00;
17'h11231:	data_out=16'h9ba;
17'h11232:	data_out=16'h44e;
17'h11233:	data_out=16'h69;
17'h11234:	data_out=16'h89af;
17'h11235:	data_out=16'h465;
17'h11236:	data_out=16'h89a7;
17'h11237:	data_out=16'h8a00;
17'h11238:	data_out=16'h89cb;
17'h11239:	data_out=16'h88d4;
17'h1123a:	data_out=16'h973;
17'h1123b:	data_out=16'h9fa;
17'h1123c:	data_out=16'h8a00;
17'h1123d:	data_out=16'h825d;
17'h1123e:	data_out=16'h92c;
17'h1123f:	data_out=16'h6f7;
17'h11240:	data_out=16'h824;
17'h11241:	data_out=16'h363;
17'h11242:	data_out=16'h89fa;
17'h11243:	data_out=16'h9f1;
17'h11244:	data_out=16'h9af;
17'h11245:	data_out=16'h4e3;
17'h11246:	data_out=16'h8a00;
17'h11247:	data_out=16'h89af;
17'h11248:	data_out=16'h5c0;
17'h11249:	data_out=16'h44a;
17'h1124a:	data_out=16'h9ff;
17'h1124b:	data_out=16'h89d4;
17'h1124c:	data_out=16'h8a00;
17'h1124d:	data_out=16'h8a00;
17'h1124e:	data_out=16'h552;
17'h1124f:	data_out=16'h87a7;
17'h11250:	data_out=16'h9ed;
17'h11251:	data_out=16'h84e7;
17'h11252:	data_out=16'h89f2;
17'h11253:	data_out=16'h280;
17'h11254:	data_out=16'h802e;
17'h11255:	data_out=16'h850b;
17'h11256:	data_out=16'h8a00;
17'h11257:	data_out=16'h8a00;
17'h11258:	data_out=16'h8156;
17'h11259:	data_out=16'h17e;
17'h1125a:	data_out=16'h8362;
17'h1125b:	data_out=16'h152;
17'h1125c:	data_out=16'h8a00;
17'h1125d:	data_out=16'h9e0;
17'h1125e:	data_out=16'ha00;
17'h1125f:	data_out=16'h89e9;
17'h11260:	data_out=16'h8a00;
17'h11261:	data_out=16'h82e8;
17'h11262:	data_out=16'h85f9;
17'h11263:	data_out=16'h62c;
17'h11264:	data_out=16'h19;
17'h11265:	data_out=16'h6df;
17'h11266:	data_out=16'ha00;
17'h11267:	data_out=16'h8a00;
17'h11268:	data_out=16'h907;
17'h11269:	data_out=16'h8a00;
17'h1126a:	data_out=16'h7de;
17'h1126b:	data_out=16'h9d6;
17'h1126c:	data_out=16'h89e9;
17'h1126d:	data_out=16'h4a7;
17'h1126e:	data_out=16'h7e1;
17'h1126f:	data_out=16'h9ee;
17'h11270:	data_out=16'h825;
17'h11271:	data_out=16'h89d4;
17'h11272:	data_out=16'h77c;
17'h11273:	data_out=16'h160;
17'h11274:	data_out=16'ha00;
17'h11275:	data_out=16'h8a00;
17'h11276:	data_out=16'h8a00;
17'h11277:	data_out=16'h347;
17'h11278:	data_out=16'h85b9;
17'h11279:	data_out=16'h8049;
17'h1127a:	data_out=16'h777;
17'h1127b:	data_out=16'h92c;
17'h1127c:	data_out=16'h89f3;
17'h1127d:	data_out=16'h9ea;
17'h1127e:	data_out=16'h967;
17'h1127f:	data_out=16'h81eb;
17'h11280:	data_out=16'h89a9;
17'h11281:	data_out=16'h88fa;
17'h11282:	data_out=16'h82c7;
17'h11283:	data_out=16'h38;
17'h11284:	data_out=16'h9f8;
17'h11285:	data_out=16'h9e1;
17'h11286:	data_out=16'h89ff;
17'h11287:	data_out=16'ha00;
17'h11288:	data_out=16'h89aa;
17'h11289:	data_out=16'h80c8;
17'h1128a:	data_out=16'h88cb;
17'h1128b:	data_out=16'h67a;
17'h1128c:	data_out=16'h83e;
17'h1128d:	data_out=16'h8a00;
17'h1128e:	data_out=16'h965;
17'h1128f:	data_out=16'h8131;
17'h11290:	data_out=16'h929;
17'h11291:	data_out=16'h89ee;
17'h11292:	data_out=16'h8a00;
17'h11293:	data_out=16'h9da;
17'h11294:	data_out=16'h167;
17'h11295:	data_out=16'h9f0;
17'h11296:	data_out=16'h9ec;
17'h11297:	data_out=16'h6f6;
17'h11298:	data_out=16'h8a00;
17'h11299:	data_out=16'ha00;
17'h1129a:	data_out=16'h9ef;
17'h1129b:	data_out=16'h9ae;
17'h1129c:	data_out=16'h8a00;
17'h1129d:	data_out=16'h445;
17'h1129e:	data_out=16'h8147;
17'h1129f:	data_out=16'h965;
17'h112a0:	data_out=16'h845;
17'h112a1:	data_out=16'h980;
17'h112a2:	data_out=16'h89fc;
17'h112a3:	data_out=16'h702;
17'h112a4:	data_out=16'h74f;
17'h112a5:	data_out=16'h841c;
17'h112a6:	data_out=16'h89ff;
17'h112a7:	data_out=16'h9e3;
17'h112a8:	data_out=16'h9c6;
17'h112a9:	data_out=16'h8941;
17'h112aa:	data_out=16'h8885;
17'h112ab:	data_out=16'h9d1;
17'h112ac:	data_out=16'h9ec;
17'h112ad:	data_out=16'h89f4;
17'h112ae:	data_out=16'h89cb;
17'h112af:	data_out=16'h9f5;
17'h112b0:	data_out=16'ha00;
17'h112b1:	data_out=16'h9e1;
17'h112b2:	data_out=16'ha00;
17'h112b3:	data_out=16'h8692;
17'h112b4:	data_out=16'h8835;
17'h112b5:	data_out=16'h9d2;
17'h112b6:	data_out=16'h8228;
17'h112b7:	data_out=16'hbb;
17'h112b8:	data_out=16'h89ee;
17'h112b9:	data_out=16'h89f5;
17'h112ba:	data_out=16'h734;
17'h112bb:	data_out=16'ha00;
17'h112bc:	data_out=16'h2d3;
17'h112bd:	data_out=16'h8172;
17'h112be:	data_out=16'h9c8;
17'h112bf:	data_out=16'h9e0;
17'h112c0:	data_out=16'h9fb;
17'h112c1:	data_out=16'h48c;
17'h112c2:	data_out=16'h89ea;
17'h112c3:	data_out=16'h9f1;
17'h112c4:	data_out=16'h9c5;
17'h112c5:	data_out=16'h9f0;
17'h112c6:	data_out=16'h89f8;
17'h112c7:	data_out=16'h89c9;
17'h112c8:	data_out=16'h4ba;
17'h112c9:	data_out=16'h929;
17'h112ca:	data_out=16'ha00;
17'h112cb:	data_out=16'h89d8;
17'h112cc:	data_out=16'h8a00;
17'h112cd:	data_out=16'h89c5;
17'h112ce:	data_out=16'h959;
17'h112cf:	data_out=16'h8925;
17'h112d0:	data_out=16'h9f2;
17'h112d1:	data_out=16'h15d;
17'h112d2:	data_out=16'h263;
17'h112d3:	data_out=16'h9f0;
17'h112d4:	data_out=16'h800f;
17'h112d5:	data_out=16'h977;
17'h112d6:	data_out=16'h8937;
17'h112d7:	data_out=16'h8a00;
17'h112d8:	data_out=16'h106;
17'h112d9:	data_out=16'h9e3;
17'h112da:	data_out=16'h810d;
17'h112db:	data_out=16'h9b0;
17'h112dc:	data_out=16'h8214;
17'h112dd:	data_out=16'h9fd;
17'h112de:	data_out=16'ha00;
17'h112df:	data_out=16'h89b5;
17'h112e0:	data_out=16'h89fa;
17'h112e1:	data_out=16'h968;
17'h112e2:	data_out=16'h490;
17'h112e3:	data_out=16'h828d;
17'h112e4:	data_out=16'h8990;
17'h112e5:	data_out=16'ha00;
17'h112e6:	data_out=16'ha00;
17'h112e7:	data_out=16'h9d9;
17'h112e8:	data_out=16'h9a1;
17'h112e9:	data_out=16'h8a00;
17'h112ea:	data_out=16'h94b;
17'h112eb:	data_out=16'h9ed;
17'h112ec:	data_out=16'h894c;
17'h112ed:	data_out=16'h83f9;
17'h112ee:	data_out=16'h94c;
17'h112ef:	data_out=16'h9fb;
17'h112f0:	data_out=16'h95b;
17'h112f1:	data_out=16'h23e;
17'h112f2:	data_out=16'h7c4;
17'h112f3:	data_out=16'h881;
17'h112f4:	data_out=16'ha00;
17'h112f5:	data_out=16'h8a00;
17'h112f6:	data_out=16'h8983;
17'h112f7:	data_out=16'h93b;
17'h112f8:	data_out=16'h800d;
17'h112f9:	data_out=16'h59f;
17'h112fa:	data_out=16'h515;
17'h112fb:	data_out=16'h9c9;
17'h112fc:	data_out=16'h89fb;
17'h112fd:	data_out=16'h9e8;
17'h112fe:	data_out=16'h2b;
17'h112ff:	data_out=16'h89f1;
17'h11300:	data_out=16'h89ef;
17'h11301:	data_out=16'h89e9;
17'h11302:	data_out=16'h8202;
17'h11303:	data_out=16'h627;
17'h11304:	data_out=16'ha00;
17'h11305:	data_out=16'h9ef;
17'h11306:	data_out=16'h89d8;
17'h11307:	data_out=16'h9fe;
17'h11308:	data_out=16'h89d4;
17'h11309:	data_out=16'h24c;
17'h1130a:	data_out=16'h392;
17'h1130b:	data_out=16'h8612;
17'h1130c:	data_out=16'h72f;
17'h1130d:	data_out=16'h89eb;
17'h1130e:	data_out=16'h9e7;
17'h1130f:	data_out=16'h87af;
17'h11310:	data_out=16'h40;
17'h11311:	data_out=16'h884c;
17'h11312:	data_out=16'h8a00;
17'h11313:	data_out=16'h9d5;
17'h11314:	data_out=16'h223;
17'h11315:	data_out=16'h9f6;
17'h11316:	data_out=16'h9f5;
17'h11317:	data_out=16'h586;
17'h11318:	data_out=16'h89ff;
17'h11319:	data_out=16'ha00;
17'h1131a:	data_out=16'h9f5;
17'h1131b:	data_out=16'h9f4;
17'h1131c:	data_out=16'h89dd;
17'h1131d:	data_out=16'h86d2;
17'h1131e:	data_out=16'h816d;
17'h1131f:	data_out=16'h4fc;
17'h11320:	data_out=16'h883b;
17'h11321:	data_out=16'h9ec;
17'h11322:	data_out=16'h893a;
17'h11323:	data_out=16'h9f5;
17'h11324:	data_out=16'h9f6;
17'h11325:	data_out=16'h60b;
17'h11326:	data_out=16'h86d2;
17'h11327:	data_out=16'h9d5;
17'h11328:	data_out=16'h9f0;
17'h11329:	data_out=16'h9bf;
17'h1132a:	data_out=16'h84cb;
17'h1132b:	data_out=16'h9e2;
17'h1132c:	data_out=16'h9f5;
17'h1132d:	data_out=16'h89e7;
17'h1132e:	data_out=16'h86ea;
17'h1132f:	data_out=16'h4fd;
17'h11330:	data_out=16'ha00;
17'h11331:	data_out=16'h9dd;
17'h11332:	data_out=16'ha00;
17'h11333:	data_out=16'h89cc;
17'h11334:	data_out=16'h89c6;
17'h11335:	data_out=16'h9e4;
17'h11336:	data_out=16'h87c0;
17'h11337:	data_out=16'h679;
17'h11338:	data_out=16'h8a00;
17'h11339:	data_out=16'h89de;
17'h1133a:	data_out=16'h460;
17'h1133b:	data_out=16'ha00;
17'h1133c:	data_out=16'h9a6;
17'h1133d:	data_out=16'h81cf;
17'h1133e:	data_out=16'h9f0;
17'h1133f:	data_out=16'h9ee;
17'h11340:	data_out=16'ha00;
17'h11341:	data_out=16'h6b6;
17'h11342:	data_out=16'h89e4;
17'h11343:	data_out=16'h9f5;
17'h11344:	data_out=16'h9e7;
17'h11345:	data_out=16'h9f6;
17'h11346:	data_out=16'h8a00;
17'h11347:	data_out=16'h89e5;
17'h11348:	data_out=16'h855f;
17'h11349:	data_out=16'h9e6;
17'h1134a:	data_out=16'ha00;
17'h1134b:	data_out=16'h89d7;
17'h1134c:	data_out=16'h89fe;
17'h1134d:	data_out=16'h88df;
17'h1134e:	data_out=16'h5c5;
17'h1134f:	data_out=16'h855d;
17'h11350:	data_out=16'h9fc;
17'h11351:	data_out=16'h5bf;
17'h11352:	data_out=16'h9f8;
17'h11353:	data_out=16'h9fa;
17'h11354:	data_out=16'h8985;
17'h11355:	data_out=16'h9e3;
17'h11356:	data_out=16'h3c4;
17'h11357:	data_out=16'h8553;
17'h11358:	data_out=16'h48b;
17'h11359:	data_out=16'h9e5;
17'h1135a:	data_out=16'h8707;
17'h1135b:	data_out=16'h9d2;
17'h1135c:	data_out=16'h3a5;
17'h1135d:	data_out=16'h9d6;
17'h1135e:	data_out=16'h9ff;
17'h1135f:	data_out=16'h89eb;
17'h11360:	data_out=16'h8489;
17'h11361:	data_out=16'h9eb;
17'h11362:	data_out=16'h9fc;
17'h11363:	data_out=16'h8747;
17'h11364:	data_out=16'h89f9;
17'h11365:	data_out=16'ha00;
17'h11366:	data_out=16'ha00;
17'h11367:	data_out=16'ha00;
17'h11368:	data_out=16'h9ef;
17'h11369:	data_out=16'h8a00;
17'h1136a:	data_out=16'h9e3;
17'h1136b:	data_out=16'h9ec;
17'h1136c:	data_out=16'h89c7;
17'h1136d:	data_out=16'h87c2;
17'h1136e:	data_out=16'h9e3;
17'h1136f:	data_out=16'ha00;
17'h11370:	data_out=16'h9e5;
17'h11371:	data_out=16'h85d3;
17'h11372:	data_out=16'h8282;
17'h11373:	data_out=16'h9a9;
17'h11374:	data_out=16'ha00;
17'h11375:	data_out=16'h89fe;
17'h11376:	data_out=16'ha00;
17'h11377:	data_out=16'h9e3;
17'h11378:	data_out=16'hf5;
17'h11379:	data_out=16'h67e;
17'h1137a:	data_out=16'h8096;
17'h1137b:	data_out=16'h9f0;
17'h1137c:	data_out=16'h89ff;
17'h1137d:	data_out=16'h9fa;
17'h1137e:	data_out=16'h89ce;
17'h1137f:	data_out=16'h89f9;
17'h11380:	data_out=16'h89f5;
17'h11381:	data_out=16'h89fb;
17'h11382:	data_out=16'h80af;
17'h11383:	data_out=16'h3f5;
17'h11384:	data_out=16'ha00;
17'h11385:	data_out=16'ha00;
17'h11386:	data_out=16'h89ce;
17'h11387:	data_out=16'h9d7;
17'h11388:	data_out=16'h89de;
17'h11389:	data_out=16'h851c;
17'h1138a:	data_out=16'h81ea;
17'h1138b:	data_out=16'h8745;
17'h1138c:	data_out=16'h984;
17'h1138d:	data_out=16'h89f1;
17'h1138e:	data_out=16'h9f9;
17'h1138f:	data_out=16'h85d7;
17'h11390:	data_out=16'h44;
17'h11391:	data_out=16'h8649;
17'h11392:	data_out=16'h8a00;
17'h11393:	data_out=16'h8865;
17'h11394:	data_out=16'h81fa;
17'h11395:	data_out=16'h410;
17'h11396:	data_out=16'h85b;
17'h11397:	data_out=16'h111;
17'h11398:	data_out=16'h89ff;
17'h11399:	data_out=16'ha00;
17'h1139a:	data_out=16'ha00;
17'h1139b:	data_out=16'h6fa;
17'h1139c:	data_out=16'h87d5;
17'h1139d:	data_out=16'h89f0;
17'h1139e:	data_out=16'h8527;
17'h1139f:	data_out=16'h8243;
17'h113a0:	data_out=16'h88a0;
17'h113a1:	data_out=16'h9fb;
17'h113a2:	data_out=16'h840e;
17'h113a3:	data_out=16'h9cf;
17'h113a4:	data_out=16'h9d2;
17'h113a5:	data_out=16'h2e2;
17'h113a6:	data_out=16'h860c;
17'h113a7:	data_out=16'h5c7;
17'h113a8:	data_out=16'h9fc;
17'h113a9:	data_out=16'h9f4;
17'h113aa:	data_out=16'h83c4;
17'h113ab:	data_out=16'h9ff;
17'h113ac:	data_out=16'h53d;
17'h113ad:	data_out=16'h8a00;
17'h113ae:	data_out=16'h86a3;
17'h113af:	data_out=16'h8014;
17'h113b0:	data_out=16'ha00;
17'h113b1:	data_out=16'h55a;
17'h113b2:	data_out=16'ha00;
17'h113b3:	data_out=16'h8992;
17'h113b4:	data_out=16'h8a00;
17'h113b5:	data_out=16'h9cf;
17'h113b6:	data_out=16'h854b;
17'h113b7:	data_out=16'h635;
17'h113b8:	data_out=16'h8a00;
17'h113b9:	data_out=16'h89c9;
17'h113ba:	data_out=16'h8441;
17'h113bb:	data_out=16'ha00;
17'h113bc:	data_out=16'h9fb;
17'h113bd:	data_out=16'h83be;
17'h113be:	data_out=16'h9fc;
17'h113bf:	data_out=16'ha00;
17'h113c0:	data_out=16'ha00;
17'h113c1:	data_out=16'h98e;
17'h113c2:	data_out=16'h8a00;
17'h113c3:	data_out=16'h9fe;
17'h113c4:	data_out=16'h9fe;
17'h113c5:	data_out=16'h711;
17'h113c6:	data_out=16'h8a00;
17'h113c7:	data_out=16'h89f2;
17'h113c8:	data_out=16'h89c4;
17'h113c9:	data_out=16'h757;
17'h113ca:	data_out=16'h9ff;
17'h113cb:	data_out=16'h8a00;
17'h113cc:	data_out=16'h8921;
17'h113cd:	data_out=16'h8480;
17'h113ce:	data_out=16'h3b1;
17'h113cf:	data_out=16'h87e7;
17'h113d0:	data_out=16'ha00;
17'h113d1:	data_out=16'h8b9;
17'h113d2:	data_out=16'h9fb;
17'h113d3:	data_out=16'h9f0;
17'h113d4:	data_out=16'h889d;
17'h113d5:	data_out=16'h9fb;
17'h113d6:	data_out=16'h9af;
17'h113d7:	data_out=16'h85f4;
17'h113d8:	data_out=16'h737;
17'h113d9:	data_out=16'h809d;
17'h113da:	data_out=16'h89c4;
17'h113db:	data_out=16'h9fd;
17'h113dc:	data_out=16'h8000;
17'h113dd:	data_out=16'h4bb;
17'h113de:	data_out=16'h486;
17'h113df:	data_out=16'h89f0;
17'h113e0:	data_out=16'h87f8;
17'h113e1:	data_out=16'h9f2;
17'h113e2:	data_out=16'h8ac;
17'h113e3:	data_out=16'h8950;
17'h113e4:	data_out=16'h8a00;
17'h113e5:	data_out=16'ha00;
17'h113e6:	data_out=16'ha00;
17'h113e7:	data_out=16'ha00;
17'h113e8:	data_out=16'h9fb;
17'h113e9:	data_out=16'h8a00;
17'h113ea:	data_out=16'h9f6;
17'h113eb:	data_out=16'h9e5;
17'h113ec:	data_out=16'h88c2;
17'h113ed:	data_out=16'h8959;
17'h113ee:	data_out=16'h9f6;
17'h113ef:	data_out=16'ha00;
17'h113f0:	data_out=16'h9f8;
17'h113f1:	data_out=16'h8715;
17'h113f2:	data_out=16'h86b5;
17'h113f3:	data_out=16'h28f;
17'h113f4:	data_out=16'ha00;
17'h113f5:	data_out=16'h8237;
17'h113f6:	data_out=16'ha00;
17'h113f7:	data_out=16'h410;
17'h113f8:	data_out=16'h984;
17'h113f9:	data_out=16'h8cf;
17'h113fa:	data_out=16'h8436;
17'h113fb:	data_out=16'h9fd;
17'h113fc:	data_out=16'h89fe;
17'h113fd:	data_out=16'h8225;
17'h113fe:	data_out=16'h89dd;
17'h113ff:	data_out=16'h89f8;
17'h11400:	data_out=16'h8981;
17'h11401:	data_out=16'h89f9;
17'h11402:	data_out=16'h89bc;
17'h11403:	data_out=16'h87b2;
17'h11404:	data_out=16'ha00;
17'h11405:	data_out=16'ha00;
17'h11406:	data_out=16'h89dd;
17'h11407:	data_out=16'h9db;
17'h11408:	data_out=16'h89eb;
17'h11409:	data_out=16'h88ec;
17'h1140a:	data_out=16'h9d1;
17'h1140b:	data_out=16'h897b;
17'h1140c:	data_out=16'h9e6;
17'h1140d:	data_out=16'h89f8;
17'h1140e:	data_out=16'h9fd;
17'h1140f:	data_out=16'h8903;
17'h11410:	data_out=16'h86e2;
17'h11411:	data_out=16'h478;
17'h11412:	data_out=16'h89fd;
17'h11413:	data_out=16'h89d8;
17'h11414:	data_out=16'h88fa;
17'h11415:	data_out=16'h9f4;
17'h11416:	data_out=16'h57;
17'h11417:	data_out=16'h8928;
17'h11418:	data_out=16'h89ff;
17'h11419:	data_out=16'ha00;
17'h1141a:	data_out=16'ha00;
17'h1141b:	data_out=16'h88cb;
17'h1141c:	data_out=16'h89de;
17'h1141d:	data_out=16'h89ef;
17'h1141e:	data_out=16'h88e6;
17'h1141f:	data_out=16'h877c;
17'h11420:	data_out=16'h88b7;
17'h11421:	data_out=16'h9fd;
17'h11422:	data_out=16'h8776;
17'h11423:	data_out=16'h9e8;
17'h11424:	data_out=16'h9ea;
17'h11425:	data_out=16'h82e6;
17'h11426:	data_out=16'h8977;
17'h11427:	data_out=16'h237;
17'h11428:	data_out=16'h9fe;
17'h11429:	data_out=16'h9ee;
17'h1142a:	data_out=16'h880b;
17'h1142b:	data_out=16'ha00;
17'h1142c:	data_out=16'h1ea;
17'h1142d:	data_out=16'h8a00;
17'h1142e:	data_out=16'h88c2;
17'h1142f:	data_out=16'h8706;
17'h11430:	data_out=16'ha00;
17'h11431:	data_out=16'h9c8;
17'h11432:	data_out=16'ha00;
17'h11433:	data_out=16'h89cd;
17'h11434:	data_out=16'h8a00;
17'h11435:	data_out=16'h9dc;
17'h11436:	data_out=16'h8811;
17'h11437:	data_out=16'h89a3;
17'h11438:	data_out=16'h8a00;
17'h11439:	data_out=16'h89d9;
17'h1143a:	data_out=16'h8701;
17'h1143b:	data_out=16'ha00;
17'h1143c:	data_out=16'h815d;
17'h1143d:	data_out=16'h84d2;
17'h1143e:	data_out=16'h9fe;
17'h1143f:	data_out=16'ha00;
17'h11440:	data_out=16'ha00;
17'h11441:	data_out=16'h5f5;
17'h11442:	data_out=16'h8a00;
17'h11443:	data_out=16'ha00;
17'h11444:	data_out=16'ha00;
17'h11445:	data_out=16'h9f3;
17'h11446:	data_out=16'h8a00;
17'h11447:	data_out=16'h89de;
17'h11448:	data_out=16'h89dc;
17'h11449:	data_out=16'h12e;
17'h1144a:	data_out=16'h9f8;
17'h1144b:	data_out=16'h89fd;
17'h1144c:	data_out=16'h89bc;
17'h1144d:	data_out=16'h874b;
17'h1144e:	data_out=16'h85a7;
17'h1144f:	data_out=16'h8836;
17'h11450:	data_out=16'h336;
17'h11451:	data_out=16'h264;
17'h11452:	data_out=16'h9f7;
17'h11453:	data_out=16'h864d;
17'h11454:	data_out=16'h896c;
17'h11455:	data_out=16'h84d4;
17'h11456:	data_out=16'h9f6;
17'h11457:	data_out=16'h85af;
17'h11458:	data_out=16'h38;
17'h11459:	data_out=16'h9b8;
17'h1145a:	data_out=16'h89e5;
17'h1145b:	data_out=16'ha00;
17'h1145c:	data_out=16'h8988;
17'h1145d:	data_out=16'h82d7;
17'h1145e:	data_out=16'h85c8;
17'h1145f:	data_out=16'h89ea;
17'h11460:	data_out=16'h89d8;
17'h11461:	data_out=16'h9f4;
17'h11462:	data_out=16'h8662;
17'h11463:	data_out=16'h89be;
17'h11464:	data_out=16'h89fe;
17'h11465:	data_out=16'ha00;
17'h11466:	data_out=16'ha00;
17'h11467:	data_out=16'ha00;
17'h11468:	data_out=16'h9fd;
17'h11469:	data_out=16'h89fe;
17'h1146a:	data_out=16'h9fb;
17'h1146b:	data_out=16'h5c7;
17'h1146c:	data_out=16'h881b;
17'h1146d:	data_out=16'h89c5;
17'h1146e:	data_out=16'h9fb;
17'h1146f:	data_out=16'ha00;
17'h11470:	data_out=16'h9fd;
17'h11471:	data_out=16'h890b;
17'h11472:	data_out=16'h8647;
17'h11473:	data_out=16'h8107;
17'h11474:	data_out=16'ha00;
17'h11475:	data_out=16'h889a;
17'h11476:	data_out=16'ha00;
17'h11477:	data_out=16'h8574;
17'h11478:	data_out=16'h9c2;
17'h11479:	data_out=16'h968;
17'h1147a:	data_out=16'h8967;
17'h1147b:	data_out=16'h9fe;
17'h1147c:	data_out=16'h89ff;
17'h1147d:	data_out=16'h850d;
17'h1147e:	data_out=16'h89fa;
17'h1147f:	data_out=16'h815b;
17'h11480:	data_out=16'h8949;
17'h11481:	data_out=16'h89fc;
17'h11482:	data_out=16'h89e6;
17'h11483:	data_out=16'h89f6;
17'h11484:	data_out=16'ha00;
17'h11485:	data_out=16'ha00;
17'h11486:	data_out=16'h89fc;
17'h11487:	data_out=16'h99f;
17'h11488:	data_out=16'h89f9;
17'h11489:	data_out=16'h89f0;
17'h1148a:	data_out=16'h9f9;
17'h1148b:	data_out=16'h89b6;
17'h1148c:	data_out=16'h813;
17'h1148d:	data_out=16'h89fc;
17'h1148e:	data_out=16'h7ee;
17'h1148f:	data_out=16'h89d8;
17'h11490:	data_out=16'h89f2;
17'h11491:	data_out=16'h9e0;
17'h11492:	data_out=16'h89fe;
17'h11493:	data_out=16'h89fb;
17'h11494:	data_out=16'h89f1;
17'h11495:	data_out=16'h9f1;
17'h11496:	data_out=16'h87d1;
17'h11497:	data_out=16'h89f2;
17'h11498:	data_out=16'h89fb;
17'h11499:	data_out=16'ha00;
17'h1149a:	data_out=16'ha00;
17'h1149b:	data_out=16'h89ea;
17'h1149c:	data_out=16'h89fa;
17'h1149d:	data_out=16'h8845;
17'h1149e:	data_out=16'h89ef;
17'h1149f:	data_out=16'h88f1;
17'h114a0:	data_out=16'h897b;
17'h114a1:	data_out=16'h7a4;
17'h114a2:	data_out=16'h88cf;
17'h114a3:	data_out=16'h9e7;
17'h114a4:	data_out=16'h9e9;
17'h114a5:	data_out=16'h8764;
17'h114a6:	data_out=16'h89b1;
17'h114a7:	data_out=16'h6f4;
17'h114a8:	data_out=16'h794;
17'h114a9:	data_out=16'h99e;
17'h114aa:	data_out=16'h89ca;
17'h114ab:	data_out=16'ha00;
17'h114ac:	data_out=16'h86f5;
17'h114ad:	data_out=16'h8a00;
17'h114ae:	data_out=16'h89d4;
17'h114af:	data_out=16'h89f1;
17'h114b0:	data_out=16'h9fd;
17'h114b1:	data_out=16'h9ea;
17'h114b2:	data_out=16'h9f8;
17'h114b3:	data_out=16'h89f1;
17'h114b4:	data_out=16'h8a00;
17'h114b5:	data_out=16'h9e5;
17'h114b6:	data_out=16'h89c1;
17'h114b7:	data_out=16'h89da;
17'h114b8:	data_out=16'h89f7;
17'h114b9:	data_out=16'h89f5;
17'h114ba:	data_out=16'h89d9;
17'h114bb:	data_out=16'ha00;
17'h114bc:	data_out=16'h89db;
17'h114bd:	data_out=16'h851c;
17'h114be:	data_out=16'h795;
17'h114bf:	data_out=16'ha00;
17'h114c0:	data_out=16'ha00;
17'h114c1:	data_out=16'h88ee;
17'h114c2:	data_out=16'h8a00;
17'h114c3:	data_out=16'ha00;
17'h114c4:	data_out=16'ha00;
17'h114c5:	data_out=16'h9ef;
17'h114c6:	data_out=16'h8a00;
17'h114c7:	data_out=16'h89fa;
17'h114c8:	data_out=16'h89f9;
17'h114c9:	data_out=16'h8415;
17'h114ca:	data_out=16'h33e;
17'h114cb:	data_out=16'h89ff;
17'h114cc:	data_out=16'h89e4;
17'h114cd:	data_out=16'h8448;
17'h114ce:	data_out=16'h859c;
17'h114cf:	data_out=16'h89f2;
17'h114d0:	data_out=16'h8372;
17'h114d1:	data_out=16'h89ec;
17'h114d2:	data_out=16'h9f7;
17'h114d3:	data_out=16'h8435;
17'h114d4:	data_out=16'h89e5;
17'h114d5:	data_out=16'h89b8;
17'h114d6:	data_out=16'h9f1;
17'h114d7:	data_out=16'h86c4;
17'h114d8:	data_out=16'h89fd;
17'h114d9:	data_out=16'h9bf;
17'h114da:	data_out=16'h89ff;
17'h114db:	data_out=16'ha00;
17'h114dc:	data_out=16'h84d2;
17'h114dd:	data_out=16'h8917;
17'h114de:	data_out=16'h89f4;
17'h114df:	data_out=16'h89fd;
17'h114e0:	data_out=16'h89e5;
17'h114e1:	data_out=16'ha00;
17'h114e2:	data_out=16'h89e8;
17'h114e3:	data_out=16'h89ef;
17'h114e4:	data_out=16'h89f8;
17'h114e5:	data_out=16'h9f4;
17'h114e6:	data_out=16'ha00;
17'h114e7:	data_out=16'ha00;
17'h114e8:	data_out=16'h78b;
17'h114e9:	data_out=16'h89ff;
17'h114ea:	data_out=16'h801;
17'h114eb:	data_out=16'h7aa;
17'h114ec:	data_out=16'h87ae;
17'h114ed:	data_out=16'h89f0;
17'h114ee:	data_out=16'h801;
17'h114ef:	data_out=16'h9fd;
17'h114f0:	data_out=16'h7fb;
17'h114f1:	data_out=16'h89d1;
17'h114f2:	data_out=16'h7e7;
17'h114f3:	data_out=16'ha00;
17'h114f4:	data_out=16'h9fa;
17'h114f5:	data_out=16'h33c;
17'h114f6:	data_out=16'ha00;
17'h114f7:	data_out=16'h89ed;
17'h114f8:	data_out=16'h9eb;
17'h114f9:	data_out=16'h24e;
17'h114fa:	data_out=16'h89f2;
17'h114fb:	data_out=16'h793;
17'h114fc:	data_out=16'h89fa;
17'h114fd:	data_out=16'h8536;
17'h114fe:	data_out=16'h8a00;
17'h114ff:	data_out=16'h81b;
17'h11500:	data_out=16'h9d9;
17'h11501:	data_out=16'h933;
17'h11502:	data_out=16'h89fc;
17'h11503:	data_out=16'h89fb;
17'h11504:	data_out=16'ha00;
17'h11505:	data_out=16'ha00;
17'h11506:	data_out=16'h89ff;
17'h11507:	data_out=16'h1d3;
17'h11508:	data_out=16'h89fd;
17'h11509:	data_out=16'h89fc;
17'h1150a:	data_out=16'h9ff;
17'h1150b:	data_out=16'h89ed;
17'h1150c:	data_out=16'h8114;
17'h1150d:	data_out=16'h89ff;
17'h1150e:	data_out=16'h9ff;
17'h1150f:	data_out=16'h89fd;
17'h11510:	data_out=16'h88e8;
17'h11511:	data_out=16'h9ff;
17'h11512:	data_out=16'h8a00;
17'h11513:	data_out=16'h89fd;
17'h11514:	data_out=16'h89fc;
17'h11515:	data_out=16'h9fe;
17'h11516:	data_out=16'h8022;
17'h11517:	data_out=16'h89fe;
17'h11518:	data_out=16'h89fc;
17'h11519:	data_out=16'ha00;
17'h1151a:	data_out=16'ha00;
17'h1151b:	data_out=16'h89fd;
17'h1151c:	data_out=16'h39f;
17'h1151d:	data_out=16'h800;
17'h1151e:	data_out=16'h89f9;
17'h1151f:	data_out=16'h89e2;
17'h11520:	data_out=16'h9e2;
17'h11521:	data_out=16'h9ff;
17'h11522:	data_out=16'ha00;
17'h11523:	data_out=16'h9c5;
17'h11524:	data_out=16'h9c6;
17'h11525:	data_out=16'h845b;
17'h11526:	data_out=16'h89f3;
17'h11527:	data_out=16'h9e0;
17'h11528:	data_out=16'h9f7;
17'h11529:	data_out=16'h780;
17'h1152a:	data_out=16'h89fd;
17'h1152b:	data_out=16'ha00;
17'h1152c:	data_out=16'h596;
17'h1152d:	data_out=16'h8a00;
17'h1152e:	data_out=16'h89ff;
17'h1152f:	data_out=16'h89fa;
17'h11530:	data_out=16'h9f8;
17'h11531:	data_out=16'h9f4;
17'h11532:	data_out=16'h9f7;
17'h11533:	data_out=16'h89fb;
17'h11534:	data_out=16'h3e0;
17'h11535:	data_out=16'ha00;
17'h11536:	data_out=16'h89f2;
17'h11537:	data_out=16'h89fc;
17'h11538:	data_out=16'h289;
17'h11539:	data_out=16'h89fa;
17'h1153a:	data_out=16'h89d7;
17'h1153b:	data_out=16'ha00;
17'h1153c:	data_out=16'h8813;
17'h1153d:	data_out=16'h9f8;
17'h1153e:	data_out=16'h9f6;
17'h1153f:	data_out=16'ha00;
17'h11540:	data_out=16'ha00;
17'h11541:	data_out=16'h89bc;
17'h11542:	data_out=16'h8a00;
17'h11543:	data_out=16'h8321;
17'h11544:	data_out=16'ha00;
17'h11545:	data_out=16'h9fc;
17'h11546:	data_out=16'h8a00;
17'h11547:	data_out=16'h89f3;
17'h11548:	data_out=16'h89ff;
17'h11549:	data_out=16'h3a;
17'h1154a:	data_out=16'h8932;
17'h1154b:	data_out=16'h89ff;
17'h1154c:	data_out=16'h89ad;
17'h1154d:	data_out=16'ha00;
17'h1154e:	data_out=16'h8578;
17'h1154f:	data_out=16'h8716;
17'h11550:	data_out=16'h708;
17'h11551:	data_out=16'h89fb;
17'h11552:	data_out=16'h9fb;
17'h11553:	data_out=16'h80cd;
17'h11554:	data_out=16'h867f;
17'h11555:	data_out=16'h89f3;
17'h11556:	data_out=16'h9eb;
17'h11557:	data_out=16'h9fb;
17'h11558:	data_out=16'h89fe;
17'h11559:	data_out=16'ha00;
17'h1155a:	data_out=16'h8a00;
17'h1155b:	data_out=16'ha00;
17'h1155c:	data_out=16'h8c9;
17'h1155d:	data_out=16'h838e;
17'h1155e:	data_out=16'h89fb;
17'h1155f:	data_out=16'h89f7;
17'h11560:	data_out=16'h8a00;
17'h11561:	data_out=16'ha00;
17'h11562:	data_out=16'h89fc;
17'h11563:	data_out=16'h89fc;
17'h11564:	data_out=16'h83f1;
17'h11565:	data_out=16'h9d7;
17'h11566:	data_out=16'ha00;
17'h11567:	data_out=16'ha00;
17'h11568:	data_out=16'h9f8;
17'h11569:	data_out=16'h8a00;
17'h1156a:	data_out=16'h9ff;
17'h1156b:	data_out=16'h9cc;
17'h1156c:	data_out=16'h3cb;
17'h1156d:	data_out=16'h89fb;
17'h1156e:	data_out=16'h9ff;
17'h1156f:	data_out=16'h9ee;
17'h11570:	data_out=16'h9ff;
17'h11571:	data_out=16'h89fd;
17'h11572:	data_out=16'h9d5;
17'h11573:	data_out=16'ha00;
17'h11574:	data_out=16'h9f5;
17'h11575:	data_out=16'h8f2;
17'h11576:	data_out=16'ha00;
17'h11577:	data_out=16'h89e5;
17'h11578:	data_out=16'h706;
17'h11579:	data_out=16'h839e;
17'h1157a:	data_out=16'h89fc;
17'h1157b:	data_out=16'h9f6;
17'h1157c:	data_out=16'h89fb;
17'h1157d:	data_out=16'h84c2;
17'h1157e:	data_out=16'h8a00;
17'h1157f:	data_out=16'ha00;
17'h11580:	data_out=16'ha00;
17'h11581:	data_out=16'h9f8;
17'h11582:	data_out=16'h89fd;
17'h11583:	data_out=16'h89ed;
17'h11584:	data_out=16'ha00;
17'h11585:	data_out=16'h9fd;
17'h11586:	data_out=16'h8a00;
17'h11587:	data_out=16'h8891;
17'h11588:	data_out=16'h89fd;
17'h11589:	data_out=16'h8fa;
17'h1158a:	data_out=16'ha00;
17'h1158b:	data_out=16'h89fb;
17'h1158c:	data_out=16'h8a00;
17'h1158d:	data_out=16'h89ff;
17'h1158e:	data_out=16'ha00;
17'h1158f:	data_out=16'h89fe;
17'h11590:	data_out=16'h9e3;
17'h11591:	data_out=16'ha00;
17'h11592:	data_out=16'h89fe;
17'h11593:	data_out=16'h859f;
17'h11594:	data_out=16'h89fd;
17'h11595:	data_out=16'ha00;
17'h11596:	data_out=16'h9f3;
17'h11597:	data_out=16'h8a00;
17'h11598:	data_out=16'h11b;
17'h11599:	data_out=16'ha00;
17'h1159a:	data_out=16'ha00;
17'h1159b:	data_out=16'h8a00;
17'h1159c:	data_out=16'h910;
17'h1159d:	data_out=16'h9c1;
17'h1159e:	data_out=16'h86ec;
17'h1159f:	data_out=16'h83ec;
17'h115a0:	data_out=16'ha00;
17'h115a1:	data_out=16'h9ff;
17'h115a2:	data_out=16'ha00;
17'h115a3:	data_out=16'h989;
17'h115a4:	data_out=16'h987;
17'h115a5:	data_out=16'h9fd;
17'h115a6:	data_out=16'h89fd;
17'h115a7:	data_out=16'ha00;
17'h115a8:	data_out=16'h9ff;
17'h115a9:	data_out=16'h502;
17'h115aa:	data_out=16'h89fd;
17'h115ab:	data_out=16'ha00;
17'h115ac:	data_out=16'h9ff;
17'h115ad:	data_out=16'h8a00;
17'h115ae:	data_out=16'h8a00;
17'h115af:	data_out=16'h1a9;
17'h115b0:	data_out=16'h9f9;
17'h115b1:	data_out=16'ha00;
17'h115b2:	data_out=16'h9ef;
17'h115b3:	data_out=16'h89f7;
17'h115b4:	data_out=16'h7c4;
17'h115b5:	data_out=16'ha00;
17'h115b6:	data_out=16'h89e4;
17'h115b7:	data_out=16'h89fe;
17'h115b8:	data_out=16'h9fe;
17'h115b9:	data_out=16'h88bc;
17'h115ba:	data_out=16'h81c;
17'h115bb:	data_out=16'h992;
17'h115bc:	data_out=16'h89ee;
17'h115bd:	data_out=16'ha00;
17'h115be:	data_out=16'h9ff;
17'h115bf:	data_out=16'h9fd;
17'h115c0:	data_out=16'ha00;
17'h115c1:	data_out=16'h89fb;
17'h115c2:	data_out=16'h8a00;
17'h115c3:	data_out=16'h86ed;
17'h115c4:	data_out=16'ha00;
17'h115c5:	data_out=16'ha00;
17'h115c6:	data_out=16'h8a00;
17'h115c7:	data_out=16'h8281;
17'h115c8:	data_out=16'h8a00;
17'h115c9:	data_out=16'ha00;
17'h115ca:	data_out=16'h89fe;
17'h115cb:	data_out=16'h8a00;
17'h115cc:	data_out=16'h817c;
17'h115cd:	data_out=16'ha00;
17'h115ce:	data_out=16'h8332;
17'h115cf:	data_out=16'h87a;
17'h115d0:	data_out=16'h9f3;
17'h115d1:	data_out=16'h89fe;
17'h115d2:	data_out=16'h9ff;
17'h115d3:	data_out=16'h853c;
17'h115d4:	data_out=16'ha00;
17'h115d5:	data_out=16'h89fe;
17'h115d6:	data_out=16'h9f5;
17'h115d7:	data_out=16'ha00;
17'h115d8:	data_out=16'h8a00;
17'h115d9:	data_out=16'ha00;
17'h115da:	data_out=16'h8a00;
17'h115db:	data_out=16'ha00;
17'h115dc:	data_out=16'h8c8;
17'h115dd:	data_out=16'h9fb;
17'h115de:	data_out=16'he3;
17'h115df:	data_out=16'h3b8;
17'h115e0:	data_out=16'h89fe;
17'h115e1:	data_out=16'ha00;
17'h115e2:	data_out=16'h89ff;
17'h115e3:	data_out=16'h89fe;
17'h115e4:	data_out=16'ha00;
17'h115e5:	data_out=16'h9e7;
17'h115e6:	data_out=16'ha00;
17'h115e7:	data_out=16'ha00;
17'h115e8:	data_out=16'h9ff;
17'h115e9:	data_out=16'h89fe;
17'h115ea:	data_out=16'ha00;
17'h115eb:	data_out=16'ha00;
17'h115ec:	data_out=16'ha00;
17'h115ed:	data_out=16'h89fc;
17'h115ee:	data_out=16'ha00;
17'h115ef:	data_out=16'h268;
17'h115f0:	data_out=16'ha00;
17'h115f1:	data_out=16'h89fe;
17'h115f2:	data_out=16'ha00;
17'h115f3:	data_out=16'ha00;
17'h115f4:	data_out=16'h9db;
17'h115f5:	data_out=16'h89da;
17'h115f6:	data_out=16'ha00;
17'h115f7:	data_out=16'h951;
17'h115f8:	data_out=16'h8110;
17'h115f9:	data_out=16'h8495;
17'h115fa:	data_out=16'h89ff;
17'h115fb:	data_out=16'h9ff;
17'h115fc:	data_out=16'h15b;
17'h115fd:	data_out=16'h19b;
17'h115fe:	data_out=16'h23a;
17'h115ff:	data_out=16'ha00;
17'h11600:	data_out=16'ha00;
17'h11601:	data_out=16'h9fd;
17'h11602:	data_out=16'h89ff;
17'h11603:	data_out=16'h9f6;
17'h11604:	data_out=16'ha00;
17'h11605:	data_out=16'h9fb;
17'h11606:	data_out=16'h80c0;
17'h11607:	data_out=16'h860a;
17'h11608:	data_out=16'h8982;
17'h11609:	data_out=16'h9e5;
17'h1160a:	data_out=16'ha00;
17'h1160b:	data_out=16'h8798;
17'h1160c:	data_out=16'h8a00;
17'h1160d:	data_out=16'h8a00;
17'h1160e:	data_out=16'h5ff;
17'h1160f:	data_out=16'h88fa;
17'h11610:	data_out=16'h9f7;
17'h11611:	data_out=16'ha00;
17'h11612:	data_out=16'h89f3;
17'h11613:	data_out=16'h9ff;
17'h11614:	data_out=16'h5b8;
17'h11615:	data_out=16'ha00;
17'h11616:	data_out=16'ha00;
17'h11617:	data_out=16'h8a00;
17'h11618:	data_out=16'h9ff;
17'h11619:	data_out=16'h8bd;
17'h1161a:	data_out=16'ha00;
17'h1161b:	data_out=16'h8a00;
17'h1161c:	data_out=16'h9fc;
17'h1161d:	data_out=16'h9fc;
17'h1161e:	data_out=16'h9fb;
17'h1161f:	data_out=16'h68a;
17'h11620:	data_out=16'ha00;
17'h11621:	data_out=16'h588;
17'h11622:	data_out=16'ha00;
17'h11623:	data_out=16'h670;
17'h11624:	data_out=16'h67d;
17'h11625:	data_out=16'ha00;
17'h11626:	data_out=16'h873;
17'h11627:	data_out=16'h9ff;
17'h11628:	data_out=16'h4e6;
17'h11629:	data_out=16'h968;
17'h1162a:	data_out=16'h81ff;
17'h1162b:	data_out=16'ha00;
17'h1162c:	data_out=16'ha00;
17'h1162d:	data_out=16'h3ca;
17'h1162e:	data_out=16'h8953;
17'h1162f:	data_out=16'h9f6;
17'h11630:	data_out=16'h9c8;
17'h11631:	data_out=16'ha00;
17'h11632:	data_out=16'h982;
17'h11633:	data_out=16'h9f0;
17'h11634:	data_out=16'h9f6;
17'h11635:	data_out=16'ha00;
17'h11636:	data_out=16'h9f1;
17'h11637:	data_out=16'h8a00;
17'h11638:	data_out=16'ha00;
17'h11639:	data_out=16'h9f9;
17'h1163a:	data_out=16'h9f9;
17'h1163b:	data_out=16'h826;
17'h1163c:	data_out=16'h8a00;
17'h1163d:	data_out=16'ha00;
17'h1163e:	data_out=16'h4e1;
17'h1163f:	data_out=16'h9fb;
17'h11640:	data_out=16'ha00;
17'h11641:	data_out=16'h894d;
17'h11642:	data_out=16'h8706;
17'h11643:	data_out=16'h852a;
17'h11644:	data_out=16'ha00;
17'h11645:	data_out=16'ha00;
17'h11646:	data_out=16'h8a00;
17'h11647:	data_out=16'h9f7;
17'h11648:	data_out=16'h80f0;
17'h11649:	data_out=16'ha00;
17'h1164a:	data_out=16'h88ab;
17'h1164b:	data_out=16'h8a00;
17'h1164c:	data_out=16'h54e;
17'h1164d:	data_out=16'ha00;
17'h1164e:	data_out=16'h818e;
17'h1164f:	data_out=16'h9fd;
17'h11650:	data_out=16'h9fe;
17'h11651:	data_out=16'h82;
17'h11652:	data_out=16'ha00;
17'h11653:	data_out=16'h87fc;
17'h11654:	data_out=16'ha00;
17'h11655:	data_out=16'h89ff;
17'h11656:	data_out=16'h9fd;
17'h11657:	data_out=16'ha00;
17'h11658:	data_out=16'h8a00;
17'h11659:	data_out=16'ha00;
17'h1165a:	data_out=16'h8a00;
17'h1165b:	data_out=16'ha00;
17'h1165c:	data_out=16'h7d8;
17'h1165d:	data_out=16'ha00;
17'h1165e:	data_out=16'h9f4;
17'h1165f:	data_out=16'ha00;
17'h11660:	data_out=16'h81b0;
17'h11661:	data_out=16'h9ff;
17'h11662:	data_out=16'h8977;
17'h11663:	data_out=16'h9e8;
17'h11664:	data_out=16'ha00;
17'h11665:	data_out=16'h9e6;
17'h11666:	data_out=16'h9cf;
17'h11667:	data_out=16'ha00;
17'h11668:	data_out=16'h54e;
17'h11669:	data_out=16'h89ff;
17'h1166a:	data_out=16'h650;
17'h1166b:	data_out=16'ha00;
17'h1166c:	data_out=16'ha00;
17'h1166d:	data_out=16'h9ea;
17'h1166e:	data_out=16'h64e;
17'h1166f:	data_out=16'h808;
17'h11670:	data_out=16'h61c;
17'h11671:	data_out=16'h89ff;
17'h11672:	data_out=16'ha00;
17'h11673:	data_out=16'ha00;
17'h11674:	data_out=16'h938;
17'h11675:	data_out=16'h89fb;
17'h11676:	data_out=16'ha00;
17'h11677:	data_out=16'h9f5;
17'h11678:	data_out=16'h8485;
17'h11679:	data_out=16'h812b;
17'h1167a:	data_out=16'h9ae;
17'h1167b:	data_out=16'h4dd;
17'h1167c:	data_out=16'h9ff;
17'h1167d:	data_out=16'h6cd;
17'h1167e:	data_out=16'h875;
17'h1167f:	data_out=16'ha00;
17'h11680:	data_out=16'ha00;
17'h11681:	data_out=16'ha00;
17'h11682:	data_out=16'h8a00;
17'h11683:	data_out=16'h9ff;
17'h11684:	data_out=16'ha00;
17'h11685:	data_out=16'h9f8;
17'h11686:	data_out=16'h9ea;
17'h11687:	data_out=16'h371;
17'h11688:	data_out=16'h8a00;
17'h11689:	data_out=16'h9fe;
17'h1168a:	data_out=16'ha00;
17'h1168b:	data_out=16'h84b1;
17'h1168c:	data_out=16'h8a00;
17'h1168d:	data_out=16'h315;
17'h1168e:	data_out=16'h50;
17'h1168f:	data_out=16'h8688;
17'h11690:	data_out=16'ha00;
17'h11691:	data_out=16'ha00;
17'h11692:	data_out=16'h8068;
17'h11693:	data_out=16'ha00;
17'h11694:	data_out=16'ha00;
17'h11695:	data_out=16'ha00;
17'h11696:	data_out=16'ha00;
17'h11697:	data_out=16'h972;
17'h11698:	data_out=16'h124;
17'h11699:	data_out=16'h506;
17'h1169a:	data_out=16'ha00;
17'h1169b:	data_out=16'h818e;
17'h1169c:	data_out=16'h9fe;
17'h1169d:	data_out=16'ha00;
17'h1169e:	data_out=16'ha00;
17'h1169f:	data_out=16'ha00;
17'h116a0:	data_out=16'ha00;
17'h116a1:	data_out=16'h3e;
17'h116a2:	data_out=16'h9fd;
17'h116a3:	data_out=16'h8a00;
17'h116a4:	data_out=16'h8a00;
17'h116a5:	data_out=16'ha00;
17'h116a6:	data_out=16'h4e1;
17'h116a7:	data_out=16'ha00;
17'h116a8:	data_out=16'h3c;
17'h116a9:	data_out=16'h9c3;
17'h116aa:	data_out=16'h8611;
17'h116ab:	data_out=16'ha00;
17'h116ac:	data_out=16'ha00;
17'h116ad:	data_out=16'h9ff;
17'h116ae:	data_out=16'h82fc;
17'h116af:	data_out=16'ha00;
17'h116b0:	data_out=16'h82be;
17'h116b1:	data_out=16'ha00;
17'h116b2:	data_out=16'h8074;
17'h116b3:	data_out=16'ha00;
17'h116b4:	data_out=16'ha00;
17'h116b5:	data_out=16'h12;
17'h116b6:	data_out=16'h82e0;
17'h116b7:	data_out=16'h8a00;
17'h116b8:	data_out=16'ha00;
17'h116b9:	data_out=16'ha00;
17'h116ba:	data_out=16'ha00;
17'h116bb:	data_out=16'h6b8;
17'h116bc:	data_out=16'h8a00;
17'h116bd:	data_out=16'ha00;
17'h116be:	data_out=16'h3c;
17'h116bf:	data_out=16'h9fa;
17'h116c0:	data_out=16'ha00;
17'h116c1:	data_out=16'h8884;
17'h116c2:	data_out=16'h894c;
17'h116c3:	data_out=16'ha00;
17'h116c4:	data_out=16'ha00;
17'h116c5:	data_out=16'ha00;
17'h116c6:	data_out=16'h8a00;
17'h116c7:	data_out=16'ha00;
17'h116c8:	data_out=16'h853;
17'h116c9:	data_out=16'ha00;
17'h116ca:	data_out=16'h78;
17'h116cb:	data_out=16'h8a00;
17'h116cc:	data_out=16'h74b;
17'h116cd:	data_out=16'h9fd;
17'h116ce:	data_out=16'h865e;
17'h116cf:	data_out=16'h9f9;
17'h116d0:	data_out=16'ha00;
17'h116d1:	data_out=16'h1dc;
17'h116d2:	data_out=16'h86c0;
17'h116d3:	data_out=16'h792;
17'h116d4:	data_out=16'ha00;
17'h116d5:	data_out=16'h8897;
17'h116d6:	data_out=16'h9f8;
17'h116d7:	data_out=16'ha00;
17'h116d8:	data_out=16'h8a00;
17'h116d9:	data_out=16'ha00;
17'h116da:	data_out=16'h8a00;
17'h116db:	data_out=16'ha00;
17'h116dc:	data_out=16'h8f4;
17'h116dd:	data_out=16'ha00;
17'h116de:	data_out=16'ha00;
17'h116df:	data_out=16'h633;
17'h116e0:	data_out=16'h8267;
17'h116e1:	data_out=16'h9fe;
17'h116e2:	data_out=16'h8710;
17'h116e3:	data_out=16'ha00;
17'h116e4:	data_out=16'ha00;
17'h116e5:	data_out=16'ha00;
17'h116e6:	data_out=16'h63c;
17'h116e7:	data_out=16'h9fe;
17'h116e8:	data_out=16'h40;
17'h116e9:	data_out=16'h8a00;
17'h116ea:	data_out=16'h5b;
17'h116eb:	data_out=16'ha00;
17'h116ec:	data_out=16'ha00;
17'h116ed:	data_out=16'ha00;
17'h116ee:	data_out=16'h5b;
17'h116ef:	data_out=16'h95c;
17'h116f0:	data_out=16'h51;
17'h116f1:	data_out=16'h8a00;
17'h116f2:	data_out=16'ha00;
17'h116f3:	data_out=16'ha00;
17'h116f4:	data_out=16'h83cb;
17'h116f5:	data_out=16'h8a00;
17'h116f6:	data_out=16'ha00;
17'h116f7:	data_out=16'h9fc;
17'h116f8:	data_out=16'h9fd;
17'h116f9:	data_out=16'h850c;
17'h116fa:	data_out=16'ha00;
17'h116fb:	data_out=16'h3a;
17'h116fc:	data_out=16'h107;
17'h116fd:	data_out=16'ha00;
17'h116fe:	data_out=16'h9fe;
17'h116ff:	data_out=16'ha00;
17'h11700:	data_out=16'h9a4;
17'h11701:	data_out=16'h480;
17'h11702:	data_out=16'h8019;
17'h11703:	data_out=16'h579;
17'h11704:	data_out=16'h2e7;
17'h11705:	data_out=16'h366;
17'h11706:	data_out=16'h20f;
17'h11707:	data_out=16'h3c3;
17'h11708:	data_out=16'h810e;
17'h11709:	data_out=16'h875;
17'h1170a:	data_out=16'h470;
17'h1170b:	data_out=16'hf9;
17'h1170c:	data_out=16'h8758;
17'h1170d:	data_out=16'h1e2;
17'h1170e:	data_out=16'hc0;
17'h1170f:	data_out=16'h1c4;
17'h11710:	data_out=16'h54f;
17'h11711:	data_out=16'h4aa;
17'h11712:	data_out=16'h2d3;
17'h11713:	data_out=16'h54c;
17'h11714:	data_out=16'h489;
17'h11715:	data_out=16'h355;
17'h11716:	data_out=16'h269;
17'h11717:	data_out=16'h345;
17'h11718:	data_out=16'h146;
17'h11719:	data_out=16'h1a2;
17'h1171a:	data_out=16'h218;
17'h1171b:	data_out=16'h2f4;
17'h1171c:	data_out=16'h79b;
17'h1171d:	data_out=16'h614;
17'h1171e:	data_out=16'h501;
17'h1171f:	data_out=16'h443;
17'h11720:	data_out=16'ha00;
17'h11721:	data_out=16'hd0;
17'h11722:	data_out=16'h7e6;
17'h11723:	data_out=16'h8301;
17'h11724:	data_out=16'h8302;
17'h11725:	data_out=16'h43b;
17'h11726:	data_out=16'h462;
17'h11727:	data_out=16'h5a1;
17'h11728:	data_out=16'he3;
17'h11729:	data_out=16'h699;
17'h1172a:	data_out=16'h243;
17'h1172b:	data_out=16'h88c;
17'h1172c:	data_out=16'h2f3;
17'h1172d:	data_out=16'h213;
17'h1172e:	data_out=16'h1f9;
17'h1172f:	data_out=16'h5c5;
17'h11730:	data_out=16'h810e;
17'h11731:	data_out=16'h81e;
17'h11732:	data_out=16'h80aa;
17'h11733:	data_out=16'h5d1;
17'h11734:	data_out=16'h7a3;
17'h11735:	data_out=16'h825a;
17'h11736:	data_out=16'h802d;
17'h11737:	data_out=16'hcc;
17'h11738:	data_out=16'ha00;
17'h11739:	data_out=16'h5be;
17'h1173a:	data_out=16'h6fb;
17'h1173b:	data_out=16'h290;
17'h1173c:	data_out=16'h82dd;
17'h1173d:	data_out=16'ha00;
17'h1173e:	data_out=16'hf0;
17'h1173f:	data_out=16'h2ff;
17'h11740:	data_out=16'h50b;
17'h11741:	data_out=16'h8253;
17'h11742:	data_out=16'h8316;
17'h11743:	data_out=16'h1d7;
17'h11744:	data_out=16'h583;
17'h11745:	data_out=16'h35c;
17'h11746:	data_out=16'hac;
17'h11747:	data_out=16'h5e2;
17'h11748:	data_out=16'h446;
17'h11749:	data_out=16'h4a8;
17'h1174a:	data_out=16'hd1;
17'h1174b:	data_out=16'h8732;
17'h1174c:	data_out=16'h1f5;
17'h1174d:	data_out=16'h7e8;
17'h1174e:	data_out=16'h20c;
17'h1174f:	data_out=16'h1d2;
17'h11750:	data_out=16'h519;
17'h11751:	data_out=16'h803e;
17'h11752:	data_out=16'h8115;
17'h11753:	data_out=16'h593;
17'h11754:	data_out=16'h7b2;
17'h11755:	data_out=16'h83db;
17'h11756:	data_out=16'h67e;
17'h11757:	data_out=16'h725;
17'h11758:	data_out=16'h8468;
17'h11759:	data_out=16'h4de;
17'h1175a:	data_out=16'h80c6;
17'h1175b:	data_out=16'h381;
17'h1175c:	data_out=16'h22c;
17'h1175d:	data_out=16'h39a;
17'h1175e:	data_out=16'h5b1;
17'h1175f:	data_out=16'h24e;
17'h11760:	data_out=16'h37f;
17'h11761:	data_out=16'h615;
17'h11762:	data_out=16'h80fb;
17'h11763:	data_out=16'h582;
17'h11764:	data_out=16'ha00;
17'h11765:	data_out=16'h40f;
17'h11766:	data_out=16'h20a;
17'h11767:	data_out=16'h47f;
17'h11768:	data_out=16'hcd;
17'h11769:	data_out=16'h81a5;
17'h1176a:	data_out=16'hae;
17'h1176b:	data_out=16'h5e9;
17'h1176c:	data_out=16'h32c;
17'h1176d:	data_out=16'h5aa;
17'h1176e:	data_out=16'hb3;
17'h1176f:	data_out=16'h2f0;
17'h11770:	data_out=16'hba;
17'h11771:	data_out=16'hd0;
17'h11772:	data_out=16'h6a6;
17'h11773:	data_out=16'h806;
17'h11774:	data_out=16'h8164;
17'h11775:	data_out=16'h8394;
17'h11776:	data_out=16'h552;
17'h11777:	data_out=16'h529;
17'h11778:	data_out=16'h201;
17'h11779:	data_out=16'h179;
17'h1177a:	data_out=16'h4d7;
17'h1177b:	data_out=16'hea;
17'h1177c:	data_out=16'h10d;
17'h1177d:	data_out=16'h219;
17'h1177e:	data_out=16'h940;
17'h1177f:	data_out=16'h3e5;
17'h11780:	data_out=16'h90;
17'h11781:	data_out=16'h2b;
17'h11782:	data_out=16'h809a;
17'h11783:	data_out=16'h8a;
17'h11784:	data_out=16'h8037;
17'h11785:	data_out=16'h4e;
17'h11786:	data_out=16'ha;
17'h11787:	data_out=16'h8007;
17'h11788:	data_out=16'h8070;
17'h11789:	data_out=16'h8032;
17'h1178a:	data_out=16'h8004;
17'h1178b:	data_out=16'h8019;
17'h1178c:	data_out=16'h8082;
17'h1178d:	data_out=16'hd5;
17'h1178e:	data_out=16'h801a;
17'h1178f:	data_out=16'h34;
17'h11790:	data_out=16'h807f;
17'h11791:	data_out=16'h806e;
17'h11792:	data_out=16'h802a;
17'h11793:	data_out=16'hcc;
17'h11794:	data_out=16'h75;
17'h11795:	data_out=16'hc4;
17'h11796:	data_out=16'h10a;
17'h11797:	data_out=16'h81;
17'h11798:	data_out=16'h8037;
17'h11799:	data_out=16'h808c;
17'h1179a:	data_out=16'h7;
17'h1179b:	data_out=16'h57;
17'h1179c:	data_out=16'ha2;
17'h1179d:	data_out=16'h8059;
17'h1179e:	data_out=16'h63;
17'h1179f:	data_out=16'h9;
17'h117a0:	data_out=16'h44;
17'h117a1:	data_out=16'h801b;
17'h117a2:	data_out=16'h8022;
17'h117a3:	data_out=16'h80d8;
17'h117a4:	data_out=16'h80e0;
17'h117a5:	data_out=16'h8066;
17'h117a6:	data_out=16'h8031;
17'h117a7:	data_out=16'h8067;
17'h117a8:	data_out=16'h800e;
17'h117a9:	data_out=16'h7d;
17'h117aa:	data_out=16'h8044;
17'h117ab:	data_out=16'h8068;
17'h117ac:	data_out=16'h8b;
17'h117ad:	data_out=16'h8070;
17'h117ae:	data_out=16'h807b;
17'h117af:	data_out=16'h75;
17'h117b0:	data_out=16'h4f;
17'h117b1:	data_out=16'h84;
17'h117b2:	data_out=16'h4f;
17'h117b3:	data_out=16'h82;
17'h117b4:	data_out=16'h9;
17'h117b5:	data_out=16'h808a;
17'h117b6:	data_out=16'h8081;
17'h117b7:	data_out=16'h806f;
17'h117b8:	data_out=16'h8012;
17'h117b9:	data_out=16'h78;
17'h117ba:	data_out=16'h806d;
17'h117bb:	data_out=16'hb;
17'h117bc:	data_out=16'h804d;
17'h117bd:	data_out=16'h59;
17'h117be:	data_out=16'h8009;
17'h117bf:	data_out=16'h48;
17'h117c0:	data_out=16'h8049;
17'h117c1:	data_out=16'h8023;
17'h117c2:	data_out=16'h8051;
17'h117c3:	data_out=16'h10;
17'h117c4:	data_out=16'h2b;
17'h117c5:	data_out=16'hce;
17'h117c6:	data_out=16'h8088;
17'h117c7:	data_out=16'h8059;
17'h117c8:	data_out=16'h8057;
17'h117c9:	data_out=16'h8065;
17'h117ca:	data_out=16'h8076;
17'h117cb:	data_out=16'h8070;
17'h117cc:	data_out=16'h8082;
17'h117cd:	data_out=16'h13;
17'h117ce:	data_out=16'h8034;
17'h117cf:	data_out=16'h8086;
17'h117d0:	data_out=16'h6;
17'h117d1:	data_out=16'hf2;
17'h117d2:	data_out=16'h809f;
17'h117d3:	data_out=16'h8025;
17'h117d4:	data_out=16'h8;
17'h117d5:	data_out=16'h8003;
17'h117d6:	data_out=16'h802f;
17'h117d7:	data_out=16'h8076;
17'h117d8:	data_out=16'h804f;
17'h117d9:	data_out=16'h806c;
17'h117da:	data_out=16'h8050;
17'h117db:	data_out=16'h14;
17'h117dc:	data_out=16'h23;
17'h117dd:	data_out=16'h14;
17'h117de:	data_out=16'h4c;
17'h117df:	data_out=16'h8018;
17'h117e0:	data_out=16'h804f;
17'h117e1:	data_out=16'h52;
17'h117e2:	data_out=16'h3f;
17'h117e3:	data_out=16'h6c;
17'h117e4:	data_out=16'h8018;
17'h117e5:	data_out=16'h8063;
17'h117e6:	data_out=16'h806f;
17'h117e7:	data_out=16'h8059;
17'h117e8:	data_out=16'h800e;
17'h117e9:	data_out=16'h8089;
17'h117ea:	data_out=16'h8015;
17'h117eb:	data_out=16'h66;
17'h117ec:	data_out=16'h4f;
17'h117ed:	data_out=16'h7d;
17'h117ee:	data_out=16'h800d;
17'h117ef:	data_out=16'hbe;
17'h117f0:	data_out=16'h8018;
17'h117f1:	data_out=16'h804b;
17'h117f2:	data_out=16'h8b;
17'h117f3:	data_out=16'h9b;
17'h117f4:	data_out=16'h4b;
17'h117f5:	data_out=16'h2a;
17'h117f6:	data_out=16'h8046;
17'h117f7:	data_out=16'h803d;
17'h117f8:	data_out=16'h4a;
17'h117f9:	data_out=16'h8074;
17'h117fa:	data_out=16'h77;
17'h117fb:	data_out=16'h800b;
17'h117fc:	data_out=16'h8022;
17'h117fd:	data_out=16'h28;
17'h117fe:	data_out=16'h8014;
17'h117ff:	data_out=16'h8023;
17'h11800:	data_out=16'h8007;
17'h11801:	data_out=16'h8008;
17'h11802:	data_out=16'h7;
17'h11803:	data_out=16'h8003;
17'h11804:	data_out=16'h2;
17'h11805:	data_out=16'h6;
17'h11806:	data_out=16'h8008;
17'h11807:	data_out=16'h8002;
17'h11808:	data_out=16'h8001;
17'h11809:	data_out=16'h2;
17'h1180a:	data_out=16'h7;
17'h1180b:	data_out=16'h7;
17'h1180c:	data_out=16'h5;
17'h1180d:	data_out=16'h6;
17'h1180e:	data_out=16'h3;
17'h1180f:	data_out=16'h8008;
17'h11810:	data_out=16'h8006;
17'h11811:	data_out=16'h8004;
17'h11812:	data_out=16'h8006;
17'h11813:	data_out=16'h8008;
17'h11814:	data_out=16'h8003;
17'h11815:	data_out=16'h8008;
17'h11816:	data_out=16'h4;
17'h11817:	data_out=16'h8001;
17'h11818:	data_out=16'h8007;
17'h11819:	data_out=16'h2;
17'h1181a:	data_out=16'h8002;
17'h1181b:	data_out=16'h8004;
17'h1181c:	data_out=16'h3;
17'h1181d:	data_out=16'h6;
17'h1181e:	data_out=16'h1;
17'h1181f:	data_out=16'h6;
17'h11820:	data_out=16'h7;
17'h11821:	data_out=16'h8001;
17'h11822:	data_out=16'h8006;
17'h11823:	data_out=16'h8000;
17'h11824:	data_out=16'h8004;
17'h11825:	data_out=16'h8004;
17'h11826:	data_out=16'h7;
17'h11827:	data_out=16'h4;
17'h11828:	data_out=16'h7;
17'h11829:	data_out=16'h4;
17'h1182a:	data_out=16'h2;
17'h1182b:	data_out=16'h2;
17'h1182c:	data_out=16'h1;
17'h1182d:	data_out=16'h8004;
17'h1182e:	data_out=16'h4;
17'h1182f:	data_out=16'h4;
17'h11830:	data_out=16'h1;
17'h11831:	data_out=16'h7;
17'h11832:	data_out=16'h5;
17'h11833:	data_out=16'h7;
17'h11834:	data_out=16'h8;
17'h11835:	data_out=16'h1;
17'h11836:	data_out=16'h8002;
17'h11837:	data_out=16'h8008;
17'h11838:	data_out=16'h8006;
17'h11839:	data_out=16'h4;
17'h1183a:	data_out=16'h8004;
17'h1183b:	data_out=16'h6;
17'h1183c:	data_out=16'h1;
17'h1183d:	data_out=16'h6;
17'h1183e:	data_out=16'h3;
17'h1183f:	data_out=16'h8001;
17'h11840:	data_out=16'h8004;
17'h11841:	data_out=16'h6;
17'h11842:	data_out=16'h8;
17'h11843:	data_out=16'h0;
17'h11844:	data_out=16'h8007;
17'h11845:	data_out=16'h5;
17'h11846:	data_out=16'h8005;
17'h11847:	data_out=16'h9;
17'h11848:	data_out=16'h0;
17'h11849:	data_out=16'h6;
17'h1184a:	data_out=16'h2;
17'h1184b:	data_out=16'h8008;
17'h1184c:	data_out=16'h8006;
17'h1184d:	data_out=16'h8004;
17'h1184e:	data_out=16'h5;
17'h1184f:	data_out=16'h4;
17'h11850:	data_out=16'h8006;
17'h11851:	data_out=16'h2;
17'h11852:	data_out=16'h2;
17'h11853:	data_out=16'h8007;
17'h11854:	data_out=16'h8007;
17'h11855:	data_out=16'h9;
17'h11856:	data_out=16'h8006;
17'h11857:	data_out=16'h8004;
17'h11858:	data_out=16'h4;
17'h11859:	data_out=16'h8000;
17'h1185a:	data_out=16'h8007;
17'h1185b:	data_out=16'h8004;
17'h1185c:	data_out=16'h8003;
17'h1185d:	data_out=16'h5;
17'h1185e:	data_out=16'h4;
17'h1185f:	data_out=16'h1;
17'h11860:	data_out=16'h2;
17'h11861:	data_out=16'h3;
17'h11862:	data_out=16'h8007;
17'h11863:	data_out=16'h4;
17'h11864:	data_out=16'h8001;
17'h11865:	data_out=16'h8003;
17'h11866:	data_out=16'h4;
17'h11867:	data_out=16'h8;
17'h11868:	data_out=16'h8006;
17'h11869:	data_out=16'h8003;
17'h1186a:	data_out=16'h8009;
17'h1186b:	data_out=16'h8003;
17'h1186c:	data_out=16'h2;
17'h1186d:	data_out=16'h6;
17'h1186e:	data_out=16'h8009;
17'h1186f:	data_out=16'h5;
17'h11870:	data_out=16'h8002;
17'h11871:	data_out=16'h3;
17'h11872:	data_out=16'h8;
17'h11873:	data_out=16'h1;
17'h11874:	data_out=16'h2;
17'h11875:	data_out=16'h8007;
17'h11876:	data_out=16'h6;
17'h11877:	data_out=16'h8003;
17'h11878:	data_out=16'h1;
17'h11879:	data_out=16'h9;
17'h1187a:	data_out=16'h2;
17'h1187b:	data_out=16'h7;
17'h1187c:	data_out=16'h5;
17'h1187d:	data_out=16'h8003;
17'h1187e:	data_out=16'h8001;
17'h1187f:	data_out=16'h8002;
17'h11880:	data_out=16'h1aa;
17'h11881:	data_out=16'h96;
17'h11882:	data_out=16'h8060;
17'h11883:	data_out=16'h814e;
17'h11884:	data_out=16'h8004;
17'h11885:	data_out=16'h8196;
17'h11886:	data_out=16'h8170;
17'h11887:	data_out=16'h60;
17'h11888:	data_out=16'h158;
17'h11889:	data_out=16'hb7;
17'h1188a:	data_out=16'h289;
17'h1188b:	data_out=16'h32;
17'h1188c:	data_out=16'h30d;
17'h1188d:	data_out=16'h8186;
17'h1188e:	data_out=16'h8051;
17'h1188f:	data_out=16'h8173;
17'h11890:	data_out=16'h801a;
17'h11891:	data_out=16'hda;
17'h11892:	data_out=16'h80ce;
17'h11893:	data_out=16'h815d;
17'h11894:	data_out=16'h81b1;
17'h11895:	data_out=16'h80c3;
17'h11896:	data_out=16'h80d2;
17'h11897:	data_out=16'h819b;
17'h11898:	data_out=16'h804f;
17'h11899:	data_out=16'h179;
17'h1189a:	data_out=16'h8027;
17'h1189b:	data_out=16'h815d;
17'h1189c:	data_out=16'h820f;
17'h1189d:	data_out=16'h131;
17'h1189e:	data_out=16'h81e3;
17'h1189f:	data_out=16'h81db;
17'h118a0:	data_out=16'h8193;
17'h118a1:	data_out=16'h8054;
17'h118a2:	data_out=16'h8120;
17'h118a3:	data_out=16'h1e6;
17'h118a4:	data_out=16'h1db;
17'h118a5:	data_out=16'h59;
17'h118a6:	data_out=16'h292;
17'h118a7:	data_out=16'hcf;
17'h118a8:	data_out=16'h8050;
17'h118a9:	data_out=16'h810d;
17'h118aa:	data_out=16'h26;
17'h118ab:	data_out=16'h1ac;
17'h118ac:	data_out=16'h8057;
17'h118ad:	data_out=16'h1ee;
17'h118ae:	data_out=16'h8161;
17'h118af:	data_out=16'h815b;
17'h118b0:	data_out=16'h5;
17'h118b1:	data_out=16'h280;
17'h118b2:	data_out=16'h8020;
17'h118b3:	data_out=16'h81d2;
17'h118b4:	data_out=16'h201;
17'h118b5:	data_out=16'h174;
17'h118b6:	data_out=16'h12;
17'h118b7:	data_out=16'h80b4;
17'h118b8:	data_out=16'h8144;
17'h118b9:	data_out=16'h8193;
17'h118ba:	data_out=16'h27;
17'h118bb:	data_out=16'h201;
17'h118bc:	data_out=16'h4;
17'h118bd:	data_out=16'h8075;
17'h118be:	data_out=16'h8054;
17'h118bf:	data_out=16'h8159;
17'h118c0:	data_out=16'h81d4;
17'h118c1:	data_out=16'h80d9;
17'h118c2:	data_out=16'h1bc;
17'h118c3:	data_out=16'h8206;
17'h118c4:	data_out=16'h9a;
17'h118c5:	data_out=16'h80a8;
17'h118c6:	data_out=16'h8052;
17'h118c7:	data_out=16'h802b;
17'h118c8:	data_out=16'h8177;
17'h118c9:	data_out=16'h24;
17'h118ca:	data_out=16'h1e;
17'h118cb:	data_out=16'h328;
17'h118cc:	data_out=16'h8017;
17'h118cd:	data_out=16'h8137;
17'h118ce:	data_out=16'h802f;
17'h118cf:	data_out=16'h49;
17'h118d0:	data_out=16'h8217;
17'h118d1:	data_out=16'h8180;
17'h118d2:	data_out=16'h178;
17'h118d3:	data_out=16'h80ae;
17'h118d4:	data_out=16'h8129;
17'h118d5:	data_out=16'h808e;
17'h118d6:	data_out=16'h8101;
17'h118d7:	data_out=16'h812d;
17'h118d8:	data_out=16'h8009;
17'h118d9:	data_out=16'h8173;
17'h118da:	data_out=16'h8149;
17'h118db:	data_out=16'h8129;
17'h118dc:	data_out=16'ha;
17'h118dd:	data_out=16'h8100;
17'h118de:	data_out=16'h813c;
17'h118df:	data_out=16'h8076;
17'h118e0:	data_out=16'h298;
17'h118e1:	data_out=16'h80cb;
17'h118e2:	data_out=16'h8132;
17'h118e3:	data_out=16'h81bf;
17'h118e4:	data_out=16'h1bf;
17'h118e5:	data_out=16'hd4;
17'h118e6:	data_out=16'h14f;
17'h118e7:	data_out=16'h81a7;
17'h118e8:	data_out=16'h8057;
17'h118e9:	data_out=16'he8;
17'h118ea:	data_out=16'h8055;
17'h118eb:	data_out=16'h80ff;
17'h118ec:	data_out=16'h245;
17'h118ed:	data_out=16'h81d5;
17'h118ee:	data_out=16'h805b;
17'h118ef:	data_out=16'h81bd;
17'h118f0:	data_out=16'h804a;
17'h118f1:	data_out=16'h80e6;
17'h118f2:	data_out=16'h81d6;
17'h118f3:	data_out=16'h81be;
17'h118f4:	data_out=16'h4;
17'h118f5:	data_out=16'h8154;
17'h118f6:	data_out=16'h18b;
17'h118f7:	data_out=16'h80fe;
17'h118f8:	data_out=16'h8174;
17'h118f9:	data_out=16'h813e;
17'h118fa:	data_out=16'h81b5;
17'h118fb:	data_out=16'h8046;
17'h118fc:	data_out=16'h8088;
17'h118fd:	data_out=16'h81fd;
17'h118fe:	data_out=16'h8e;
17'h118ff:	data_out=16'h810f;
17'h11900:	data_out=16'h876c;
17'h11901:	data_out=16'h1d0;
17'h11902:	data_out=16'h475;
17'h11903:	data_out=16'h71;
17'h11904:	data_out=16'h2a0;
17'h11905:	data_out=16'h733;
17'h11906:	data_out=16'h4cb;
17'h11907:	data_out=16'h3b6;
17'h11908:	data_out=16'h4d5;
17'h11909:	data_out=16'h11;
17'h1190a:	data_out=16'h8097;
17'h1190b:	data_out=16'h50d;
17'h1190c:	data_out=16'h65f;
17'h1190d:	data_out=16'h8004;
17'h1190e:	data_out=16'h1ed;
17'h1190f:	data_out=16'h625;
17'h11910:	data_out=16'hb8;
17'h11911:	data_out=16'h509;
17'h11912:	data_out=16'h474;
17'h11913:	data_out=16'h6d;
17'h11914:	data_out=16'h3d4;
17'h11915:	data_out=16'h80c4;
17'h11916:	data_out=16'h1b;
17'h11917:	data_out=16'h2d5;
17'h11918:	data_out=16'h237;
17'h11919:	data_out=16'h4f0;
17'h1191a:	data_out=16'h308;
17'h1191b:	data_out=16'h46c;
17'h1191c:	data_out=16'h52f;
17'h1191d:	data_out=16'h352;
17'h1191e:	data_out=16'h4c4;
17'h1191f:	data_out=16'h778;
17'h11920:	data_out=16'h60c;
17'h11921:	data_out=16'h1f6;
17'h11922:	data_out=16'h810e;
17'h11923:	data_out=16'h123;
17'h11924:	data_out=16'h123;
17'h11925:	data_out=16'hee;
17'h11926:	data_out=16'h27;
17'h11927:	data_out=16'h4fb;
17'h11928:	data_out=16'h212;
17'h11929:	data_out=16'h839e;
17'h1192a:	data_out=16'h316;
17'h1192b:	data_out=16'h78e;
17'h1192c:	data_out=16'h30;
17'h1192d:	data_out=16'h893b;
17'h1192e:	data_out=16'h65f;
17'h1192f:	data_out=16'h4d5;
17'h11930:	data_out=16'h202;
17'h11931:	data_out=16'h29a;
17'h11932:	data_out=16'h1f2;
17'h11933:	data_out=16'h534;
17'h11934:	data_out=16'h28d;
17'h11935:	data_out=16'h9ff;
17'h11936:	data_out=16'h5b3;
17'h11937:	data_out=16'h4e2;
17'h11938:	data_out=16'h3d2;
17'h11939:	data_out=16'h541;
17'h1193a:	data_out=16'h804e;
17'h1193b:	data_out=16'h27e;
17'h1193c:	data_out=16'h35c;
17'h1193d:	data_out=16'h149;
17'h1193e:	data_out=16'h213;
17'h1193f:	data_out=16'h72f;
17'h11940:	data_out=16'h387;
17'h11941:	data_out=16'h718;
17'h11942:	data_out=16'h85dd;
17'h11943:	data_out=16'h43a;
17'h11944:	data_out=16'h25c;
17'h11945:	data_out=16'h80bc;
17'h11946:	data_out=16'h55;
17'h11947:	data_out=16'hac;
17'h11948:	data_out=16'h57e;
17'h11949:	data_out=16'hd7;
17'h1194a:	data_out=16'h5d9;
17'h1194b:	data_out=16'hf9;
17'h1194c:	data_out=16'h20;
17'h1194d:	data_out=16'h8109;
17'h1194e:	data_out=16'h602;
17'h1194f:	data_out=16'h90;
17'h11950:	data_out=16'h32f;
17'h11951:	data_out=16'h5ea;
17'h11952:	data_out=16'h15;
17'h11953:	data_out=16'h711;
17'h11954:	data_out=16'h453;
17'h11955:	data_out=16'h708;
17'h11956:	data_out=16'h278;
17'h11957:	data_out=16'h1c4;
17'h11958:	data_out=16'h574;
17'h11959:	data_out=16'h2ed;
17'h1195a:	data_out=16'h165;
17'h1195b:	data_out=16'h6ee;
17'h1195c:	data_out=16'h62c;
17'h1195d:	data_out=16'h74;
17'h1195e:	data_out=16'h46d;
17'h1195f:	data_out=16'h105;
17'h11960:	data_out=16'h81e0;
17'h11961:	data_out=16'h485;
17'h11962:	data_out=16'h2c7;
17'h11963:	data_out=16'h56d;
17'h11964:	data_out=16'h3a9;
17'h11965:	data_out=16'h41f;
17'h11966:	data_out=16'h668;
17'h11967:	data_out=16'h280;
17'h11968:	data_out=16'h1ff;
17'h11969:	data_out=16'h4b4;
17'h1196a:	data_out=16'h1e7;
17'h1196b:	data_out=16'h432;
17'h1196c:	data_out=16'h8952;
17'h1196d:	data_out=16'h55a;
17'h1196e:	data_out=16'h1e7;
17'h1196f:	data_out=16'h12d;
17'h11970:	data_out=16'h1eb;
17'h11971:	data_out=16'h7f1;
17'h11972:	data_out=16'hb9;
17'h11973:	data_out=16'h3b9;
17'h11974:	data_out=16'h1f6;
17'h11975:	data_out=16'h39f;
17'h11976:	data_out=16'h583;
17'h11977:	data_out=16'h178;
17'h11978:	data_out=16'h3b4;
17'h11979:	data_out=16'h80a;
17'h1197a:	data_out=16'h4a2;
17'h1197b:	data_out=16'h213;
17'h1197c:	data_out=16'h24f;
17'h1197d:	data_out=16'h76a;
17'h1197e:	data_out=16'h13b;
17'h1197f:	data_out=16'h336;
17'h11980:	data_out=16'h8a00;
17'h11981:	data_out=16'h519;
17'h11982:	data_out=16'h9fc;
17'h11983:	data_out=16'h262;
17'h11984:	data_out=16'ha00;
17'h11985:	data_out=16'ha00;
17'h11986:	data_out=16'h9f2;
17'h11987:	data_out=16'h87dd;
17'h11988:	data_out=16'h8331;
17'h11989:	data_out=16'h8a00;
17'h1198a:	data_out=16'h8a00;
17'h1198b:	data_out=16'h99d;
17'h1198c:	data_out=16'h196;
17'h1198d:	data_out=16'h3c6;
17'h1198e:	data_out=16'h4a4;
17'h1198f:	data_out=16'h8a2;
17'h11990:	data_out=16'h89fd;
17'h11991:	data_out=16'ha00;
17'h11992:	data_out=16'h7a4;
17'h11993:	data_out=16'h81b4;
17'h11994:	data_out=16'ha00;
17'h11995:	data_out=16'ha9;
17'h11996:	data_out=16'h8a00;
17'h11997:	data_out=16'h9f3;
17'h11998:	data_out=16'h1f6;
17'h11999:	data_out=16'ha00;
17'h1199a:	data_out=16'ha00;
17'h1199b:	data_out=16'ha00;
17'h1199c:	data_out=16'h9fa;
17'h1199d:	data_out=16'h994;
17'h1199e:	data_out=16'h9f3;
17'h1199f:	data_out=16'ha00;
17'h119a0:	data_out=16'ha00;
17'h119a1:	data_out=16'h50b;
17'h119a2:	data_out=16'h8a00;
17'h119a3:	data_out=16'h8a00;
17'h119a4:	data_out=16'h8a00;
17'h119a5:	data_out=16'h89ff;
17'h119a6:	data_out=16'h8a00;
17'h119a7:	data_out=16'ha00;
17'h119a8:	data_out=16'h619;
17'h119a9:	data_out=16'h8a00;
17'h119aa:	data_out=16'h8a00;
17'h119ab:	data_out=16'ha00;
17'h119ac:	data_out=16'h8952;
17'h119ad:	data_out=16'h8a00;
17'h119ae:	data_out=16'h591;
17'h119af:	data_out=16'ha00;
17'h119b0:	data_out=16'h89bf;
17'h119b1:	data_out=16'ha00;
17'h119b2:	data_out=16'h8800;
17'h119b3:	data_out=16'ha00;
17'h119b4:	data_out=16'h80d8;
17'h119b5:	data_out=16'h9fe;
17'h119b6:	data_out=16'h409;
17'h119b7:	data_out=16'h9fc;
17'h119b8:	data_out=16'ha00;
17'h119b9:	data_out=16'ha00;
17'h119ba:	data_out=16'h8a00;
17'h119bb:	data_out=16'h8f1;
17'h119bc:	data_out=16'h9fa;
17'h119bd:	data_out=16'h9e9;
17'h119be:	data_out=16'h623;
17'h119bf:	data_out=16'ha00;
17'h119c0:	data_out=16'h58e;
17'h119c1:	data_out=16'h9fa;
17'h119c2:	data_out=16'h8a00;
17'h119c3:	data_out=16'ha00;
17'h119c4:	data_out=16'ha00;
17'h119c5:	data_out=16'h39;
17'h119c6:	data_out=16'h89ff;
17'h119c7:	data_out=16'h8a00;
17'h119c8:	data_out=16'h9fe;
17'h119c9:	data_out=16'h8a00;
17'h119ca:	data_out=16'h79b;
17'h119cb:	data_out=16'h8a00;
17'h119cc:	data_out=16'h8a00;
17'h119cd:	data_out=16'h8a00;
17'h119ce:	data_out=16'h179;
17'h119cf:	data_out=16'h8a00;
17'h119d0:	data_out=16'h989;
17'h119d1:	data_out=16'h9f8;
17'h119d2:	data_out=16'h8a00;
17'h119d3:	data_out=16'ha00;
17'h119d4:	data_out=16'ha00;
17'h119d5:	data_out=16'h9e8;
17'h119d6:	data_out=16'h8a00;
17'h119d7:	data_out=16'h89ab;
17'h119d8:	data_out=16'ha00;
17'h119d9:	data_out=16'h869b;
17'h119da:	data_out=16'ha00;
17'h119db:	data_out=16'ha00;
17'h119dc:	data_out=16'ha00;
17'h119dd:	data_out=16'h89ff;
17'h119de:	data_out=16'ha00;
17'h119df:	data_out=16'h818f;
17'h119e0:	data_out=16'h8a00;
17'h119e1:	data_out=16'ha00;
17'h119e2:	data_out=16'h736;
17'h119e3:	data_out=16'ha00;
17'h119e4:	data_out=16'h3f5;
17'h119e5:	data_out=16'ha00;
17'h119e6:	data_out=16'ha00;
17'h119e7:	data_out=16'h83c2;
17'h119e8:	data_out=16'h560;
17'h119e9:	data_out=16'h8927;
17'h119ea:	data_out=16'h462;
17'h119eb:	data_out=16'ha00;
17'h119ec:	data_out=16'h8a00;
17'h119ed:	data_out=16'ha00;
17'h119ee:	data_out=16'h462;
17'h119ef:	data_out=16'h735;
17'h119f0:	data_out=16'h488;
17'h119f1:	data_out=16'h9f6;
17'h119f2:	data_out=16'h82b;
17'h119f3:	data_out=16'h9fb;
17'h119f4:	data_out=16'h89ff;
17'h119f5:	data_out=16'ha00;
17'h119f6:	data_out=16'ha00;
17'h119f7:	data_out=16'h81df;
17'h119f8:	data_out=16'ha00;
17'h119f9:	data_out=16'h187;
17'h119fa:	data_out=16'ha00;
17'h119fb:	data_out=16'h626;
17'h119fc:	data_out=16'h78b;
17'h119fd:	data_out=16'ha00;
17'h119fe:	data_out=16'h89fa;
17'h119ff:	data_out=16'h18b;
17'h11a00:	data_out=16'h89d3;
17'h11a01:	data_out=16'h9ef;
17'h11a02:	data_out=16'h9d6;
17'h11a03:	data_out=16'h8a00;
17'h11a04:	data_out=16'ha00;
17'h11a05:	data_out=16'h9ef;
17'h11a06:	data_out=16'h608;
17'h11a07:	data_out=16'h87c6;
17'h11a08:	data_out=16'h759;
17'h11a09:	data_out=16'h89fd;
17'h11a0a:	data_out=16'h742;
17'h11a0b:	data_out=16'h7b7;
17'h11a0c:	data_out=16'h8a00;
17'h11a0d:	data_out=16'h8a00;
17'h11a0e:	data_out=16'h9a4;
17'h11a0f:	data_out=16'h30e;
17'h11a10:	data_out=16'h89fa;
17'h11a11:	data_out=16'ha00;
17'h11a12:	data_out=16'h9e2;
17'h11a13:	data_out=16'h8403;
17'h11a14:	data_out=16'h9e6;
17'h11a15:	data_out=16'h9f5;
17'h11a16:	data_out=16'h8a00;
17'h11a17:	data_out=16'h4f4;
17'h11a18:	data_out=16'h3d9;
17'h11a19:	data_out=16'ha00;
17'h11a1a:	data_out=16'h9f2;
17'h11a1b:	data_out=16'h9e9;
17'h11a1c:	data_out=16'h9ad;
17'h11a1d:	data_out=16'h9f5;
17'h11a1e:	data_out=16'h9b0;
17'h11a1f:	data_out=16'h9fd;
17'h11a20:	data_out=16'ha00;
17'h11a21:	data_out=16'h9fe;
17'h11a22:	data_out=16'h89fd;
17'h11a23:	data_out=16'h83f3;
17'h11a24:	data_out=16'h83e7;
17'h11a25:	data_out=16'h89f2;
17'h11a26:	data_out=16'h8a00;
17'h11a27:	data_out=16'ha00;
17'h11a28:	data_out=16'h9ff;
17'h11a29:	data_out=16'h8a00;
17'h11a2a:	data_out=16'h89fc;
17'h11a2b:	data_out=16'ha00;
17'h11a2c:	data_out=16'h89ff;
17'h11a2d:	data_out=16'h8a00;
17'h11a2e:	data_out=16'h56;
17'h11a2f:	data_out=16'h9ed;
17'h11a30:	data_out=16'h839f;
17'h11a31:	data_out=16'h9ff;
17'h11a32:	data_out=16'h273;
17'h11a33:	data_out=16'h9f8;
17'h11a34:	data_out=16'h6ff;
17'h11a35:	data_out=16'h9ff;
17'h11a36:	data_out=16'h9ee;
17'h11a37:	data_out=16'h9da;
17'h11a38:	data_out=16'h9f9;
17'h11a39:	data_out=16'h9f5;
17'h11a3a:	data_out=16'h89fb;
17'h11a3b:	data_out=16'ha00;
17'h11a3c:	data_out=16'h9e8;
17'h11a3d:	data_out=16'h9df;
17'h11a3e:	data_out=16'h9ff;
17'h11a3f:	data_out=16'h9ef;
17'h11a40:	data_out=16'h9ea;
17'h11a41:	data_out=16'h9c0;
17'h11a42:	data_out=16'h8a00;
17'h11a43:	data_out=16'h9f3;
17'h11a44:	data_out=16'ha00;
17'h11a45:	data_out=16'h9bb;
17'h11a46:	data_out=16'h8999;
17'h11a47:	data_out=16'h89fc;
17'h11a48:	data_out=16'h9dc;
17'h11a49:	data_out=16'h89f9;
17'h11a4a:	data_out=16'ha00;
17'h11a4b:	data_out=16'h8a00;
17'h11a4c:	data_out=16'h8a00;
17'h11a4d:	data_out=16'h89fc;
17'h11a4e:	data_out=16'h261;
17'h11a4f:	data_out=16'h8a00;
17'h11a50:	data_out=16'h1cd;
17'h11a51:	data_out=16'h6c9;
17'h11a52:	data_out=16'h8a00;
17'h11a53:	data_out=16'ha00;
17'h11a54:	data_out=16'h9f4;
17'h11a55:	data_out=16'h3b6;
17'h11a56:	data_out=16'h9df;
17'h11a57:	data_out=16'h51c;
17'h11a58:	data_out=16'h9e1;
17'h11a59:	data_out=16'h82c;
17'h11a5a:	data_out=16'h9fe;
17'h11a5b:	data_out=16'ha00;
17'h11a5c:	data_out=16'h9fb;
17'h11a5d:	data_out=16'h89f9;
17'h11a5e:	data_out=16'h9e8;
17'h11a5f:	data_out=16'h81c9;
17'h11a60:	data_out=16'h8a00;
17'h11a61:	data_out=16'h9f1;
17'h11a62:	data_out=16'h8689;
17'h11a63:	data_out=16'h9f9;
17'h11a64:	data_out=16'h9ff;
17'h11a65:	data_out=16'h9ff;
17'h11a66:	data_out=16'ha00;
17'h11a67:	data_out=16'h8958;
17'h11a68:	data_out=16'h9fe;
17'h11a69:	data_out=16'h88d5;
17'h11a6a:	data_out=16'h94b;
17'h11a6b:	data_out=16'h9e7;
17'h11a6c:	data_out=16'h89f8;
17'h11a6d:	data_out=16'h9f8;
17'h11a6e:	data_out=16'h949;
17'h11a6f:	data_out=16'h83a5;
17'h11a70:	data_out=16'h97f;
17'h11a71:	data_out=16'h9b8;
17'h11a72:	data_out=16'h9ed;
17'h11a73:	data_out=16'h9ee;
17'h11a74:	data_out=16'h864f;
17'h11a75:	data_out=16'h9c2;
17'h11a76:	data_out=16'ha00;
17'h11a77:	data_out=16'h89fe;
17'h11a78:	data_out=16'h6e2;
17'h11a79:	data_out=16'h8407;
17'h11a7a:	data_out=16'h9f0;
17'h11a7b:	data_out=16'h9ff;
17'h11a7c:	data_out=16'h9ff;
17'h11a7d:	data_out=16'ha00;
17'h11a7e:	data_out=16'h8795;
17'h11a7f:	data_out=16'h837;
17'h11a80:	data_out=16'h89cb;
17'h11a81:	data_out=16'ha00;
17'h11a82:	data_out=16'h8da;
17'h11a83:	data_out=16'h89fe;
17'h11a84:	data_out=16'h9df;
17'h11a85:	data_out=16'h979;
17'h11a86:	data_out=16'h82c;
17'h11a87:	data_out=16'h89da;
17'h11a88:	data_out=16'ha00;
17'h11a89:	data_out=16'h89fa;
17'h11a8a:	data_out=16'h9ff;
17'h11a8b:	data_out=16'h9fc;
17'h11a8c:	data_out=16'h89f6;
17'h11a8d:	data_out=16'h8a00;
17'h11a8e:	data_out=16'h9fb;
17'h11a8f:	data_out=16'h89fb;
17'h11a90:	data_out=16'h89f8;
17'h11a91:	data_out=16'ha00;
17'h11a92:	data_out=16'h734;
17'h11a93:	data_out=16'h6b7;
17'h11a94:	data_out=16'h4ef;
17'h11a95:	data_out=16'h3d6;
17'h11a96:	data_out=16'h89ff;
17'h11a97:	data_out=16'h834a;
17'h11a98:	data_out=16'h85e2;
17'h11a99:	data_out=16'ha00;
17'h11a9a:	data_out=16'h9cf;
17'h11a9b:	data_out=16'h97d;
17'h11a9c:	data_out=16'h45d;
17'h11a9d:	data_out=16'ha00;
17'h11a9e:	data_out=16'h8430;
17'h11a9f:	data_out=16'h9fc;
17'h11aa0:	data_out=16'h9da;
17'h11aa1:	data_out=16'h9fb;
17'h11aa2:	data_out=16'h89fe;
17'h11aa3:	data_out=16'ha00;
17'h11aa4:	data_out=16'ha00;
17'h11aa5:	data_out=16'h89f9;
17'h11aa6:	data_out=16'h89d6;
17'h11aa7:	data_out=16'ha00;
17'h11aa8:	data_out=16'h9fb;
17'h11aa9:	data_out=16'h89ec;
17'h11aaa:	data_out=16'h89fb;
17'h11aab:	data_out=16'ha00;
17'h11aac:	data_out=16'h89fe;
17'h11aad:	data_out=16'h89d9;
17'h11aae:	data_out=16'h830c;
17'h11aaf:	data_out=16'h61f;
17'h11ab0:	data_out=16'h96d;
17'h11ab1:	data_out=16'ha00;
17'h11ab2:	data_out=16'h9f8;
17'h11ab3:	data_out=16'h9eb;
17'h11ab4:	data_out=16'ha00;
17'h11ab5:	data_out=16'ha00;
17'h11ab6:	data_out=16'h6d8;
17'h11ab7:	data_out=16'h9f4;
17'h11ab8:	data_out=16'h9e7;
17'h11ab9:	data_out=16'h9e0;
17'h11aba:	data_out=16'h89f8;
17'h11abb:	data_out=16'ha00;
17'h11abc:	data_out=16'h9f2;
17'h11abd:	data_out=16'h50f;
17'h11abe:	data_out=16'h9fb;
17'h11abf:	data_out=16'h95c;
17'h11ac0:	data_out=16'h9d0;
17'h11ac1:	data_out=16'h80a1;
17'h11ac2:	data_out=16'h8a00;
17'h11ac3:	data_out=16'h8853;
17'h11ac4:	data_out=16'ha00;
17'h11ac5:	data_out=16'h310;
17'h11ac6:	data_out=16'h9ee;
17'h11ac7:	data_out=16'h89f9;
17'h11ac8:	data_out=16'h86bf;
17'h11ac9:	data_out=16'h89f9;
17'h11aca:	data_out=16'ha00;
17'h11acb:	data_out=16'h8a00;
17'h11acc:	data_out=16'h8a00;
17'h11acd:	data_out=16'h89fe;
17'h11ace:	data_out=16'h3cf;
17'h11acf:	data_out=16'h8a00;
17'h11ad0:	data_out=16'h89fc;
17'h11ad1:	data_out=16'h8552;
17'h11ad2:	data_out=16'h1ae;
17'h11ad3:	data_out=16'ha00;
17'h11ad4:	data_out=16'h9d5;
17'h11ad5:	data_out=16'h8081;
17'h11ad6:	data_out=16'h9ee;
17'h11ad7:	data_out=16'h9c8;
17'h11ad8:	data_out=16'h9e7;
17'h11ad9:	data_out=16'h9bf;
17'h11ada:	data_out=16'h9fd;
17'h11adb:	data_out=16'ha00;
17'h11adc:	data_out=16'h9f8;
17'h11add:	data_out=16'h89fa;
17'h11ade:	data_out=16'h80e3;
17'h11adf:	data_out=16'h89e7;
17'h11ae0:	data_out=16'h89b9;
17'h11ae1:	data_out=16'h9eb;
17'h11ae2:	data_out=16'h89bc;
17'h11ae3:	data_out=16'h9f1;
17'h11ae4:	data_out=16'ha00;
17'h11ae5:	data_out=16'ha00;
17'h11ae6:	data_out=16'ha00;
17'h11ae7:	data_out=16'h89b7;
17'h11ae8:	data_out=16'h9fb;
17'h11ae9:	data_out=16'h22f;
17'h11aea:	data_out=16'h9fb;
17'h11aeb:	data_out=16'h914;
17'h11aec:	data_out=16'h89f3;
17'h11aed:	data_out=16'h9f0;
17'h11aee:	data_out=16'h9fb;
17'h11aef:	data_out=16'h652;
17'h11af0:	data_out=16'h9fb;
17'h11af1:	data_out=16'h158;
17'h11af2:	data_out=16'h9bc;
17'h11af3:	data_out=16'h9db;
17'h11af4:	data_out=16'h924;
17'h11af5:	data_out=16'h9bd;
17'h11af6:	data_out=16'ha00;
17'h11af7:	data_out=16'h89fd;
17'h11af8:	data_out=16'h89f9;
17'h11af9:	data_out=16'h89f6;
17'h11afa:	data_out=16'h9c7;
17'h11afb:	data_out=16'h9fb;
17'h11afc:	data_out=16'h92c;
17'h11afd:	data_out=16'h9dd;
17'h11afe:	data_out=16'h8466;
17'h11aff:	data_out=16'h89fd;
17'h11b00:	data_out=16'h89ba;
17'h11b01:	data_out=16'ha00;
17'h11b02:	data_out=16'h1e8;
17'h11b03:	data_out=16'h89fa;
17'h11b04:	data_out=16'h9e8;
17'h11b05:	data_out=16'h9cc;
17'h11b06:	data_out=16'h9b9;
17'h11b07:	data_out=16'h89df;
17'h11b08:	data_out=16'h8959;
17'h11b09:	data_out=16'h89fb;
17'h11b0a:	data_out=16'ha00;
17'h11b0b:	data_out=16'h724;
17'h11b0c:	data_out=16'h89f5;
17'h11b0d:	data_out=16'h8a00;
17'h11b0e:	data_out=16'h9f8;
17'h11b0f:	data_out=16'h89fd;
17'h11b10:	data_out=16'h89f9;
17'h11b11:	data_out=16'ha00;
17'h11b12:	data_out=16'h8696;
17'h11b13:	data_out=16'ha00;
17'h11b14:	data_out=16'h8631;
17'h11b15:	data_out=16'h18e;
17'h11b16:	data_out=16'h89fc;
17'h11b17:	data_out=16'h8973;
17'h11b18:	data_out=16'h89fe;
17'h11b19:	data_out=16'ha00;
17'h11b1a:	data_out=16'h9d3;
17'h11b1b:	data_out=16'h8739;
17'h11b1c:	data_out=16'hdc;
17'h11b1d:	data_out=16'ha00;
17'h11b1e:	data_out=16'h89c7;
17'h11b1f:	data_out=16'ha00;
17'h11b20:	data_out=16'h9d4;
17'h11b21:	data_out=16'h9f7;
17'h11b22:	data_out=16'h89fd;
17'h11b23:	data_out=16'ha00;
17'h11b24:	data_out=16'ha00;
17'h11b25:	data_out=16'h89ea;
17'h11b26:	data_out=16'h89d7;
17'h11b27:	data_out=16'ha00;
17'h11b28:	data_out=16'h9f8;
17'h11b29:	data_out=16'h89e8;
17'h11b2a:	data_out=16'h89e3;
17'h11b2b:	data_out=16'ha00;
17'h11b2c:	data_out=16'h89fc;
17'h11b2d:	data_out=16'h89bd;
17'h11b2e:	data_out=16'h858c;
17'h11b2f:	data_out=16'h823f;
17'h11b30:	data_out=16'h9fc;
17'h11b31:	data_out=16'ha00;
17'h11b32:	data_out=16'ha00;
17'h11b33:	data_out=16'h827f;
17'h11b34:	data_out=16'ha00;
17'h11b35:	data_out=16'h9ff;
17'h11b36:	data_out=16'h894e;
17'h11b37:	data_out=16'h902;
17'h11b38:	data_out=16'h9fe;
17'h11b39:	data_out=16'h89a6;
17'h11b3a:	data_out=16'h89fc;
17'h11b3b:	data_out=16'h9fe;
17'h11b3c:	data_out=16'h9fc;
17'h11b3d:	data_out=16'h804c;
17'h11b3e:	data_out=16'h9f8;
17'h11b3f:	data_out=16'h9c9;
17'h11b40:	data_out=16'h9d9;
17'h11b41:	data_out=16'h89ff;
17'h11b42:	data_out=16'h8a00;
17'h11b43:	data_out=16'h8154;
17'h11b44:	data_out=16'ha00;
17'h11b45:	data_out=16'hc7;
17'h11b46:	data_out=16'h9e9;
17'h11b47:	data_out=16'h89fe;
17'h11b48:	data_out=16'h898b;
17'h11b49:	data_out=16'h89f7;
17'h11b4a:	data_out=16'h85e9;
17'h11b4b:	data_out=16'h8a00;
17'h11b4c:	data_out=16'h8a00;
17'h11b4d:	data_out=16'h89fe;
17'h11b4e:	data_out=16'h834b;
17'h11b4f:	data_out=16'h8a00;
17'h11b50:	data_out=16'h89f9;
17'h11b51:	data_out=16'h89fd;
17'h11b52:	data_out=16'h336;
17'h11b53:	data_out=16'ha00;
17'h11b54:	data_out=16'h9cd;
17'h11b55:	data_out=16'h8999;
17'h11b56:	data_out=16'h9e3;
17'h11b57:	data_out=16'h9a5;
17'h11b58:	data_out=16'h8746;
17'h11b59:	data_out=16'h9be;
17'h11b5a:	data_out=16'h9f0;
17'h11b5b:	data_out=16'ha00;
17'h11b5c:	data_out=16'h9f9;
17'h11b5d:	data_out=16'h89f4;
17'h11b5e:	data_out=16'h87cb;
17'h11b5f:	data_out=16'h89f5;
17'h11b60:	data_out=16'h89b4;
17'h11b61:	data_out=16'h9f6;
17'h11b62:	data_out=16'h8902;
17'h11b63:	data_out=16'h7a8;
17'h11b64:	data_out=16'ha00;
17'h11b65:	data_out=16'ha00;
17'h11b66:	data_out=16'ha00;
17'h11b67:	data_out=16'h89d1;
17'h11b68:	data_out=16'h9f7;
17'h11b69:	data_out=16'h89ff;
17'h11b6a:	data_out=16'h9f8;
17'h11b6b:	data_out=16'h9cb;
17'h11b6c:	data_out=16'h89e0;
17'h11b6d:	data_out=16'h6f9;
17'h11b6e:	data_out=16'h9f8;
17'h11b6f:	data_out=16'h9d5;
17'h11b70:	data_out=16'h9f8;
17'h11b71:	data_out=16'h89ab;
17'h11b72:	data_out=16'h9c5;
17'h11b73:	data_out=16'h9f9;
17'h11b74:	data_out=16'h9ee;
17'h11b75:	data_out=16'h9ea;
17'h11b76:	data_out=16'h9fd;
17'h11b77:	data_out=16'h8a00;
17'h11b78:	data_out=16'h813c;
17'h11b79:	data_out=16'h8a00;
17'h11b7a:	data_out=16'h27e;
17'h11b7b:	data_out=16'h9f8;
17'h11b7c:	data_out=16'h89ed;
17'h11b7d:	data_out=16'h9e2;
17'h11b7e:	data_out=16'h75f;
17'h11b7f:	data_out=16'h89fe;
17'h11b80:	data_out=16'h896a;
17'h11b81:	data_out=16'ha00;
17'h11b82:	data_out=16'h8a00;
17'h11b83:	data_out=16'h89f9;
17'h11b84:	data_out=16'ha00;
17'h11b85:	data_out=16'h9d9;
17'h11b86:	data_out=16'h993;
17'h11b87:	data_out=16'h8a00;
17'h11b88:	data_out=16'h89fe;
17'h11b89:	data_out=16'h89fb;
17'h11b8a:	data_out=16'ha00;
17'h11b8b:	data_out=16'h89a2;
17'h11b8c:	data_out=16'h8a00;
17'h11b8d:	data_out=16'h8a00;
17'h11b8e:	data_out=16'h9f8;
17'h11b8f:	data_out=16'h8a00;
17'h11b90:	data_out=16'h89f6;
17'h11b91:	data_out=16'ha00;
17'h11b92:	data_out=16'h8a00;
17'h11b93:	data_out=16'ha00;
17'h11b94:	data_out=16'h89ec;
17'h11b95:	data_out=16'h8294;
17'h11b96:	data_out=16'h89f8;
17'h11b97:	data_out=16'h89e3;
17'h11b98:	data_out=16'h8a00;
17'h11b99:	data_out=16'h9ff;
17'h11b9a:	data_out=16'h9f2;
17'h11b9b:	data_out=16'h89ff;
17'h11b9c:	data_out=16'h8937;
17'h11b9d:	data_out=16'ha00;
17'h11b9e:	data_out=16'h89f7;
17'h11b9f:	data_out=16'h866a;
17'h11ba0:	data_out=16'h9db;
17'h11ba1:	data_out=16'h9f7;
17'h11ba2:	data_out=16'h89fa;
17'h11ba3:	data_out=16'ha00;
17'h11ba4:	data_out=16'ha00;
17'h11ba5:	data_out=16'h8992;
17'h11ba6:	data_out=16'h89e6;
17'h11ba7:	data_out=16'ha00;
17'h11ba8:	data_out=16'h9f7;
17'h11ba9:	data_out=16'h8a00;
17'h11baa:	data_out=16'h89d1;
17'h11bab:	data_out=16'h9fb;
17'h11bac:	data_out=16'h89ee;
17'h11bad:	data_out=16'h884e;
17'h11bae:	data_out=16'h88e4;
17'h11baf:	data_out=16'h88fe;
17'h11bb0:	data_out=16'h9f8;
17'h11bb1:	data_out=16'ha00;
17'h11bb2:	data_out=16'ha00;
17'h11bb3:	data_out=16'h89f7;
17'h11bb4:	data_out=16'ha00;
17'h11bb5:	data_out=16'h9fd;
17'h11bb6:	data_out=16'h89bc;
17'h11bb7:	data_out=16'h89bf;
17'h11bb8:	data_out=16'ha00;
17'h11bb9:	data_out=16'h89fc;
17'h11bba:	data_out=16'h89fc;
17'h11bbb:	data_out=16'h9f7;
17'h11bbc:	data_out=16'ha00;
17'h11bbd:	data_out=16'h880d;
17'h11bbe:	data_out=16'h9f7;
17'h11bbf:	data_out=16'h9d6;
17'h11bc0:	data_out=16'ha00;
17'h11bc1:	data_out=16'h8a00;
17'h11bc2:	data_out=16'h8a00;
17'h11bc3:	data_out=16'h3e4;
17'h11bc4:	data_out=16'ha00;
17'h11bc5:	data_out=16'h8383;
17'h11bc6:	data_out=16'h812;
17'h11bc7:	data_out=16'h8a00;
17'h11bc8:	data_out=16'h89aa;
17'h11bc9:	data_out=16'h89c8;
17'h11bca:	data_out=16'h8991;
17'h11bcb:	data_out=16'h8a00;
17'h11bcc:	data_out=16'h8a00;
17'h11bcd:	data_out=16'h89f8;
17'h11bce:	data_out=16'h89f1;
17'h11bcf:	data_out=16'h89ff;
17'h11bd0:	data_out=16'h89f4;
17'h11bd1:	data_out=16'h8a00;
17'h11bd2:	data_out=16'h73b;
17'h11bd3:	data_out=16'h9fc;
17'h11bd4:	data_out=16'h8018;
17'h11bd5:	data_out=16'h89fa;
17'h11bd6:	data_out=16'h97d;
17'h11bd7:	data_out=16'h6be;
17'h11bd8:	data_out=16'h8a00;
17'h11bd9:	data_out=16'h9f9;
17'h11bda:	data_out=16'h1a2;
17'h11bdb:	data_out=16'ha00;
17'h11bdc:	data_out=16'h9eb;
17'h11bdd:	data_out=16'h8974;
17'h11bde:	data_out=16'h8859;
17'h11bdf:	data_out=16'h89f1;
17'h11be0:	data_out=16'h89e4;
17'h11be1:	data_out=16'ha00;
17'h11be2:	data_out=16'h894a;
17'h11be3:	data_out=16'h89e8;
17'h11be4:	data_out=16'ha00;
17'h11be5:	data_out=16'ha00;
17'h11be6:	data_out=16'h9fa;
17'h11be7:	data_out=16'h89b7;
17'h11be8:	data_out=16'h9f7;
17'h11be9:	data_out=16'h8a00;
17'h11bea:	data_out=16'h9f9;
17'h11beb:	data_out=16'h9ef;
17'h11bec:	data_out=16'h896a;
17'h11bed:	data_out=16'h89eb;
17'h11bee:	data_out=16'h9f9;
17'h11bef:	data_out=16'ha00;
17'h11bf0:	data_out=16'h9f9;
17'h11bf1:	data_out=16'h89f0;
17'h11bf2:	data_out=16'h9fc;
17'h11bf3:	data_out=16'ha00;
17'h11bf4:	data_out=16'h9e8;
17'h11bf5:	data_out=16'h9e1;
17'h11bf6:	data_out=16'h9fc;
17'h11bf7:	data_out=16'h8a00;
17'h11bf8:	data_out=16'h99f;
17'h11bf9:	data_out=16'h8a00;
17'h11bfa:	data_out=16'h89e9;
17'h11bfb:	data_out=16'h9f7;
17'h11bfc:	data_out=16'h8a00;
17'h11bfd:	data_out=16'h8178;
17'h11bfe:	data_out=16'h93d;
17'h11bff:	data_out=16'h89fa;
17'h11c00:	data_out=16'h314;
17'h11c01:	data_out=16'ha00;
17'h11c02:	data_out=16'h89e7;
17'h11c03:	data_out=16'h89f3;
17'h11c04:	data_out=16'ha00;
17'h11c05:	data_out=16'h9ef;
17'h11c06:	data_out=16'h990;
17'h11c07:	data_out=16'h8a00;
17'h11c08:	data_out=16'h89be;
17'h11c09:	data_out=16'h89f5;
17'h11c0a:	data_out=16'ha00;
17'h11c0b:	data_out=16'h89a1;
17'h11c0c:	data_out=16'h8a00;
17'h11c0d:	data_out=16'h8a00;
17'h11c0e:	data_out=16'h9fe;
17'h11c0f:	data_out=16'h89ea;
17'h11c10:	data_out=16'h89e5;
17'h11c11:	data_out=16'ha00;
17'h11c12:	data_out=16'h8a00;
17'h11c13:	data_out=16'ha00;
17'h11c14:	data_out=16'h89ea;
17'h11c15:	data_out=16'h346;
17'h11c16:	data_out=16'h8982;
17'h11c17:	data_out=16'h89e9;
17'h11c18:	data_out=16'h8a00;
17'h11c19:	data_out=16'h9ef;
17'h11c1a:	data_out=16'h9f2;
17'h11c1b:	data_out=16'h89e0;
17'h11c1c:	data_out=16'h89f7;
17'h11c1d:	data_out=16'ha00;
17'h11c1e:	data_out=16'h89da;
17'h11c1f:	data_out=16'h8995;
17'h11c20:	data_out=16'ha00;
17'h11c21:	data_out=16'h940;
17'h11c22:	data_out=16'h89ba;
17'h11c23:	data_out=16'ha00;
17'h11c24:	data_out=16'ha00;
17'h11c25:	data_out=16'h8992;
17'h11c26:	data_out=16'h89bf;
17'h11c27:	data_out=16'ha00;
17'h11c28:	data_out=16'h8e1;
17'h11c29:	data_out=16'h8a00;
17'h11c2a:	data_out=16'h8949;
17'h11c2b:	data_out=16'h9f5;
17'h11c2c:	data_out=16'h8971;
17'h11c2d:	data_out=16'hcd;
17'h11c2e:	data_out=16'h8925;
17'h11c2f:	data_out=16'h86b3;
17'h11c30:	data_out=16'h9da;
17'h11c31:	data_out=16'ha00;
17'h11c32:	data_out=16'ha00;
17'h11c33:	data_out=16'h89ec;
17'h11c34:	data_out=16'ha00;
17'h11c35:	data_out=16'ha00;
17'h11c36:	data_out=16'h8960;
17'h11c37:	data_out=16'h89c2;
17'h11c38:	data_out=16'ha00;
17'h11c39:	data_out=16'h89f8;
17'h11c3a:	data_out=16'h89f5;
17'h11c3b:	data_out=16'h9be;
17'h11c3c:	data_out=16'ha00;
17'h11c3d:	data_out=16'h715;
17'h11c3e:	data_out=16'h8e2;
17'h11c3f:	data_out=16'h9ed;
17'h11c40:	data_out=16'ha00;
17'h11c41:	data_out=16'h8a00;
17'h11c42:	data_out=16'h89ff;
17'h11c43:	data_out=16'h89f5;
17'h11c44:	data_out=16'ha00;
17'h11c45:	data_out=16'h29d;
17'h11c46:	data_out=16'h84f5;
17'h11c47:	data_out=16'h89fe;
17'h11c48:	data_out=16'h8852;
17'h11c49:	data_out=16'h8988;
17'h11c4a:	data_out=16'h88ea;
17'h11c4b:	data_out=16'h89fa;
17'h11c4c:	data_out=16'h89fa;
17'h11c4d:	data_out=16'h89ac;
17'h11c4e:	data_out=16'h89f3;
17'h11c4f:	data_out=16'h89ef;
17'h11c50:	data_out=16'h89ad;
17'h11c51:	data_out=16'h89ff;
17'h11c52:	data_out=16'h95f;
17'h11c53:	data_out=16'h9f9;
17'h11c54:	data_out=16'h66a;
17'h11c55:	data_out=16'h89ff;
17'h11c56:	data_out=16'h871c;
17'h11c57:	data_out=16'h8910;
17'h11c58:	data_out=16'h8a00;
17'h11c59:	data_out=16'ha00;
17'h11c5a:	data_out=16'h8a00;
17'h11c5b:	data_out=16'ha00;
17'h11c5c:	data_out=16'h9e9;
17'h11c5d:	data_out=16'h8602;
17'h11c5e:	data_out=16'h853f;
17'h11c5f:	data_out=16'h89bd;
17'h11c60:	data_out=16'h89d8;
17'h11c61:	data_out=16'ha00;
17'h11c62:	data_out=16'h8909;
17'h11c63:	data_out=16'h89dc;
17'h11c64:	data_out=16'ha00;
17'h11c65:	data_out=16'ha00;
17'h11c66:	data_out=16'h6f;
17'h11c67:	data_out=16'h8983;
17'h11c68:	data_out=16'h8fc;
17'h11c69:	data_out=16'h8a00;
17'h11c6a:	data_out=16'h9ff;
17'h11c6b:	data_out=16'h9fe;
17'h11c6c:	data_out=16'h864;
17'h11c6d:	data_out=16'h89de;
17'h11c6e:	data_out=16'h9ff;
17'h11c6f:	data_out=16'ha00;
17'h11c70:	data_out=16'h9fe;
17'h11c71:	data_out=16'h89de;
17'h11c72:	data_out=16'ha00;
17'h11c73:	data_out=16'ha00;
17'h11c74:	data_out=16'h9c1;
17'h11c75:	data_out=16'h9ea;
17'h11c76:	data_out=16'h8096;
17'h11c77:	data_out=16'h89ff;
17'h11c78:	data_out=16'h9aa;
17'h11c79:	data_out=16'h8a00;
17'h11c7a:	data_out=16'h89e1;
17'h11c7b:	data_out=16'h8e0;
17'h11c7c:	data_out=16'h8a00;
17'h11c7d:	data_out=16'h89ec;
17'h11c7e:	data_out=16'h19e;
17'h11c7f:	data_out=16'h89f4;
17'h11c80:	data_out=16'h9f1;
17'h11c81:	data_out=16'ha00;
17'h11c82:	data_out=16'h8a00;
17'h11c83:	data_out=16'h89b2;
17'h11c84:	data_out=16'ha00;
17'h11c85:	data_out=16'h9e9;
17'h11c86:	data_out=16'h9fd;
17'h11c87:	data_out=16'h8a00;
17'h11c88:	data_out=16'h89d7;
17'h11c89:	data_out=16'h8993;
17'h11c8a:	data_out=16'ha00;
17'h11c8b:	data_out=16'h8976;
17'h11c8c:	data_out=16'h8a00;
17'h11c8d:	data_out=16'h8a00;
17'h11c8e:	data_out=16'h89c2;
17'h11c8f:	data_out=16'h89f0;
17'h11c90:	data_out=16'h8757;
17'h11c91:	data_out=16'ha00;
17'h11c92:	data_out=16'h8a00;
17'h11c93:	data_out=16'ha00;
17'h11c94:	data_out=16'h89de;
17'h11c95:	data_out=16'h964;
17'h11c96:	data_out=16'h805b;
17'h11c97:	data_out=16'h89db;
17'h11c98:	data_out=16'h8a00;
17'h11c99:	data_out=16'h9f0;
17'h11c9a:	data_out=16'ha00;
17'h11c9b:	data_out=16'h89d0;
17'h11c9c:	data_out=16'h89e2;
17'h11c9d:	data_out=16'ha00;
17'h11c9e:	data_out=16'h89bb;
17'h11c9f:	data_out=16'h89cd;
17'h11ca0:	data_out=16'h9fe;
17'h11ca1:	data_out=16'h89dd;
17'h11ca2:	data_out=16'h8959;
17'h11ca3:	data_out=16'h9fc;
17'h11ca4:	data_out=16'h9fb;
17'h11ca5:	data_out=16'h88f9;
17'h11ca6:	data_out=16'h89b6;
17'h11ca7:	data_out=16'ha00;
17'h11ca8:	data_out=16'h89e8;
17'h11ca9:	data_out=16'h8a00;
17'h11caa:	data_out=16'h8916;
17'h11cab:	data_out=16'h747;
17'h11cac:	data_out=16'h40c;
17'h11cad:	data_out=16'h598;
17'h11cae:	data_out=16'h88e5;
17'h11caf:	data_out=16'h9c1;
17'h11cb0:	data_out=16'h940;
17'h11cb1:	data_out=16'ha00;
17'h11cb2:	data_out=16'ha00;
17'h11cb3:	data_out=16'h89f3;
17'h11cb4:	data_out=16'ha00;
17'h11cb5:	data_out=16'ha00;
17'h11cb6:	data_out=16'h8951;
17'h11cb7:	data_out=16'h89d0;
17'h11cb8:	data_out=16'ha00;
17'h11cb9:	data_out=16'h89fd;
17'h11cba:	data_out=16'h89b4;
17'h11cbb:	data_out=16'h9b0;
17'h11cbc:	data_out=16'h8298;
17'h11cbd:	data_out=16'h9f9;
17'h11cbe:	data_out=16'h89e8;
17'h11cbf:	data_out=16'h9e7;
17'h11cc0:	data_out=16'ha00;
17'h11cc1:	data_out=16'h8a00;
17'h11cc2:	data_out=16'h8301;
17'h11cc3:	data_out=16'h89fe;
17'h11cc4:	data_out=16'ha00;
17'h11cc5:	data_out=16'h921;
17'h11cc6:	data_out=16'h897d;
17'h11cc7:	data_out=16'h89fc;
17'h11cc8:	data_out=16'h1ae;
17'h11cc9:	data_out=16'h875d;
17'h11cca:	data_out=16'h808a;
17'h11ccb:	data_out=16'h58b;
17'h11ccc:	data_out=16'h89c4;
17'h11ccd:	data_out=16'h8760;
17'h11cce:	data_out=16'h8a00;
17'h11ccf:	data_out=16'h89a4;
17'h11cd0:	data_out=16'h83be;
17'h11cd1:	data_out=16'h8a00;
17'h11cd2:	data_out=16'h9c3;
17'h11cd3:	data_out=16'h81ff;
17'h11cd4:	data_out=16'ha00;
17'h11cd5:	data_out=16'h8a00;
17'h11cd6:	data_out=16'h8972;
17'h11cd7:	data_out=16'h8977;
17'h11cd8:	data_out=16'h8a00;
17'h11cd9:	data_out=16'ha00;
17'h11cda:	data_out=16'h8a00;
17'h11cdb:	data_out=16'ha00;
17'h11cdc:	data_out=16'h7d4;
17'h11cdd:	data_out=16'ha00;
17'h11cde:	data_out=16'ha00;
17'h11cdf:	data_out=16'h892e;
17'h11ce0:	data_out=16'h89a9;
17'h11ce1:	data_out=16'ha00;
17'h11ce2:	data_out=16'h87e3;
17'h11ce3:	data_out=16'h89e2;
17'h11ce4:	data_out=16'ha00;
17'h11ce5:	data_out=16'ha00;
17'h11ce6:	data_out=16'h89e2;
17'h11ce7:	data_out=16'h8996;
17'h11ce8:	data_out=16'h89e8;
17'h11ce9:	data_out=16'h8a00;
17'h11cea:	data_out=16'h89b0;
17'h11ceb:	data_out=16'ha00;
17'h11cec:	data_out=16'ha00;
17'h11ced:	data_out=16'h89e3;
17'h11cee:	data_out=16'h89b1;
17'h11cef:	data_out=16'ha00;
17'h11cf0:	data_out=16'h89bb;
17'h11cf1:	data_out=16'h89fe;
17'h11cf2:	data_out=16'ha00;
17'h11cf3:	data_out=16'ha00;
17'h11cf4:	data_out=16'h91c;
17'h11cf5:	data_out=16'h9f4;
17'h11cf6:	data_out=16'h88b2;
17'h11cf7:	data_out=16'h89c6;
17'h11cf8:	data_out=16'hd2;
17'h11cf9:	data_out=16'h8a00;
17'h11cfa:	data_out=16'h89da;
17'h11cfb:	data_out=16'h89e8;
17'h11cfc:	data_out=16'h8a00;
17'h11cfd:	data_out=16'h89f6;
17'h11cfe:	data_out=16'h8242;
17'h11cff:	data_out=16'h8941;
17'h11d00:	data_out=16'h9eb;
17'h11d01:	data_out=16'ha00;
17'h11d02:	data_out=16'h8a00;
17'h11d03:	data_out=16'h87ad;
17'h11d04:	data_out=16'ha00;
17'h11d05:	data_out=16'h9ea;
17'h11d06:	data_out=16'h9fd;
17'h11d07:	data_out=16'h89fb;
17'h11d08:	data_out=16'h89f1;
17'h11d09:	data_out=16'h853b;
17'h11d0a:	data_out=16'ha00;
17'h11d0b:	data_out=16'h876f;
17'h11d0c:	data_out=16'h76b;
17'h11d0d:	data_out=16'h8a00;
17'h11d0e:	data_out=16'h89fa;
17'h11d0f:	data_out=16'h89ff;
17'h11d10:	data_out=16'ha00;
17'h11d11:	data_out=16'ha00;
17'h11d12:	data_out=16'h8a00;
17'h11d13:	data_out=16'h8ef;
17'h11d14:	data_out=16'h89e8;
17'h11d15:	data_out=16'h9ed;
17'h11d16:	data_out=16'h9ec;
17'h11d17:	data_out=16'h89c3;
17'h11d18:	data_out=16'h8a00;
17'h11d19:	data_out=16'h52e;
17'h11d1a:	data_out=16'ha00;
17'h11d1b:	data_out=16'h89c9;
17'h11d1c:	data_out=16'h89eb;
17'h11d1d:	data_out=16'ha00;
17'h11d1e:	data_out=16'h89d9;
17'h11d1f:	data_out=16'h89f6;
17'h11d20:	data_out=16'ha00;
17'h11d21:	data_out=16'h89fd;
17'h11d22:	data_out=16'h877c;
17'h11d23:	data_out=16'ha00;
17'h11d24:	data_out=16'ha00;
17'h11d25:	data_out=16'h19b;
17'h11d26:	data_out=16'h899b;
17'h11d27:	data_out=16'ha00;
17'h11d28:	data_out=16'h89fe;
17'h11d29:	data_out=16'h8a00;
17'h11d2a:	data_out=16'h874b;
17'h11d2b:	data_out=16'h48e;
17'h11d2c:	data_out=16'h9f0;
17'h11d2d:	data_out=16'h3d3;
17'h11d2e:	data_out=16'h8907;
17'h11d2f:	data_out=16'ha00;
17'h11d30:	data_out=16'h68a;
17'h11d31:	data_out=16'ha00;
17'h11d32:	data_out=16'ha00;
17'h11d33:	data_out=16'h89fc;
17'h11d34:	data_out=16'ha00;
17'h11d35:	data_out=16'ha00;
17'h11d36:	data_out=16'h887e;
17'h11d37:	data_out=16'h89ff;
17'h11d38:	data_out=16'h9fc;
17'h11d39:	data_out=16'h89fb;
17'h11d3a:	data_out=16'h8153;
17'h11d3b:	data_out=16'h9f0;
17'h11d3c:	data_out=16'h8749;
17'h11d3d:	data_out=16'h9f3;
17'h11d3e:	data_out=16'h89fe;
17'h11d3f:	data_out=16'h9e9;
17'h11d40:	data_out=16'ha00;
17'h11d41:	data_out=16'h899b;
17'h11d42:	data_out=16'h9f3;
17'h11d43:	data_out=16'h89ff;
17'h11d44:	data_out=16'ha00;
17'h11d45:	data_out=16'h9ec;
17'h11d46:	data_out=16'h8954;
17'h11d47:	data_out=16'h89f7;
17'h11d48:	data_out=16'ha00;
17'h11d49:	data_out=16'h9f8;
17'h11d4a:	data_out=16'h9fc;
17'h11d4b:	data_out=16'h9f7;
17'h11d4c:	data_out=16'h854a;
17'h11d4d:	data_out=16'h5a2;
17'h11d4e:	data_out=16'h8a00;
17'h11d4f:	data_out=16'h9f7;
17'h11d50:	data_out=16'ha00;
17'h11d51:	data_out=16'h89ff;
17'h11d52:	data_out=16'h9e3;
17'h11d53:	data_out=16'h870e;
17'h11d54:	data_out=16'ha00;
17'h11d55:	data_out=16'h89f7;
17'h11d56:	data_out=16'h89a8;
17'h11d57:	data_out=16'h89ef;
17'h11d58:	data_out=16'h8a00;
17'h11d59:	data_out=16'ha00;
17'h11d5a:	data_out=16'h8a00;
17'h11d5b:	data_out=16'ha00;
17'h11d5c:	data_out=16'h8989;
17'h11d5d:	data_out=16'ha00;
17'h11d5e:	data_out=16'ha00;
17'h11d5f:	data_out=16'h8856;
17'h11d60:	data_out=16'h8945;
17'h11d61:	data_out=16'ha00;
17'h11d62:	data_out=16'h870f;
17'h11d63:	data_out=16'h89fc;
17'h11d64:	data_out=16'ha00;
17'h11d65:	data_out=16'ha00;
17'h11d66:	data_out=16'h89ef;
17'h11d67:	data_out=16'h8a00;
17'h11d68:	data_out=16'h89fe;
17'h11d69:	data_out=16'h8a00;
17'h11d6a:	data_out=16'h89f8;
17'h11d6b:	data_out=16'ha00;
17'h11d6c:	data_out=16'ha00;
17'h11d6d:	data_out=16'h89fc;
17'h11d6e:	data_out=16'h89f8;
17'h11d6f:	data_out=16'ha00;
17'h11d70:	data_out=16'h89f9;
17'h11d71:	data_out=16'h8a00;
17'h11d72:	data_out=16'ha00;
17'h11d73:	data_out=16'ha00;
17'h11d74:	data_out=16'h68b;
17'h11d75:	data_out=16'h8630;
17'h11d76:	data_out=16'h898a;
17'h11d77:	data_out=16'h88ff;
17'h11d78:	data_out=16'h821e;
17'h11d79:	data_out=16'h8a00;
17'h11d7a:	data_out=16'h89f3;
17'h11d7b:	data_out=16'h89fe;
17'h11d7c:	data_out=16'h8a00;
17'h11d7d:	data_out=16'h89f3;
17'h11d7e:	data_out=16'h80e9;
17'h11d7f:	data_out=16'h825b;
17'h11d80:	data_out=16'h9fe;
17'h11d81:	data_out=16'ha00;
17'h11d82:	data_out=16'h8a00;
17'h11d83:	data_out=16'h84cb;
17'h11d84:	data_out=16'ha00;
17'h11d85:	data_out=16'ha00;
17'h11d86:	data_out=16'h9fc;
17'h11d87:	data_out=16'h6cf;
17'h11d88:	data_out=16'h89bb;
17'h11d89:	data_out=16'h959;
17'h11d8a:	data_out=16'ha00;
17'h11d8b:	data_out=16'h8942;
17'h11d8c:	data_out=16'h9fe;
17'h11d8d:	data_out=16'h8a00;
17'h11d8e:	data_out=16'h8a00;
17'h11d8f:	data_out=16'h8a00;
17'h11d90:	data_out=16'ha00;
17'h11d91:	data_out=16'ha00;
17'h11d92:	data_out=16'h8a00;
17'h11d93:	data_out=16'h20c;
17'h11d94:	data_out=16'h89f8;
17'h11d95:	data_out=16'h9fd;
17'h11d96:	data_out=16'ha00;
17'h11d97:	data_out=16'h89e1;
17'h11d98:	data_out=16'h8a00;
17'h11d99:	data_out=16'h89d7;
17'h11d9a:	data_out=16'ha00;
17'h11d9b:	data_out=16'h89ea;
17'h11d9c:	data_out=16'h89ff;
17'h11d9d:	data_out=16'ha00;
17'h11d9e:	data_out=16'h89ef;
17'h11d9f:	data_out=16'h89fa;
17'h11da0:	data_out=16'ha00;
17'h11da1:	data_out=16'h8a00;
17'h11da2:	data_out=16'h88f0;
17'h11da3:	data_out=16'h686;
17'h11da4:	data_out=16'h66b;
17'h11da5:	data_out=16'h84fe;
17'h11da6:	data_out=16'h89b8;
17'h11da7:	data_out=16'ha00;
17'h11da8:	data_out=16'h8a00;
17'h11da9:	data_out=16'h8a00;
17'h11daa:	data_out=16'h8369;
17'h11dab:	data_out=16'h899b;
17'h11dac:	data_out=16'ha00;
17'h11dad:	data_out=16'h89b9;
17'h11dae:	data_out=16'h89a8;
17'h11daf:	data_out=16'ha00;
17'h11db0:	data_out=16'h6e;
17'h11db1:	data_out=16'ha00;
17'h11db2:	data_out=16'ha00;
17'h11db3:	data_out=16'h89ff;
17'h11db4:	data_out=16'ha00;
17'h11db5:	data_out=16'ha00;
17'h11db6:	data_out=16'h87ea;
17'h11db7:	data_out=16'h8a00;
17'h11db8:	data_out=16'h9f8;
17'h11db9:	data_out=16'h8a00;
17'h11dba:	data_out=16'ha00;
17'h11dbb:	data_out=16'h9ff;
17'h11dbc:	data_out=16'h897d;
17'h11dbd:	data_out=16'h9eb;
17'h11dbe:	data_out=16'h8a00;
17'h11dbf:	data_out=16'ha00;
17'h11dc0:	data_out=16'ha00;
17'h11dc1:	data_out=16'h849c;
17'h11dc2:	data_out=16'h9fc;
17'h11dc3:	data_out=16'h8a00;
17'h11dc4:	data_out=16'ha00;
17'h11dc5:	data_out=16'h9fd;
17'h11dc6:	data_out=16'h89a8;
17'h11dc7:	data_out=16'h89e9;
17'h11dc8:	data_out=16'ha00;
17'h11dc9:	data_out=16'h318;
17'h11dca:	data_out=16'ha00;
17'h11dcb:	data_out=16'h9fb;
17'h11dcc:	data_out=16'h85d8;
17'h11dcd:	data_out=16'h998;
17'h11dce:	data_out=16'h886a;
17'h11dcf:	data_out=16'h9f7;
17'h11dd0:	data_out=16'ha00;
17'h11dd1:	data_out=16'h8a00;
17'h11dd2:	data_out=16'h9f8;
17'h11dd3:	data_out=16'h8944;
17'h11dd4:	data_out=16'h9fa;
17'h11dd5:	data_out=16'h89fb;
17'h11dd6:	data_out=16'h89c8;
17'h11dd7:	data_out=16'h89f9;
17'h11dd8:	data_out=16'h8a00;
17'h11dd9:	data_out=16'ha00;
17'h11dda:	data_out=16'h8a00;
17'h11ddb:	data_out=16'h883a;
17'h11ddc:	data_out=16'h89f7;
17'h11ddd:	data_out=16'ha00;
17'h11dde:	data_out=16'ha00;
17'h11ddf:	data_out=16'h48;
17'h11de0:	data_out=16'h8964;
17'h11de1:	data_out=16'ha00;
17'h11de2:	data_out=16'h894a;
17'h11de3:	data_out=16'h8a00;
17'h11de4:	data_out=16'h9f6;
17'h11de5:	data_out=16'ha00;
17'h11de6:	data_out=16'h89f8;
17'h11de7:	data_out=16'h8a00;
17'h11de8:	data_out=16'h8a00;
17'h11de9:	data_out=16'h8a00;
17'h11dea:	data_out=16'h8a00;
17'h11deb:	data_out=16'ha00;
17'h11dec:	data_out=16'ha00;
17'h11ded:	data_out=16'h8a00;
17'h11dee:	data_out=16'h8a00;
17'h11def:	data_out=16'ha00;
17'h11df0:	data_out=16'h8a00;
17'h11df1:	data_out=16'h8a00;
17'h11df2:	data_out=16'ha00;
17'h11df3:	data_out=16'h9fd;
17'h11df4:	data_out=16'h5a;
17'h11df5:	data_out=16'h8955;
17'h11df6:	data_out=16'h89c3;
17'h11df7:	data_out=16'h83be;
17'h11df8:	data_out=16'h8887;
17'h11df9:	data_out=16'h89e1;
17'h11dfa:	data_out=16'h89fc;
17'h11dfb:	data_out=16'h8a00;
17'h11dfc:	data_out=16'h8a00;
17'h11dfd:	data_out=16'h89ee;
17'h11dfe:	data_out=16'h89b7;
17'h11dff:	data_out=16'h9e1;
17'h11e00:	data_out=16'h998;
17'h11e01:	data_out=16'h9e6;
17'h11e02:	data_out=16'h8a00;
17'h11e03:	data_out=16'h87e6;
17'h11e04:	data_out=16'h9fd;
17'h11e05:	data_out=16'h9f9;
17'h11e06:	data_out=16'h78d;
17'h11e07:	data_out=16'h9fc;
17'h11e08:	data_out=16'h89fe;
17'h11e09:	data_out=16'h9f4;
17'h11e0a:	data_out=16'ha00;
17'h11e0b:	data_out=16'h89d9;
17'h11e0c:	data_out=16'h9fe;
17'h11e0d:	data_out=16'h8a00;
17'h11e0e:	data_out=16'h89ff;
17'h11e0f:	data_out=16'h89ff;
17'h11e10:	data_out=16'h9fc;
17'h11e11:	data_out=16'ha00;
17'h11e12:	data_out=16'h8a00;
17'h11e13:	data_out=16'h8a5;
17'h11e14:	data_out=16'h89ff;
17'h11e15:	data_out=16'h9dc;
17'h11e16:	data_out=16'ha00;
17'h11e17:	data_out=16'h89fe;
17'h11e18:	data_out=16'h8a00;
17'h11e19:	data_out=16'h89ac;
17'h11e1a:	data_out=16'h9fa;
17'h11e1b:	data_out=16'h8a00;
17'h11e1c:	data_out=16'h8a00;
17'h11e1d:	data_out=16'ha00;
17'h11e1e:	data_out=16'h89fe;
17'h11e1f:	data_out=16'h8a00;
17'h11e20:	data_out=16'h994;
17'h11e21:	data_out=16'h8a00;
17'h11e22:	data_out=16'h1e2;
17'h11e23:	data_out=16'h8953;
17'h11e24:	data_out=16'h8959;
17'h11e25:	data_out=16'h87c4;
17'h11e26:	data_out=16'h89fd;
17'h11e27:	data_out=16'h9dc;
17'h11e28:	data_out=16'h8a00;
17'h11e29:	data_out=16'h8a00;
17'h11e2a:	data_out=16'h824e;
17'h11e2b:	data_out=16'h89ea;
17'h11e2c:	data_out=16'ha00;
17'h11e2d:	data_out=16'h89fe;
17'h11e2e:	data_out=16'h89fe;
17'h11e2f:	data_out=16'h9fb;
17'h11e30:	data_out=16'h388;
17'h11e31:	data_out=16'h9f4;
17'h11e32:	data_out=16'ha00;
17'h11e33:	data_out=16'h89ff;
17'h11e34:	data_out=16'h9f6;
17'h11e35:	data_out=16'h8fd;
17'h11e36:	data_out=16'h89ba;
17'h11e37:	data_out=16'h8a00;
17'h11e38:	data_out=16'h9dd;
17'h11e39:	data_out=16'h89ff;
17'h11e3a:	data_out=16'h9fd;
17'h11e3b:	data_out=16'h9f8;
17'h11e3c:	data_out=16'h89ff;
17'h11e3d:	data_out=16'h968;
17'h11e3e:	data_out=16'h8a00;
17'h11e3f:	data_out=16'h9f8;
17'h11e40:	data_out=16'ha00;
17'h11e41:	data_out=16'h12;
17'h11e42:	data_out=16'h9fc;
17'h11e43:	data_out=16'h8a00;
17'h11e44:	data_out=16'h280;
17'h11e45:	data_out=16'h9dd;
17'h11e46:	data_out=16'h89f3;
17'h11e47:	data_out=16'h89f9;
17'h11e48:	data_out=16'h9fe;
17'h11e49:	data_out=16'h8191;
17'h11e4a:	data_out=16'h9ff;
17'h11e4b:	data_out=16'h9f9;
17'h11e4c:	data_out=16'h48;
17'h11e4d:	data_out=16'h9f8;
17'h11e4e:	data_out=16'h2f7;
17'h11e4f:	data_out=16'h9f4;
17'h11e50:	data_out=16'h9fe;
17'h11e51:	data_out=16'h8a00;
17'h11e52:	data_out=16'h83d7;
17'h11e53:	data_out=16'h89b4;
17'h11e54:	data_out=16'h9bd;
17'h11e55:	data_out=16'h8a00;
17'h11e56:	data_out=16'h89f8;
17'h11e57:	data_out=16'h89ff;
17'h11e58:	data_out=16'h8a00;
17'h11e59:	data_out=16'ha00;
17'h11e5a:	data_out=16'h8a00;
17'h11e5b:	data_out=16'h89dc;
17'h11e5c:	data_out=16'h89ff;
17'h11e5d:	data_out=16'ha00;
17'h11e5e:	data_out=16'ha00;
17'h11e5f:	data_out=16'h618;
17'h11e60:	data_out=16'h89f9;
17'h11e61:	data_out=16'h9e7;
17'h11e62:	data_out=16'h89fd;
17'h11e63:	data_out=16'h89ff;
17'h11e64:	data_out=16'h9c2;
17'h11e65:	data_out=16'ha00;
17'h11e66:	data_out=16'h8999;
17'h11e67:	data_out=16'h8a00;
17'h11e68:	data_out=16'h8a00;
17'h11e69:	data_out=16'h8a00;
17'h11e6a:	data_out=16'h89ff;
17'h11e6b:	data_out=16'ha00;
17'h11e6c:	data_out=16'h9b4;
17'h11e6d:	data_out=16'h89ff;
17'h11e6e:	data_out=16'h89ff;
17'h11e6f:	data_out=16'ha00;
17'h11e70:	data_out=16'h89ff;
17'h11e71:	data_out=16'h89ff;
17'h11e72:	data_out=16'h9ff;
17'h11e73:	data_out=16'h9dd;
17'h11e74:	data_out=16'h387;
17'h11e75:	data_out=16'h89d4;
17'h11e76:	data_out=16'h89d5;
17'h11e77:	data_out=16'h1f;
17'h11e78:	data_out=16'h8522;
17'h11e79:	data_out=16'h5f9;
17'h11e7a:	data_out=16'h89ff;
17'h11e7b:	data_out=16'h8a00;
17'h11e7c:	data_out=16'h8a00;
17'h11e7d:	data_out=16'h89fb;
17'h11e7e:	data_out=16'h8a00;
17'h11e7f:	data_out=16'h9d3;
17'h11e80:	data_out=16'h7d1;
17'h11e81:	data_out=16'h844;
17'h11e82:	data_out=16'h89ff;
17'h11e83:	data_out=16'h84b8;
17'h11e84:	data_out=16'h9bd;
17'h11e85:	data_out=16'h9c7;
17'h11e86:	data_out=16'h9ec;
17'h11e87:	data_out=16'h9fb;
17'h11e88:	data_out=16'h89fb;
17'h11e89:	data_out=16'h9f6;
17'h11e8a:	data_out=16'h9ea;
17'h11e8b:	data_out=16'h89d8;
17'h11e8c:	data_out=16'h9fc;
17'h11e8d:	data_out=16'h88a1;
17'h11e8e:	data_out=16'h89ff;
17'h11e8f:	data_out=16'h89f2;
17'h11e90:	data_out=16'h9fa;
17'h11e91:	data_out=16'ha00;
17'h11e92:	data_out=16'h8a00;
17'h11e93:	data_out=16'h9c9;
17'h11e94:	data_out=16'h89fe;
17'h11e95:	data_out=16'h986;
17'h11e96:	data_out=16'h9d5;
17'h11e97:	data_out=16'h89fb;
17'h11e98:	data_out=16'h8a00;
17'h11e99:	data_out=16'h8981;
17'h11e9a:	data_out=16'h9c4;
17'h11e9b:	data_out=16'h8a00;
17'h11e9c:	data_out=16'h89ff;
17'h11e9d:	data_out=16'h9da;
17'h11e9e:	data_out=16'h89f8;
17'h11e9f:	data_out=16'h89fe;
17'h11ea0:	data_out=16'h778;
17'h11ea1:	data_out=16'h89ff;
17'h11ea2:	data_out=16'h8632;
17'h11ea3:	data_out=16'h89e5;
17'h11ea4:	data_out=16'h89e6;
17'h11ea5:	data_out=16'h83f5;
17'h11ea6:	data_out=16'h89fe;
17'h11ea7:	data_out=16'h8770;
17'h11ea8:	data_out=16'h89ff;
17'h11ea9:	data_out=16'h89e7;
17'h11eaa:	data_out=16'h811;
17'h11eab:	data_out=16'h89de;
17'h11eac:	data_out=16'h9d5;
17'h11ead:	data_out=16'h8a00;
17'h11eae:	data_out=16'h89fa;
17'h11eaf:	data_out=16'h9ea;
17'h11eb0:	data_out=16'h9fe;
17'h11eb1:	data_out=16'h89c3;
17'h11eb2:	data_out=16'h9f7;
17'h11eb3:	data_out=16'h89ff;
17'h11eb4:	data_out=16'h9c9;
17'h11eb5:	data_out=16'h8037;
17'h11eb6:	data_out=16'h8820;
17'h11eb7:	data_out=16'h89ff;
17'h11eb8:	data_out=16'h9df;
17'h11eb9:	data_out=16'h89ff;
17'h11eba:	data_out=16'h9fb;
17'h11ebb:	data_out=16'h2c2;
17'h11ebc:	data_out=16'h8a00;
17'h11ebd:	data_out=16'h77d;
17'h11ebe:	data_out=16'h89ff;
17'h11ebf:	data_out=16'h9c6;
17'h11ec0:	data_out=16'h9eb;
17'h11ec1:	data_out=16'h9f5;
17'h11ec2:	data_out=16'h9f0;
17'h11ec3:	data_out=16'h89cc;
17'h11ec4:	data_out=16'h89a0;
17'h11ec5:	data_out=16'h9a0;
17'h11ec6:	data_out=16'h89ec;
17'h11ec7:	data_out=16'h89e8;
17'h11ec8:	data_out=16'h9ff;
17'h11ec9:	data_out=16'ha;
17'h11eca:	data_out=16'h9fd;
17'h11ecb:	data_out=16'h9f5;
17'h11ecc:	data_out=16'h85d8;
17'h11ecd:	data_out=16'h83a1;
17'h11ece:	data_out=16'h7ef;
17'h11ecf:	data_out=16'h539;
17'h11ed0:	data_out=16'h9fb;
17'h11ed1:	data_out=16'h8a00;
17'h11ed2:	data_out=16'h89da;
17'h11ed3:	data_out=16'h54f;
17'h11ed4:	data_out=16'h932;
17'h11ed5:	data_out=16'h89fd;
17'h11ed6:	data_out=16'h89fa;
17'h11ed7:	data_out=16'h89ff;
17'h11ed8:	data_out=16'h8a00;
17'h11ed9:	data_out=16'h9d2;
17'h11eda:	data_out=16'h8a00;
17'h11edb:	data_out=16'h8a00;
17'h11edc:	data_out=16'h8a00;
17'h11edd:	data_out=16'ha00;
17'h11ede:	data_out=16'ha00;
17'h11edf:	data_out=16'h11d;
17'h11ee0:	data_out=16'h8a00;
17'h11ee1:	data_out=16'h8425;
17'h11ee2:	data_out=16'h89fc;
17'h11ee3:	data_out=16'h89ff;
17'h11ee4:	data_out=16'h91d;
17'h11ee5:	data_out=16'h9fc;
17'h11ee6:	data_out=16'h9e3;
17'h11ee7:	data_out=16'h8a00;
17'h11ee8:	data_out=16'h89ff;
17'h11ee9:	data_out=16'h8a00;
17'h11eea:	data_out=16'h89ff;
17'h11eeb:	data_out=16'h9e6;
17'h11eec:	data_out=16'h8c6;
17'h11eed:	data_out=16'h89ff;
17'h11eee:	data_out=16'h89ff;
17'h11eef:	data_out=16'h9fd;
17'h11ef0:	data_out=16'h89ff;
17'h11ef1:	data_out=16'h89f5;
17'h11ef2:	data_out=16'h9c0;
17'h11ef3:	data_out=16'h9a6;
17'h11ef4:	data_out=16'h9fd;
17'h11ef5:	data_out=16'h89fc;
17'h11ef6:	data_out=16'h89d5;
17'h11ef7:	data_out=16'h9e7;
17'h11ef8:	data_out=16'h8399;
17'h11ef9:	data_out=16'h9e9;
17'h11efa:	data_out=16'h89fe;
17'h11efb:	data_out=16'h89ff;
17'h11efc:	data_out=16'h8a00;
17'h11efd:	data_out=16'h89e2;
17'h11efe:	data_out=16'h8890;
17'h11eff:	data_out=16'h9a6;
17'h11f00:	data_out=16'h89f8;
17'h11f01:	data_out=16'h8a00;
17'h11f02:	data_out=16'h8a00;
17'h11f03:	data_out=16'h878f;
17'h11f04:	data_out=16'h210;
17'h11f05:	data_out=16'h80d;
17'h11f06:	data_out=16'h9ca;
17'h11f07:	data_out=16'h9fe;
17'h11f08:	data_out=16'h89f9;
17'h11f09:	data_out=16'h9eb;
17'h11f0a:	data_out=16'h8a00;
17'h11f0b:	data_out=16'h89e7;
17'h11f0c:	data_out=16'h9fc;
17'h11f0d:	data_out=16'h6be;
17'h11f0e:	data_out=16'h8a00;
17'h11f0f:	data_out=16'h8010;
17'h11f10:	data_out=16'h9af;
17'h11f11:	data_out=16'h8a00;
17'h11f12:	data_out=16'h89fe;
17'h11f13:	data_out=16'h9fd;
17'h11f14:	data_out=16'h8749;
17'h11f15:	data_out=16'h872a;
17'h11f16:	data_out=16'h9ab;
17'h11f17:	data_out=16'h9ad;
17'h11f18:	data_out=16'h8a00;
17'h11f19:	data_out=16'h8985;
17'h11f1a:	data_out=16'h7bc;
17'h11f1b:	data_out=16'h89ff;
17'h11f1c:	data_out=16'h89fd;
17'h11f1d:	data_out=16'h89fe;
17'h11f1e:	data_out=16'h8212;
17'h11f1f:	data_out=16'h868d;
17'h11f20:	data_out=16'h257;
17'h11f21:	data_out=16'h8a00;
17'h11f22:	data_out=16'h89d9;
17'h11f23:	data_out=16'h89f6;
17'h11f24:	data_out=16'h89f7;
17'h11f25:	data_out=16'h84a9;
17'h11f26:	data_out=16'h8a00;
17'h11f27:	data_out=16'h8a00;
17'h11f28:	data_out=16'h88d3;
17'h11f29:	data_out=16'h89f3;
17'h11f2a:	data_out=16'h6ac;
17'h11f2b:	data_out=16'h89c0;
17'h11f2c:	data_out=16'h9ae;
17'h11f2d:	data_out=16'h8a00;
17'h11f2e:	data_out=16'h89f7;
17'h11f2f:	data_out=16'h9ad;
17'h11f30:	data_out=16'ha00;
17'h11f31:	data_out=16'h8a00;
17'h11f32:	data_out=16'h8c1;
17'h11f33:	data_out=16'h887f;
17'h11f34:	data_out=16'h8056;
17'h11f35:	data_out=16'h89f2;
17'h11f36:	data_out=16'h8785;
17'h11f37:	data_out=16'h8a00;
17'h11f38:	data_out=16'h984;
17'h11f39:	data_out=16'h89f3;
17'h11f3a:	data_out=16'h9f9;
17'h11f3b:	data_out=16'h8a00;
17'h11f3c:	data_out=16'h8a00;
17'h11f3d:	data_out=16'h89fc;
17'h11f3e:	data_out=16'h88b0;
17'h11f3f:	data_out=16'h7f8;
17'h11f40:	data_out=16'h968;
17'h11f41:	data_out=16'h70f;
17'h11f42:	data_out=16'h923;
17'h11f43:	data_out=16'hf4;
17'h11f44:	data_out=16'h8a00;
17'h11f45:	data_out=16'h84e7;
17'h11f46:	data_out=16'h8a00;
17'h11f47:	data_out=16'h8904;
17'h11f48:	data_out=16'h9f6;
17'h11f49:	data_out=16'h82c7;
17'h11f4a:	data_out=16'h9f7;
17'h11f4b:	data_out=16'h9c9;
17'h11f4c:	data_out=16'h89f9;
17'h11f4d:	data_out=16'h8950;
17'h11f4e:	data_out=16'h676;
17'h11f4f:	data_out=16'h813b;
17'h11f50:	data_out=16'h9d4;
17'h11f51:	data_out=16'h89fb;
17'h11f52:	data_out=16'h89f1;
17'h11f53:	data_out=16'h651;
17'h11f54:	data_out=16'h63c;
17'h11f55:	data_out=16'h897f;
17'h11f56:	data_out=16'h8a00;
17'h11f57:	data_out=16'h8a00;
17'h11f58:	data_out=16'h89fe;
17'h11f59:	data_out=16'h89da;
17'h11f5a:	data_out=16'h89f9;
17'h11f5b:	data_out=16'h8a00;
17'h11f5c:	data_out=16'h848b;
17'h11f5d:	data_out=16'h9aa;
17'h11f5e:	data_out=16'ha00;
17'h11f5f:	data_out=16'h874d;
17'h11f60:	data_out=16'h8a00;
17'h11f61:	data_out=16'h8a00;
17'h11f62:	data_out=16'h344;
17'h11f63:	data_out=16'h8715;
17'h11f64:	data_out=16'h39b;
17'h11f65:	data_out=16'h9a4;
17'h11f66:	data_out=16'h9f1;
17'h11f67:	data_out=16'h8a00;
17'h11f68:	data_out=16'h8a00;
17'h11f69:	data_out=16'h89fd;
17'h11f6a:	data_out=16'h8a00;
17'h11f6b:	data_out=16'h9c0;
17'h11f6c:	data_out=16'h89fc;
17'h11f6d:	data_out=16'h876f;
17'h11f6e:	data_out=16'h8a00;
17'h11f6f:	data_out=16'h9d6;
17'h11f70:	data_out=16'h8a00;
17'h11f71:	data_out=16'h840b;
17'h11f72:	data_out=16'h43a;
17'h11f73:	data_out=16'h56d;
17'h11f74:	data_out=16'ha00;
17'h11f75:	data_out=16'h89ff;
17'h11f76:	data_out=16'h8a00;
17'h11f77:	data_out=16'h9d3;
17'h11f78:	data_out=16'h9ec;
17'h11f79:	data_out=16'h398;
17'h11f7a:	data_out=16'h8684;
17'h11f7b:	data_out=16'h889f;
17'h11f7c:	data_out=16'h89ff;
17'h11f7d:	data_out=16'h98d;
17'h11f7e:	data_out=16'h922;
17'h11f7f:	data_out=16'h89fc;
17'h11f80:	data_out=16'h89d8;
17'h11f81:	data_out=16'h863e;
17'h11f82:	data_out=16'h89ff;
17'h11f83:	data_out=16'h884f;
17'h11f84:	data_out=16'h4b5;
17'h11f85:	data_out=16'h8bc;
17'h11f86:	data_out=16'h7c4;
17'h11f87:	data_out=16'h9ff;
17'h11f88:	data_out=16'h89d0;
17'h11f89:	data_out=16'h9cc;
17'h11f8a:	data_out=16'h8a00;
17'h11f8b:	data_out=16'h89d7;
17'h11f8c:	data_out=16'h9fd;
17'h11f8d:	data_out=16'h25e;
17'h11f8e:	data_out=16'h747;
17'h11f8f:	data_out=16'h60c;
17'h11f90:	data_out=16'h16e;
17'h11f91:	data_out=16'h8a00;
17'h11f92:	data_out=16'h89c4;
17'h11f93:	data_out=16'h9ef;
17'h11f94:	data_out=16'h8704;
17'h11f95:	data_out=16'h1c3;
17'h11f96:	data_out=16'h9de;
17'h11f97:	data_out=16'h98b;
17'h11f98:	data_out=16'h89ef;
17'h11f99:	data_out=16'h9aa;
17'h11f9a:	data_out=16'h78d;
17'h11f9b:	data_out=16'h80d6;
17'h11f9c:	data_out=16'h8a00;
17'h11f9d:	data_out=16'h546;
17'h11f9e:	data_out=16'h1a4;
17'h11f9f:	data_out=16'h83c6;
17'h11fa0:	data_out=16'h42e;
17'h11fa1:	data_out=16'h7fa;
17'h11fa2:	data_out=16'h8a00;
17'h11fa3:	data_out=16'h89e9;
17'h11fa4:	data_out=16'h89eb;
17'h11fa5:	data_out=16'h80e7;
17'h11fa6:	data_out=16'h89fd;
17'h11fa7:	data_out=16'h376;
17'h11fa8:	data_out=16'h8b1;
17'h11fa9:	data_out=16'h89fe;
17'h11faa:	data_out=16'h7ee;
17'h11fab:	data_out=16'h89b1;
17'h11fac:	data_out=16'h9e8;
17'h11fad:	data_out=16'h89fb;
17'h11fae:	data_out=16'h89be;
17'h11faf:	data_out=16'h97b;
17'h11fb0:	data_out=16'ha00;
17'h11fb1:	data_out=16'h327;
17'h11fb2:	data_out=16'h60c;
17'h11fb3:	data_out=16'h8993;
17'h11fb4:	data_out=16'hf7;
17'h11fb5:	data_out=16'h1f3;
17'h11fb6:	data_out=16'h842f;
17'h11fb7:	data_out=16'h8a00;
17'h11fb8:	data_out=16'h8a00;
17'h11fb9:	data_out=16'h89e5;
17'h11fba:	data_out=16'h9fd;
17'h11fbb:	data_out=16'h50e;
17'h11fbc:	data_out=16'h8a00;
17'h11fbd:	data_out=16'h89fb;
17'h11fbe:	data_out=16'h8b5;
17'h11fbf:	data_out=16'h894;
17'h11fc0:	data_out=16'h94e;
17'h11fc1:	data_out=16'h541;
17'h11fc2:	data_out=16'h2da;
17'h11fc3:	data_out=16'h9ff;
17'h11fc4:	data_out=16'h2b3;
17'h11fc5:	data_out=16'h58f;
17'h11fc6:	data_out=16'h8a00;
17'h11fc7:	data_out=16'h824d;
17'h11fc8:	data_out=16'h9d7;
17'h11fc9:	data_out=16'h52f;
17'h11fca:	data_out=16'h9f9;
17'h11fcb:	data_out=16'h975;
17'h11fcc:	data_out=16'h8a00;
17'h11fcd:	data_out=16'h8a00;
17'h11fce:	data_out=16'h473;
17'h11fcf:	data_out=16'h8f4;
17'h11fd0:	data_out=16'h5dc;
17'h11fd1:	data_out=16'h89e9;
17'h11fd2:	data_out=16'h89b6;
17'h11fd3:	data_out=16'h5f5;
17'h11fd4:	data_out=16'h234;
17'h11fd5:	data_out=16'h84de;
17'h11fd6:	data_out=16'h89ff;
17'h11fd7:	data_out=16'h8a00;
17'h11fd8:	data_out=16'h89ff;
17'h11fd9:	data_out=16'h3cc;
17'h11fda:	data_out=16'h853e;
17'h11fdb:	data_out=16'h8a00;
17'h11fdc:	data_out=16'h8027;
17'h11fdd:	data_out=16'h9ab;
17'h11fde:	data_out=16'ha00;
17'h11fdf:	data_out=16'h89ec;
17'h11fe0:	data_out=16'h8a00;
17'h11fe1:	data_out=16'h158;
17'h11fe2:	data_out=16'h9a2;
17'h11fe3:	data_out=16'h896a;
17'h11fe4:	data_out=16'h821e;
17'h11fe5:	data_out=16'h88b;
17'h11fe6:	data_out=16'ha00;
17'h11fe7:	data_out=16'h89fc;
17'h11fe8:	data_out=16'h857;
17'h11fe9:	data_out=16'h89f3;
17'h11fea:	data_out=16'h6bc;
17'h11feb:	data_out=16'h9ce;
17'h11fec:	data_out=16'h89f8;
17'h11fed:	data_out=16'h897d;
17'h11fee:	data_out=16'h6c1;
17'h11fef:	data_out=16'h9d3;
17'h11ff0:	data_out=16'h712;
17'h11ff1:	data_out=16'h761;
17'h11ff2:	data_out=16'h95a;
17'h11ff3:	data_out=16'h782;
17'h11ff4:	data_out=16'ha00;
17'h11ff5:	data_out=16'h8618;
17'h11ff6:	data_out=16'h89fe;
17'h11ff7:	data_out=16'h950;
17'h11ff8:	data_out=16'h97a;
17'h11ff9:	data_out=16'h82a9;
17'h11ffa:	data_out=16'h857a;
17'h11ffb:	data_out=16'h8b8;
17'h11ffc:	data_out=16'h89ed;
17'h11ffd:	data_out=16'h9f8;
17'h11ffe:	data_out=16'h9b4;
17'h11fff:	data_out=16'h8a00;
17'h12000:	data_out=16'h88fc;
17'h12001:	data_out=16'h897a;
17'h12002:	data_out=16'h873d;
17'h12003:	data_out=16'h9cb;
17'h12004:	data_out=16'h9db;
17'h12005:	data_out=16'h9e5;
17'h12006:	data_out=16'h8a00;
17'h12007:	data_out=16'h9fb;
17'h12008:	data_out=16'h89ae;
17'h12009:	data_out=16'h8138;
17'h1200a:	data_out=16'h887b;
17'h1200b:	data_out=16'h89e2;
17'h1200c:	data_out=16'h98d;
17'h1200d:	data_out=16'h963;
17'h1200e:	data_out=16'h908;
17'h1200f:	data_out=16'h56c;
17'h12010:	data_out=16'h83d1;
17'h12011:	data_out=16'h8a00;
17'h12012:	data_out=16'h89e5;
17'h12013:	data_out=16'h9ce;
17'h12014:	data_out=16'h9b5;
17'h12015:	data_out=16'h9f4;
17'h12016:	data_out=16'h9f7;
17'h12017:	data_out=16'h9c0;
17'h12018:	data_out=16'h89f5;
17'h12019:	data_out=16'h9f0;
17'h1201a:	data_out=16'h9e0;
17'h1201b:	data_out=16'h862;
17'h1201c:	data_out=16'h89eb;
17'h1201d:	data_out=16'h8537;
17'h1201e:	data_out=16'h9b8;
17'h1201f:	data_out=16'h998;
17'h12020:	data_out=16'h90b;
17'h12021:	data_out=16'h946;
17'h12022:	data_out=16'h8a00;
17'h12023:	data_out=16'h89dd;
17'h12024:	data_out=16'h89dd;
17'h12025:	data_out=16'h89eb;
17'h12026:	data_out=16'h89fe;
17'h12027:	data_out=16'h705;
17'h12028:	data_out=16'h973;
17'h12029:	data_out=16'h84b;
17'h1202a:	data_out=16'h84d0;
17'h1202b:	data_out=16'h887a;
17'h1202c:	data_out=16'h9fa;
17'h1202d:	data_out=16'h89fe;
17'h1202e:	data_out=16'h89ee;
17'h1202f:	data_out=16'h9e5;
17'h12030:	data_out=16'ha00;
17'h12031:	data_out=16'h9d7;
17'h12032:	data_out=16'h768;
17'h12033:	data_out=16'h84b7;
17'h12034:	data_out=16'h8880;
17'h12035:	data_out=16'h649;
17'h12036:	data_out=16'h8094;
17'h12037:	data_out=16'h88b2;
17'h12038:	data_out=16'h8a00;
17'h12039:	data_out=16'h89ef;
17'h1203a:	data_out=16'h99b;
17'h1203b:	data_out=16'h9f8;
17'h1203c:	data_out=16'h8a00;
17'h1203d:	data_out=16'h326;
17'h1203e:	data_out=16'h974;
17'h1203f:	data_out=16'h9e5;
17'h12040:	data_out=16'h9d3;
17'h12041:	data_out=16'h872;
17'h12042:	data_out=16'h89ee;
17'h12043:	data_out=16'ha00;
17'h12044:	data_out=16'h9c5;
17'h12045:	data_out=16'h9f3;
17'h12046:	data_out=16'h8a00;
17'h12047:	data_out=16'h89d6;
17'h12048:	data_out=16'h8918;
17'h12049:	data_out=16'h76a;
17'h1204a:	data_out=16'ha00;
17'h1204b:	data_out=16'h89c4;
17'h1204c:	data_out=16'h8a00;
17'h1204d:	data_out=16'h8a00;
17'h1204e:	data_out=16'h4a5;
17'h1204f:	data_out=16'h8744;
17'h12050:	data_out=16'h9f7;
17'h12051:	data_out=16'h8ac;
17'h12052:	data_out=16'h858e;
17'h12053:	data_out=16'h93c;
17'h12054:	data_out=16'h8976;
17'h12055:	data_out=16'h9c9;
17'h12056:	data_out=16'h89fb;
17'h12057:	data_out=16'h89ff;
17'h12058:	data_out=16'h403;
17'h12059:	data_out=16'h367;
17'h1205a:	data_out=16'h8139;
17'h1205b:	data_out=16'h4d8;
17'h1205c:	data_out=16'h88a;
17'h1205d:	data_out=16'h9f2;
17'h1205e:	data_out=16'ha00;
17'h1205f:	data_out=16'h89e6;
17'h12060:	data_out=16'h8a00;
17'h12061:	data_out=16'h663;
17'h12062:	data_out=16'h9c6;
17'h12063:	data_out=16'h5;
17'h12064:	data_out=16'h89e1;
17'h12065:	data_out=16'h832;
17'h12066:	data_out=16'ha00;
17'h12067:	data_out=16'h8ea;
17'h12068:	data_out=16'h962;
17'h12069:	data_out=16'h89fe;
17'h1206a:	data_out=16'h8cb;
17'h1206b:	data_out=16'h9ea;
17'h1206c:	data_out=16'h875f;
17'h1206d:	data_out=16'h8134;
17'h1206e:	data_out=16'h8ce;
17'h1206f:	data_out=16'h9f8;
17'h12070:	data_out=16'h8f6;
17'h12071:	data_out=16'h8ec;
17'h12072:	data_out=16'h8fa;
17'h12073:	data_out=16'h8fa;
17'h12074:	data_out=16'ha00;
17'h12075:	data_out=16'h70a;
17'h12076:	data_out=16'h89f9;
17'h12077:	data_out=16'h6fc;
17'h12078:	data_out=16'h44d;
17'h12079:	data_out=16'h3ea;
17'h1207a:	data_out=16'h9aa;
17'h1207b:	data_out=16'h975;
17'h1207c:	data_out=16'h89f0;
17'h1207d:	data_out=16'h9fd;
17'h1207e:	data_out=16'h2e0;
17'h1207f:	data_out=16'h8486;
17'h12080:	data_out=16'h88cb;
17'h12081:	data_out=16'h85ea;
17'h12082:	data_out=16'h86fa;
17'h12083:	data_out=16'h7e4;
17'h12084:	data_out=16'h9f6;
17'h12085:	data_out=16'ha00;
17'h12086:	data_out=16'h8a00;
17'h12087:	data_out=16'h9f6;
17'h12088:	data_out=16'h89d0;
17'h12089:	data_out=16'h89d8;
17'h1208a:	data_out=16'h8f7;
17'h1208b:	data_out=16'h89f0;
17'h1208c:	data_out=16'h8d8;
17'h1208d:	data_out=16'h7e0;
17'h1208e:	data_out=16'h9b6;
17'h1208f:	data_out=16'h8175;
17'h12090:	data_out=16'h89d0;
17'h12091:	data_out=16'h89fd;
17'h12092:	data_out=16'h89ff;
17'h12093:	data_out=16'h935;
17'h12094:	data_out=16'h22c;
17'h12095:	data_out=16'h9f5;
17'h12096:	data_out=16'h9f8;
17'h12097:	data_out=16'h9cb;
17'h12098:	data_out=16'h89fe;
17'h12099:	data_out=16'ha00;
17'h1209a:	data_out=16'ha00;
17'h1209b:	data_out=16'h70f;
17'h1209c:	data_out=16'h896d;
17'h1209d:	data_out=16'h877c;
17'h1209e:	data_out=16'hf2;
17'h1209f:	data_out=16'h3d9;
17'h120a0:	data_out=16'h8710;
17'h120a1:	data_out=16'h9c9;
17'h120a2:	data_out=16'h8a00;
17'h120a3:	data_out=16'h253;
17'h120a4:	data_out=16'h270;
17'h120a5:	data_out=16'h87ec;
17'h120a6:	data_out=16'h8a00;
17'h120a7:	data_out=16'h9c8;
17'h120a8:	data_out=16'h9dd;
17'h120a9:	data_out=16'h9e8;
17'h120aa:	data_out=16'h84a8;
17'h120ab:	data_out=16'h8782;
17'h120ac:	data_out=16'h9fa;
17'h120ad:	data_out=16'h89fe;
17'h120ae:	data_out=16'h89f8;
17'h120af:	data_out=16'h9f2;
17'h120b0:	data_out=16'ha00;
17'h120b1:	data_out=16'h9f8;
17'h120b2:	data_out=16'ha00;
17'h120b3:	data_out=16'h89f4;
17'h120b4:	data_out=16'h87ea;
17'h120b5:	data_out=16'h9bf;
17'h120b6:	data_out=16'h88f9;
17'h120b7:	data_out=16'h8288;
17'h120b8:	data_out=16'h8a00;
17'h120b9:	data_out=16'h89f7;
17'h120ba:	data_out=16'h8475;
17'h120bb:	data_out=16'ha00;
17'h120bc:	data_out=16'h20;
17'h120bd:	data_out=16'h81f5;
17'h120be:	data_out=16'h9de;
17'h120bf:	data_out=16'ha00;
17'h120c0:	data_out=16'h9f8;
17'h120c1:	data_out=16'h830;
17'h120c2:	data_out=16'h89db;
17'h120c3:	data_out=16'h9fa;
17'h120c4:	data_out=16'h9d2;
17'h120c5:	data_out=16'h9f5;
17'h120c6:	data_out=16'h89fe;
17'h120c7:	data_out=16'h8a00;
17'h120c8:	data_out=16'h89dc;
17'h120c9:	data_out=16'h81bc;
17'h120ca:	data_out=16'ha00;
17'h120cb:	data_out=16'h89e5;
17'h120cc:	data_out=16'h8a00;
17'h120cd:	data_out=16'h8a00;
17'h120ce:	data_out=16'h3e6;
17'h120cf:	data_out=16'h89f8;
17'h120d0:	data_out=16'h9f9;
17'h120d1:	data_out=16'h84b;
17'h120d2:	data_out=16'h816;
17'h120d3:	data_out=16'h9ed;
17'h120d4:	data_out=16'h88f6;
17'h120d5:	data_out=16'h9c8;
17'h120d6:	data_out=16'h86c5;
17'h120d7:	data_out=16'h8a00;
17'h120d8:	data_out=16'h642;
17'h120d9:	data_out=16'h95f;
17'h120da:	data_out=16'h8947;
17'h120db:	data_out=16'h9b2;
17'h120dc:	data_out=16'h9db;
17'h120dd:	data_out=16'ha00;
17'h120de:	data_out=16'ha00;
17'h120df:	data_out=16'h89f4;
17'h120e0:	data_out=16'h89f0;
17'h120e1:	data_out=16'h9ec;
17'h120e2:	data_out=16'h421;
17'h120e3:	data_out=16'h877f;
17'h120e4:	data_out=16'h89f3;
17'h120e5:	data_out=16'ha00;
17'h120e6:	data_out=16'ha00;
17'h120e7:	data_out=16'h9ff;
17'h120e8:	data_out=16'h9d2;
17'h120e9:	data_out=16'h89ff;
17'h120ea:	data_out=16'h9a0;
17'h120eb:	data_out=16'h9f4;
17'h120ec:	data_out=16'h83ea;
17'h120ed:	data_out=16'h8858;
17'h120ee:	data_out=16'h9a1;
17'h120ef:	data_out=16'ha00;
17'h120f0:	data_out=16'h9ae;
17'h120f1:	data_out=16'h989;
17'h120f2:	data_out=16'h482;
17'h120f3:	data_out=16'h9de;
17'h120f4:	data_out=16'ha00;
17'h120f5:	data_out=16'h9e5;
17'h120f6:	data_out=16'h8851;
17'h120f7:	data_out=16'h86e7;
17'h120f8:	data_out=16'h80a0;
17'h120f9:	data_out=16'h45f;
17'h120fa:	data_out=16'h3;
17'h120fb:	data_out=16'h9de;
17'h120fc:	data_out=16'h89fd;
17'h120fd:	data_out=16'h9f4;
17'h120fe:	data_out=16'h89fc;
17'h120ff:	data_out=16'h8823;
17'h12100:	data_out=16'h89a0;
17'h12101:	data_out=16'h89dc;
17'h12102:	data_out=16'h89f9;
17'h12103:	data_out=16'h2aa;
17'h12104:	data_out=16'ha00;
17'h12105:	data_out=16'ha00;
17'h12106:	data_out=16'h89dd;
17'h12107:	data_out=16'h9e6;
17'h12108:	data_out=16'h89de;
17'h12109:	data_out=16'h89a8;
17'h1210a:	data_out=16'h8be;
17'h1210b:	data_out=16'h89e6;
17'h1210c:	data_out=16'h3bc;
17'h1210d:	data_out=16'h85dd;
17'h1210e:	data_out=16'h9f8;
17'h1210f:	data_out=16'h89b6;
17'h12110:	data_out=16'h8829;
17'h12111:	data_out=16'h89ff;
17'h12112:	data_out=16'h89fe;
17'h12113:	data_out=16'h846d;
17'h12114:	data_out=16'h820f;
17'h12115:	data_out=16'h9fe;
17'h12116:	data_out=16'ha00;
17'h12117:	data_out=16'h177;
17'h12118:	data_out=16'h89f9;
17'h12119:	data_out=16'ha00;
17'h1211a:	data_out=16'ha00;
17'h1211b:	data_out=16'h857d;
17'h1211c:	data_out=16'h85de;
17'h1211d:	data_out=16'h89ff;
17'h1211e:	data_out=16'h82e4;
17'h1211f:	data_out=16'h21a;
17'h12120:	data_out=16'h8277;
17'h12121:	data_out=16'h9f9;
17'h12122:	data_out=16'h89eb;
17'h12123:	data_out=16'h698;
17'h12124:	data_out=16'h69e;
17'h12125:	data_out=16'h8333;
17'h12126:	data_out=16'h8a00;
17'h12127:	data_out=16'h81a0;
17'h12128:	data_out=16'h9fa;
17'h12129:	data_out=16'h9f2;
17'h1212a:	data_out=16'h893f;
17'h1212b:	data_out=16'h489;
17'h1212c:	data_out=16'h9ff;
17'h1212d:	data_out=16'h8a00;
17'h1212e:	data_out=16'h89e7;
17'h1212f:	data_out=16'h2ec;
17'h12130:	data_out=16'ha00;
17'h12131:	data_out=16'h9f1;
17'h12132:	data_out=16'ha00;
17'h12133:	data_out=16'h89cd;
17'h12134:	data_out=16'h89e9;
17'h12135:	data_out=16'h9b0;
17'h12136:	data_out=16'h895f;
17'h12137:	data_out=16'h89f8;
17'h12138:	data_out=16'h8a00;
17'h12139:	data_out=16'h89df;
17'h1213a:	data_out=16'h8555;
17'h1213b:	data_out=16'ha00;
17'h1213c:	data_out=16'hfc;
17'h1213d:	data_out=16'h3aa;
17'h1213e:	data_out=16'h9fa;
17'h1213f:	data_out=16'ha00;
17'h12140:	data_out=16'ha00;
17'h12141:	data_out=16'h1af;
17'h12142:	data_out=16'h8a00;
17'h12143:	data_out=16'h9f0;
17'h12144:	data_out=16'h9f9;
17'h12145:	data_out=16'h9fe;
17'h12146:	data_out=16'h8a00;
17'h12147:	data_out=16'h8a00;
17'h12148:	data_out=16'h89d8;
17'h12149:	data_out=16'h398;
17'h1214a:	data_out=16'ha00;
17'h1214b:	data_out=16'h89f7;
17'h1214c:	data_out=16'h89ff;
17'h1214d:	data_out=16'h89a9;
17'h1214e:	data_out=16'h8379;
17'h1214f:	data_out=16'h89f0;
17'h12150:	data_out=16'ha00;
17'h12151:	data_out=16'h933;
17'h12152:	data_out=16'h70d;
17'h12153:	data_out=16'h84ac;
17'h12154:	data_out=16'h883b;
17'h12155:	data_out=16'h9e8;
17'h12156:	data_out=16'h8432;
17'h12157:	data_out=16'h86a2;
17'h12158:	data_out=16'h82d;
17'h12159:	data_out=16'h4f2;
17'h1215a:	data_out=16'h89d8;
17'h1215b:	data_out=16'h9ea;
17'h1215c:	data_out=16'h9eb;
17'h1215d:	data_out=16'h926;
17'h1215e:	data_out=16'h7aa;
17'h1215f:	data_out=16'h89e6;
17'h12160:	data_out=16'h8a00;
17'h12161:	data_out=16'ha00;
17'h12162:	data_out=16'h84ef;
17'h12163:	data_out=16'h891d;
17'h12164:	data_out=16'h8a00;
17'h12165:	data_out=16'ha00;
17'h12166:	data_out=16'ha00;
17'h12167:	data_out=16'ha00;
17'h12168:	data_out=16'h9f9;
17'h12169:	data_out=16'h8a00;
17'h1216a:	data_out=16'h9f4;
17'h1216b:	data_out=16'ha00;
17'h1216c:	data_out=16'h84b2;
17'h1216d:	data_out=16'h8955;
17'h1216e:	data_out=16'h9f5;
17'h1216f:	data_out=16'ha00;
17'h12170:	data_out=16'h9f7;
17'h12171:	data_out=16'h8502;
17'h12172:	data_out=16'h8230;
17'h12173:	data_out=16'h9f5;
17'h12174:	data_out=16'ha00;
17'h12175:	data_out=16'h9f0;
17'h12176:	data_out=16'ha00;
17'h12177:	data_out=16'h85ea;
17'h12178:	data_out=16'h8e;
17'h12179:	data_out=16'hcd;
17'h1217a:	data_out=16'h8437;
17'h1217b:	data_out=16'h9fa;
17'h1217c:	data_out=16'h89ee;
17'h1217d:	data_out=16'ha00;
17'h1217e:	data_out=16'h89e7;
17'h1217f:	data_out=16'h732;
17'h12180:	data_out=16'h891b;
17'h12181:	data_out=16'h89dc;
17'h12182:	data_out=16'h89f0;
17'h12183:	data_out=16'h8614;
17'h12184:	data_out=16'ha00;
17'h12185:	data_out=16'ha00;
17'h12186:	data_out=16'h89d1;
17'h12187:	data_out=16'h821b;
17'h12188:	data_out=16'h89f6;
17'h12189:	data_out=16'h89c1;
17'h1218a:	data_out=16'h99f;
17'h1218b:	data_out=16'h89da;
17'h1218c:	data_out=16'h80aa;
17'h1218d:	data_out=16'h89d6;
17'h1218e:	data_out=16'h9fc;
17'h1218f:	data_out=16'h89e8;
17'h12190:	data_out=16'h85e0;
17'h12191:	data_out=16'h89e9;
17'h12192:	data_out=16'h89fc;
17'h12193:	data_out=16'h89b9;
17'h12194:	data_out=16'h879a;
17'h12195:	data_out=16'ha00;
17'h12196:	data_out=16'ha00;
17'h12197:	data_out=16'h87ac;
17'h12198:	data_out=16'h89f6;
17'h12199:	data_out=16'ha00;
17'h1219a:	data_out=16'ha00;
17'h1219b:	data_out=16'h8890;
17'h1219c:	data_out=16'h8785;
17'h1219d:	data_out=16'h89f4;
17'h1219e:	data_out=16'h8828;
17'h1219f:	data_out=16'h8591;
17'h121a0:	data_out=16'h846a;
17'h121a1:	data_out=16'h9fd;
17'h121a2:	data_out=16'h8812;
17'h121a3:	data_out=16'h91f;
17'h121a4:	data_out=16'h92b;
17'h121a5:	data_out=16'h8521;
17'h121a6:	data_out=16'h8a00;
17'h121a7:	data_out=16'h8749;
17'h121a8:	data_out=16'h9fd;
17'h121a9:	data_out=16'h9f9;
17'h121aa:	data_out=16'h89cf;
17'h121ab:	data_out=16'ha00;
17'h121ac:	data_out=16'ha00;
17'h121ad:	data_out=16'h8a00;
17'h121ae:	data_out=16'h89c8;
17'h121af:	data_out=16'h84c3;
17'h121b0:	data_out=16'ha00;
17'h121b1:	data_out=16'h9fc;
17'h121b2:	data_out=16'h9f1;
17'h121b3:	data_out=16'h8975;
17'h121b4:	data_out=16'h89f8;
17'h121b5:	data_out=16'h9e8;
17'h121b6:	data_out=16'h89b6;
17'h121b7:	data_out=16'h89ed;
17'h121b8:	data_out=16'h8a00;
17'h121b9:	data_out=16'h89ba;
17'h121ba:	data_out=16'h8796;
17'h121bb:	data_out=16'ha00;
17'h121bc:	data_out=16'h6b3;
17'h121bd:	data_out=16'h8063;
17'h121be:	data_out=16'h9fd;
17'h121bf:	data_out=16'ha00;
17'h121c0:	data_out=16'ha00;
17'h121c1:	data_out=16'h86c9;
17'h121c2:	data_out=16'h8a00;
17'h121c3:	data_out=16'ha00;
17'h121c4:	data_out=16'h9ff;
17'h121c5:	data_out=16'ha00;
17'h121c6:	data_out=16'h8a00;
17'h121c7:	data_out=16'h8a00;
17'h121c8:	data_out=16'h89de;
17'h121c9:	data_out=16'hcc;
17'h121ca:	data_out=16'h863b;
17'h121cb:	data_out=16'h8a00;
17'h121cc:	data_out=16'h89ff;
17'h121cd:	data_out=16'h873c;
17'h121ce:	data_out=16'h8a00;
17'h121cf:	data_out=16'h89fe;
17'h121d0:	data_out=16'ha00;
17'h121d1:	data_out=16'h91f;
17'h121d2:	data_out=16'h9ea;
17'h121d3:	data_out=16'h86b9;
17'h121d4:	data_out=16'h888a;
17'h121d5:	data_out=16'h4d;
17'h121d6:	data_out=16'h446;
17'h121d7:	data_out=16'h84cd;
17'h121d8:	data_out=16'h1e5;
17'h121d9:	data_out=16'h812b;
17'h121da:	data_out=16'h89c8;
17'h121db:	data_out=16'ha00;
17'h121dc:	data_out=16'h816b;
17'h121dd:	data_out=16'h80eb;
17'h121de:	data_out=16'h8342;
17'h121df:	data_out=16'h89f6;
17'h121e0:	data_out=16'h8a00;
17'h121e1:	data_out=16'ha00;
17'h121e2:	data_out=16'h881b;
17'h121e3:	data_out=16'h895f;
17'h121e4:	data_out=16'h89ff;
17'h121e5:	data_out=16'h887;
17'h121e6:	data_out=16'ha00;
17'h121e7:	data_out=16'ha00;
17'h121e8:	data_out=16'h9fd;
17'h121e9:	data_out=16'h8a00;
17'h121ea:	data_out=16'h9fc;
17'h121eb:	data_out=16'ha00;
17'h121ec:	data_out=16'h873d;
17'h121ed:	data_out=16'h8962;
17'h121ee:	data_out=16'h9fc;
17'h121ef:	data_out=16'ha00;
17'h121f0:	data_out=16'h9fc;
17'h121f1:	data_out=16'h8998;
17'h121f2:	data_out=16'h8761;
17'h121f3:	data_out=16'ha00;
17'h121f4:	data_out=16'h9fe;
17'h121f5:	data_out=16'h9ff;
17'h121f6:	data_out=16'ha00;
17'h121f7:	data_out=16'h889d;
17'h121f8:	data_out=16'h92d;
17'h121f9:	data_out=16'h8247;
17'h121fa:	data_out=16'h8873;
17'h121fb:	data_out=16'h9fd;
17'h121fc:	data_out=16'h89f2;
17'h121fd:	data_out=16'h2df;
17'h121fe:	data_out=16'h89f2;
17'h121ff:	data_out=16'h5ba;
17'h12200:	data_out=16'h89ca;
17'h12201:	data_out=16'h8963;
17'h12202:	data_out=16'h89d4;
17'h12203:	data_out=16'h89a2;
17'h12204:	data_out=16'ha00;
17'h12205:	data_out=16'ha00;
17'h12206:	data_out=16'h89f7;
17'h12207:	data_out=16'h8693;
17'h12208:	data_out=16'h89f6;
17'h12209:	data_out=16'h89f2;
17'h1220a:	data_out=16'h9ed;
17'h1220b:	data_out=16'h89e0;
17'h1220c:	data_out=16'h89f2;
17'h1220d:	data_out=16'h89f8;
17'h1220e:	data_out=16'h9fe;
17'h1220f:	data_out=16'h89ec;
17'h12210:	data_out=16'h89e6;
17'h12211:	data_out=16'h4e6;
17'h12212:	data_out=16'h89fb;
17'h12213:	data_out=16'h89e7;
17'h12214:	data_out=16'h895e;
17'h12215:	data_out=16'ha00;
17'h12216:	data_out=16'h8411;
17'h12217:	data_out=16'h8969;
17'h12218:	data_out=16'h89fb;
17'h12219:	data_out=16'ha00;
17'h1221a:	data_out=16'ha00;
17'h1221b:	data_out=16'h8988;
17'h1221c:	data_out=16'h895a;
17'h1221d:	data_out=16'h89f4;
17'h1221e:	data_out=16'h89ab;
17'h1221f:	data_out=16'h87ed;
17'h12220:	data_out=16'h88ea;
17'h12221:	data_out=16'h9fe;
17'h12222:	data_out=16'h88f6;
17'h12223:	data_out=16'h9c1;
17'h12224:	data_out=16'h9c5;
17'h12225:	data_out=16'h88c7;
17'h12226:	data_out=16'h89d3;
17'h12227:	data_out=16'h885b;
17'h12228:	data_out=16'h9fe;
17'h12229:	data_out=16'h9fe;
17'h1222a:	data_out=16'h89f3;
17'h1222b:	data_out=16'ha00;
17'h1222c:	data_out=16'h3e0;
17'h1222d:	data_out=16'h8a00;
17'h1222e:	data_out=16'h89d6;
17'h1222f:	data_out=16'h8934;
17'h12230:	data_out=16'ha00;
17'h12231:	data_out=16'h9fb;
17'h12232:	data_out=16'h9f7;
17'h12233:	data_out=16'h89cf;
17'h12234:	data_out=16'h8a00;
17'h12235:	data_out=16'ha00;
17'h12236:	data_out=16'h89c2;
17'h12237:	data_out=16'h89d2;
17'h12238:	data_out=16'h89fc;
17'h12239:	data_out=16'h89d9;
17'h1223a:	data_out=16'h89dd;
17'h1223b:	data_out=16'ha00;
17'h1223c:	data_out=16'h22e;
17'h1223d:	data_out=16'h87d8;
17'h1223e:	data_out=16'h9fe;
17'h1223f:	data_out=16'ha00;
17'h12240:	data_out=16'h235;
17'h12241:	data_out=16'h87cf;
17'h12242:	data_out=16'h8a00;
17'h12243:	data_out=16'ha00;
17'h12244:	data_out=16'ha00;
17'h12245:	data_out=16'ha00;
17'h12246:	data_out=16'h89c2;
17'h12247:	data_out=16'h89ff;
17'h12248:	data_out=16'h89f6;
17'h12249:	data_out=16'h8528;
17'h1224a:	data_out=16'h8914;
17'h1224b:	data_out=16'h8a00;
17'h1224c:	data_out=16'h8a00;
17'h1224d:	data_out=16'h8857;
17'h1224e:	data_out=16'h8a00;
17'h1224f:	data_out=16'h89ff;
17'h12250:	data_out=16'h1f3;
17'h12251:	data_out=16'h409;
17'h12252:	data_out=16'h9dc;
17'h12253:	data_out=16'h8750;
17'h12254:	data_out=16'h89e0;
17'h12255:	data_out=16'h889d;
17'h12256:	data_out=16'h9e6;
17'h12257:	data_out=16'h86d9;
17'h12258:	data_out=16'h807f;
17'h12259:	data_out=16'h637;
17'h1225a:	data_out=16'h89e1;
17'h1225b:	data_out=16'ha00;
17'h1225c:	data_out=16'h30d;
17'h1225d:	data_out=16'h87f3;
17'h1225e:	data_out=16'h8944;
17'h1225f:	data_out=16'h89fe;
17'h12260:	data_out=16'h8a00;
17'h12261:	data_out=16'ha00;
17'h12262:	data_out=16'h8971;
17'h12263:	data_out=16'h89c3;
17'h12264:	data_out=16'h8a00;
17'h12265:	data_out=16'h2cd;
17'h12266:	data_out=16'ha00;
17'h12267:	data_out=16'ha00;
17'h12268:	data_out=16'h9fe;
17'h12269:	data_out=16'h89fd;
17'h1226a:	data_out=16'h9fe;
17'h1226b:	data_out=16'h342;
17'h1226c:	data_out=16'h893a;
17'h1226d:	data_out=16'h89cd;
17'h1226e:	data_out=16'h9fe;
17'h1226f:	data_out=16'ha00;
17'h12270:	data_out=16'h9fe;
17'h12271:	data_out=16'h89db;
17'h12272:	data_out=16'h376;
17'h12273:	data_out=16'ha00;
17'h12274:	data_out=16'h9ff;
17'h12275:	data_out=16'ha00;
17'h12276:	data_out=16'ha00;
17'h12277:	data_out=16'h89e2;
17'h12278:	data_out=16'h9ce;
17'h12279:	data_out=16'h824c;
17'h1227a:	data_out=16'h898c;
17'h1227b:	data_out=16'h9fe;
17'h1227c:	data_out=16'h89f6;
17'h1227d:	data_out=16'h831c;
17'h1227e:	data_out=16'h8a00;
17'h1227f:	data_out=16'h7da;
17'h12280:	data_out=16'h17f;
17'h12281:	data_out=16'h14f;
17'h12282:	data_out=16'h89f4;
17'h12283:	data_out=16'h89f4;
17'h12284:	data_out=16'ha00;
17'h12285:	data_out=16'ha00;
17'h12286:	data_out=16'h89fe;
17'h12287:	data_out=16'h880a;
17'h12288:	data_out=16'h89f8;
17'h12289:	data_out=16'h89f3;
17'h1228a:	data_out=16'h9fe;
17'h1228b:	data_out=16'h89e2;
17'h1228c:	data_out=16'h89fd;
17'h1228d:	data_out=16'h89fb;
17'h1228e:	data_out=16'ha00;
17'h1228f:	data_out=16'h89f5;
17'h12290:	data_out=16'h89e4;
17'h12291:	data_out=16'h9fb;
17'h12292:	data_out=16'h89fc;
17'h12293:	data_out=16'h89f6;
17'h12294:	data_out=16'h89f1;
17'h12295:	data_out=16'ha00;
17'h12296:	data_out=16'h89b2;
17'h12297:	data_out=16'h89f8;
17'h12298:	data_out=16'h89fb;
17'h12299:	data_out=16'ha00;
17'h1229a:	data_out=16'ha00;
17'h1229b:	data_out=16'h89f3;
17'h1229c:	data_out=16'h8825;
17'h1229d:	data_out=16'h83cd;
17'h1229e:	data_out=16'h89ec;
17'h1229f:	data_out=16'h8980;
17'h122a0:	data_out=16'h85a3;
17'h122a1:	data_out=16'ha00;
17'h122a2:	data_out=16'ha00;
17'h122a3:	data_out=16'h9f8;
17'h122a4:	data_out=16'h9f8;
17'h122a5:	data_out=16'h84b7;
17'h122a6:	data_out=16'h89ac;
17'h122a7:	data_out=16'h8298;
17'h122a8:	data_out=16'ha00;
17'h122a9:	data_out=16'h9fe;
17'h122aa:	data_out=16'h89f5;
17'h122ab:	data_out=16'ha00;
17'h122ac:	data_out=16'h1c9;
17'h122ad:	data_out=16'h8a00;
17'h122ae:	data_out=16'h89f8;
17'h122af:	data_out=16'h89f3;
17'h122b0:	data_out=16'h9fe;
17'h122b1:	data_out=16'h9fa;
17'h122b2:	data_out=16'ha00;
17'h122b3:	data_out=16'h89f5;
17'h122b4:	data_out=16'h89fe;
17'h122b5:	data_out=16'ha00;
17'h122b6:	data_out=16'h89e8;
17'h122b7:	data_out=16'h89ee;
17'h122b8:	data_out=16'h8903;
17'h122b9:	data_out=16'h89f5;
17'h122ba:	data_out=16'h89e3;
17'h122bb:	data_out=16'ha00;
17'h122bc:	data_out=16'h8900;
17'h122bd:	data_out=16'h9f7;
17'h122be:	data_out=16'ha00;
17'h122bf:	data_out=16'ha00;
17'h122c0:	data_out=16'ha00;
17'h122c1:	data_out=16'h899d;
17'h122c2:	data_out=16'h89ff;
17'h122c3:	data_out=16'h1f8;
17'h122c4:	data_out=16'ha00;
17'h122c5:	data_out=16'ha00;
17'h122c6:	data_out=16'h8812;
17'h122c7:	data_out=16'h89fc;
17'h122c8:	data_out=16'h89fa;
17'h122c9:	data_out=16'h15b;
17'h122ca:	data_out=16'h89de;
17'h122cb:	data_out=16'h8a00;
17'h122cc:	data_out=16'h89e1;
17'h122cd:	data_out=16'ha00;
17'h122ce:	data_out=16'h89ff;
17'h122cf:	data_out=16'h89b4;
17'h122d0:	data_out=16'h1c0;
17'h122d1:	data_out=16'h89eb;
17'h122d2:	data_out=16'h9fb;
17'h122d3:	data_out=16'h88b5;
17'h122d4:	data_out=16'h89ee;
17'h122d5:	data_out=16'h89bc;
17'h122d6:	data_out=16'h9fa;
17'h122d7:	data_out=16'h9ff;
17'h122d8:	data_out=16'h89f9;
17'h122d9:	data_out=16'h9d3;
17'h122da:	data_out=16'h89fe;
17'h122db:	data_out=16'ha00;
17'h122dc:	data_out=16'h83b2;
17'h122dd:	data_out=16'h89c6;
17'h122de:	data_out=16'h89f6;
17'h122df:	data_out=16'h89fb;
17'h122e0:	data_out=16'h89d4;
17'h122e1:	data_out=16'ha00;
17'h122e2:	data_out=16'h89f0;
17'h122e3:	data_out=16'h89f5;
17'h122e4:	data_out=16'h89e7;
17'h122e5:	data_out=16'h99e;
17'h122e6:	data_out=16'h9fb;
17'h122e7:	data_out=16'ha00;
17'h122e8:	data_out=16'ha00;
17'h122e9:	data_out=16'h89fc;
17'h122ea:	data_out=16'ha00;
17'h122eb:	data_out=16'h885;
17'h122ec:	data_out=16'h85b5;
17'h122ed:	data_out=16'h89f5;
17'h122ee:	data_out=16'ha00;
17'h122ef:	data_out=16'h425;
17'h122f0:	data_out=16'ha00;
17'h122f1:	data_out=16'h89f6;
17'h122f2:	data_out=16'h92e;
17'h122f3:	data_out=16'ha00;
17'h122f4:	data_out=16'h9fd;
17'h122f5:	data_out=16'h9fa;
17'h122f6:	data_out=16'ha00;
17'h122f7:	data_out=16'h89f4;
17'h122f8:	data_out=16'h87a;
17'h122f9:	data_out=16'h8628;
17'h122fa:	data_out=16'h89f5;
17'h122fb:	data_out=16'ha00;
17'h122fc:	data_out=16'h89fa;
17'h122fd:	data_out=16'h834d;
17'h122fe:	data_out=16'h8a00;
17'h122ff:	data_out=16'h9fd;
17'h12300:	data_out=16'h9fb;
17'h12301:	data_out=16'h9a6;
17'h12302:	data_out=16'h89d0;
17'h12303:	data_out=16'h89e7;
17'h12304:	data_out=16'ha00;
17'h12305:	data_out=16'ha00;
17'h12306:	data_out=16'h89ff;
17'h12307:	data_out=16'h89f3;
17'h12308:	data_out=16'h89fa;
17'h12309:	data_out=16'h8666;
17'h1230a:	data_out=16'ha00;
17'h1230b:	data_out=16'h89fa;
17'h1230c:	data_out=16'h89fe;
17'h1230d:	data_out=16'h89fb;
17'h1230e:	data_out=16'ha00;
17'h1230f:	data_out=16'h89df;
17'h12310:	data_out=16'h1f9;
17'h12311:	data_out=16'h9f8;
17'h12312:	data_out=16'h89fd;
17'h12313:	data_out=16'h89dd;
17'h12314:	data_out=16'h89f8;
17'h12315:	data_out=16'ha00;
17'h12316:	data_out=16'h9e3;
17'h12317:	data_out=16'h89fd;
17'h12318:	data_out=16'h29b;
17'h12319:	data_out=16'h9f7;
17'h1231a:	data_out=16'ha00;
17'h1231b:	data_out=16'h89ee;
17'h1231c:	data_out=16'h933;
17'h1231d:	data_out=16'h6ce;
17'h1231e:	data_out=16'h89d1;
17'h1231f:	data_out=16'h8986;
17'h12320:	data_out=16'ha00;
17'h12321:	data_out=16'ha00;
17'h12322:	data_out=16'ha00;
17'h12323:	data_out=16'h9fc;
17'h12324:	data_out=16'h9fc;
17'h12325:	data_out=16'h92a;
17'h12326:	data_out=16'h88fc;
17'h12327:	data_out=16'h9ec;
17'h12328:	data_out=16'ha00;
17'h12329:	data_out=16'h9fa;
17'h1232a:	data_out=16'h89df;
17'h1232b:	data_out=16'ha00;
17'h1232c:	data_out=16'h9fe;
17'h1232d:	data_out=16'h8a00;
17'h1232e:	data_out=16'h89ff;
17'h1232f:	data_out=16'h89f9;
17'h12330:	data_out=16'h9fb;
17'h12331:	data_out=16'h76c;
17'h12332:	data_out=16'h9f6;
17'h12333:	data_out=16'h89f9;
17'h12334:	data_out=16'h2f4;
17'h12335:	data_out=16'ha00;
17'h12336:	data_out=16'h89d9;
17'h12337:	data_out=16'h89cf;
17'h12338:	data_out=16'h858;
17'h12339:	data_out=16'h89f4;
17'h1233a:	data_out=16'h84d5;
17'h1233b:	data_out=16'ha00;
17'h1233c:	data_out=16'h85c1;
17'h1233d:	data_out=16'ha00;
17'h1233e:	data_out=16'ha00;
17'h1233f:	data_out=16'ha00;
17'h12340:	data_out=16'ha00;
17'h12341:	data_out=16'h89bb;
17'h12342:	data_out=16'h89fe;
17'h12343:	data_out=16'h8476;
17'h12344:	data_out=16'ha00;
17'h12345:	data_out=16'ha00;
17'h12346:	data_out=16'h81c0;
17'h12347:	data_out=16'h89dd;
17'h12348:	data_out=16'h89fe;
17'h12349:	data_out=16'ha00;
17'h1234a:	data_out=16'h89fa;
17'h1234b:	data_out=16'h89ff;
17'h1234c:	data_out=16'h8482;
17'h1234d:	data_out=16'ha00;
17'h1234e:	data_out=16'h880f;
17'h1234f:	data_out=16'h54e;
17'h12350:	data_out=16'h9e6;
17'h12351:	data_out=16'h89de;
17'h12352:	data_out=16'ha00;
17'h12353:	data_out=16'h8890;
17'h12354:	data_out=16'h518;
17'h12355:	data_out=16'h89b6;
17'h12356:	data_out=16'ha00;
17'h12357:	data_out=16'ha00;
17'h12358:	data_out=16'h89ef;
17'h12359:	data_out=16'ha00;
17'h1235a:	data_out=16'h8a00;
17'h1235b:	data_out=16'ha00;
17'h1235c:	data_out=16'h8707;
17'h1235d:	data_out=16'h8372;
17'h1235e:	data_out=16'h89fb;
17'h1235f:	data_out=16'h8977;
17'h12360:	data_out=16'h89d6;
17'h12361:	data_out=16'ha00;
17'h12362:	data_out=16'h89fb;
17'h12363:	data_out=16'h89fb;
17'h12364:	data_out=16'h39f;
17'h12365:	data_out=16'h83a0;
17'h12366:	data_out=16'h9f0;
17'h12367:	data_out=16'ha00;
17'h12368:	data_out=16'ha00;
17'h12369:	data_out=16'h89fc;
17'h1236a:	data_out=16'ha00;
17'h1236b:	data_out=16'h9ea;
17'h1236c:	data_out=16'h9ff;
17'h1236d:	data_out=16'h89fa;
17'h1236e:	data_out=16'ha00;
17'h1236f:	data_out=16'h8495;
17'h12370:	data_out=16'ha00;
17'h12371:	data_out=16'h89fb;
17'h12372:	data_out=16'h9fa;
17'h12373:	data_out=16'ha00;
17'h12374:	data_out=16'h9fc;
17'h12375:	data_out=16'h9ff;
17'h12376:	data_out=16'ha00;
17'h12377:	data_out=16'h3d8;
17'h12378:	data_out=16'h261;
17'h12379:	data_out=16'h84e2;
17'h1237a:	data_out=16'h89fb;
17'h1237b:	data_out=16'ha00;
17'h1237c:	data_out=16'h81c5;
17'h1237d:	data_out=16'h81b8;
17'h1237e:	data_out=16'h8a00;
17'h1237f:	data_out=16'ha00;
17'h12380:	data_out=16'ha00;
17'h12381:	data_out=16'h9d2;
17'h12382:	data_out=16'h89f4;
17'h12383:	data_out=16'h858d;
17'h12384:	data_out=16'ha00;
17'h12385:	data_out=16'h9f9;
17'h12386:	data_out=16'h8a00;
17'h12387:	data_out=16'h88b3;
17'h12388:	data_out=16'h89fc;
17'h12389:	data_out=16'h93d;
17'h1238a:	data_out=16'ha00;
17'h1238b:	data_out=16'h89f9;
17'h1238c:	data_out=16'h8a00;
17'h1238d:	data_out=16'h89fe;
17'h1238e:	data_out=16'ha00;
17'h1238f:	data_out=16'h89fe;
17'h12390:	data_out=16'ha00;
17'h12391:	data_out=16'h9fd;
17'h12392:	data_out=16'h89fe;
17'h12393:	data_out=16'h830e;
17'h12394:	data_out=16'h89eb;
17'h12395:	data_out=16'ha00;
17'h12396:	data_out=16'h9f3;
17'h12397:	data_out=16'h8a00;
17'h12398:	data_out=16'h9ff;
17'h12399:	data_out=16'h9fd;
17'h1239a:	data_out=16'ha00;
17'h1239b:	data_out=16'h89ff;
17'h1239c:	data_out=16'h9dc;
17'h1239d:	data_out=16'h8ff;
17'h1239e:	data_out=16'h82ef;
17'h1239f:	data_out=16'h4b0;
17'h123a0:	data_out=16'ha00;
17'h123a1:	data_out=16'ha00;
17'h123a2:	data_out=16'ha00;
17'h123a3:	data_out=16'h9d5;
17'h123a4:	data_out=16'h9d4;
17'h123a5:	data_out=16'ha00;
17'h123a6:	data_out=16'h85ed;
17'h123a7:	data_out=16'ha00;
17'h123a8:	data_out=16'ha00;
17'h123a9:	data_out=16'h7af;
17'h123aa:	data_out=16'h89fe;
17'h123ab:	data_out=16'ha00;
17'h123ac:	data_out=16'h9ff;
17'h123ad:	data_out=16'h87cd;
17'h123ae:	data_out=16'h8a00;
17'h123af:	data_out=16'h9ea;
17'h123b0:	data_out=16'h9f3;
17'h123b1:	data_out=16'h307;
17'h123b2:	data_out=16'h9f0;
17'h123b3:	data_out=16'h792;
17'h123b4:	data_out=16'h70b;
17'h123b5:	data_out=16'ha00;
17'h123b6:	data_out=16'h87ec;
17'h123b7:	data_out=16'h89f9;
17'h123b8:	data_out=16'h9fd;
17'h123b9:	data_out=16'h661;
17'h123ba:	data_out=16'ha00;
17'h123bb:	data_out=16'h91f;
17'h123bc:	data_out=16'h89e2;
17'h123bd:	data_out=16'ha00;
17'h123be:	data_out=16'ha00;
17'h123bf:	data_out=16'h9fa;
17'h123c0:	data_out=16'h9ff;
17'h123c1:	data_out=16'h89e8;
17'h123c2:	data_out=16'h8a00;
17'h123c3:	data_out=16'h888a;
17'h123c4:	data_out=16'ha00;
17'h123c5:	data_out=16'ha00;
17'h123c6:	data_out=16'h86d6;
17'h123c7:	data_out=16'h435;
17'h123c8:	data_out=16'h89ff;
17'h123c9:	data_out=16'ha00;
17'h123ca:	data_out=16'h89fd;
17'h123cb:	data_out=16'h8a00;
17'h123cc:	data_out=16'h82b8;
17'h123cd:	data_out=16'ha00;
17'h123ce:	data_out=16'h854a;
17'h123cf:	data_out=16'h9fe;
17'h123d0:	data_out=16'h9f8;
17'h123d1:	data_out=16'h82a1;
17'h123d2:	data_out=16'ha00;
17'h123d3:	data_out=16'h873e;
17'h123d4:	data_out=16'ha00;
17'h123d5:	data_out=16'h8543;
17'h123d6:	data_out=16'ha00;
17'h123d7:	data_out=16'ha00;
17'h123d8:	data_out=16'h84c1;
17'h123d9:	data_out=16'ha00;
17'h123da:	data_out=16'h8a00;
17'h123db:	data_out=16'ha00;
17'h123dc:	data_out=16'h837;
17'h123dd:	data_out=16'h9fc;
17'h123de:	data_out=16'h9c7;
17'h123df:	data_out=16'ha00;
17'h123e0:	data_out=16'h89ff;
17'h123e1:	data_out=16'h9fd;
17'h123e2:	data_out=16'h89ff;
17'h123e3:	data_out=16'hd5;
17'h123e4:	data_out=16'ha00;
17'h123e5:	data_out=16'h83b7;
17'h123e6:	data_out=16'h9f6;
17'h123e7:	data_out=16'ha00;
17'h123e8:	data_out=16'ha00;
17'h123e9:	data_out=16'h89fe;
17'h123ea:	data_out=16'ha00;
17'h123eb:	data_out=16'ha00;
17'h123ec:	data_out=16'ha00;
17'h123ed:	data_out=16'h3a7;
17'h123ee:	data_out=16'ha00;
17'h123ef:	data_out=16'h89ff;
17'h123f0:	data_out=16'ha00;
17'h123f1:	data_out=16'h89fe;
17'h123f2:	data_out=16'ha00;
17'h123f3:	data_out=16'ha00;
17'h123f4:	data_out=16'h9ed;
17'h123f5:	data_out=16'h898f;
17'h123f6:	data_out=16'ha00;
17'h123f7:	data_out=16'h9cb;
17'h123f8:	data_out=16'h851d;
17'h123f9:	data_out=16'h8466;
17'h123fa:	data_out=16'h89f9;
17'h123fb:	data_out=16'ha00;
17'h123fc:	data_out=16'h9ff;
17'h123fd:	data_out=16'h11b;
17'h123fe:	data_out=16'h5f9;
17'h123ff:	data_out=16'ha00;
17'h12400:	data_out=16'ha00;
17'h12401:	data_out=16'h9dd;
17'h12402:	data_out=16'h89f6;
17'h12403:	data_out=16'h9fc;
17'h12404:	data_out=16'h9ff;
17'h12405:	data_out=16'h979;
17'h12406:	data_out=16'h7fe;
17'h12407:	data_out=16'h8172;
17'h12408:	data_out=16'h89d5;
17'h12409:	data_out=16'h9f4;
17'h1240a:	data_out=16'h9fe;
17'h1240b:	data_out=16'h1fd;
17'h1240c:	data_out=16'h8a00;
17'h1240d:	data_out=16'h81bb;
17'h1240e:	data_out=16'h34b;
17'h1240f:	data_out=16'h86aa;
17'h12410:	data_out=16'ha00;
17'h12411:	data_out=16'h9fe;
17'h12412:	data_out=16'h89c7;
17'h12413:	data_out=16'h9fc;
17'h12414:	data_out=16'h9f2;
17'h12415:	data_out=16'ha00;
17'h12416:	data_out=16'ha00;
17'h12417:	data_out=16'h3bc;
17'h12418:	data_out=16'h98f;
17'h12419:	data_out=16'h9fa;
17'h1241a:	data_out=16'h9fb;
17'h1241b:	data_out=16'h89e0;
17'h1241c:	data_out=16'h9ff;
17'h1241d:	data_out=16'h9cf;
17'h1241e:	data_out=16'h9fb;
17'h1241f:	data_out=16'h9f1;
17'h12420:	data_out=16'ha00;
17'h12421:	data_out=16'h30d;
17'h12422:	data_out=16'ha00;
17'h12423:	data_out=16'h82bc;
17'h12424:	data_out=16'h82b9;
17'h12425:	data_out=16'ha00;
17'h12426:	data_out=16'h9ee;
17'h12427:	data_out=16'h9f4;
17'h12428:	data_out=16'h2db;
17'h12429:	data_out=16'h9fa;
17'h1242a:	data_out=16'h8159;
17'h1242b:	data_out=16'h9fd;
17'h1242c:	data_out=16'ha00;
17'h1242d:	data_out=16'h9fb;
17'h1242e:	data_out=16'h83d8;
17'h1242f:	data_out=16'h9f2;
17'h12430:	data_out=16'h89fe;
17'h12431:	data_out=16'h9ed;
17'h12432:	data_out=16'h8a00;
17'h12433:	data_out=16'h9f5;
17'h12434:	data_out=16'h9a5;
17'h12435:	data_out=16'h802;
17'h12436:	data_out=16'h396;
17'h12437:	data_out=16'h89fc;
17'h12438:	data_out=16'ha00;
17'h12439:	data_out=16'h9fb;
17'h1243a:	data_out=16'ha00;
17'h1243b:	data_out=16'h4f9;
17'h1243c:	data_out=16'h88a1;
17'h1243d:	data_out=16'ha00;
17'h1243e:	data_out=16'h2d9;
17'h1243f:	data_out=16'h98b;
17'h12440:	data_out=16'h9f7;
17'h12441:	data_out=16'h8434;
17'h12442:	data_out=16'h8551;
17'h12443:	data_out=16'h726;
17'h12444:	data_out=16'h9f9;
17'h12445:	data_out=16'ha00;
17'h12446:	data_out=16'h89f3;
17'h12447:	data_out=16'h9fc;
17'h12448:	data_out=16'h45a;
17'h12449:	data_out=16'ha00;
17'h1244a:	data_out=16'h8a00;
17'h1244b:	data_out=16'h89ff;
17'h1244c:	data_out=16'h9fc;
17'h1244d:	data_out=16'ha00;
17'h1244e:	data_out=16'h841c;
17'h1244f:	data_out=16'h9fd;
17'h12450:	data_out=16'h9fd;
17'h12451:	data_out=16'h9f5;
17'h12452:	data_out=16'h942;
17'h12453:	data_out=16'h89a5;
17'h12454:	data_out=16'h9fe;
17'h12455:	data_out=16'h83b2;
17'h12456:	data_out=16'h9ff;
17'h12457:	data_out=16'ha00;
17'h12458:	data_out=16'h89d8;
17'h12459:	data_out=16'h9fd;
17'h1245a:	data_out=16'h8a00;
17'h1245b:	data_out=16'ha00;
17'h1245c:	data_out=16'h73b;
17'h1245d:	data_out=16'ha00;
17'h1245e:	data_out=16'h9f1;
17'h1245f:	data_out=16'ha00;
17'h12460:	data_out=16'h39c;
17'h12461:	data_out=16'h9f9;
17'h12462:	data_out=16'h84e3;
17'h12463:	data_out=16'h9ef;
17'h12464:	data_out=16'ha00;
17'h12465:	data_out=16'h8af;
17'h12466:	data_out=16'h999;
17'h12467:	data_out=16'h9ff;
17'h12468:	data_out=16'h300;
17'h12469:	data_out=16'h89f3;
17'h1246a:	data_out=16'h378;
17'h1246b:	data_out=16'ha00;
17'h1246c:	data_out=16'ha00;
17'h1246d:	data_out=16'h9f0;
17'h1246e:	data_out=16'h376;
17'h1246f:	data_out=16'h4fb;
17'h12470:	data_out=16'h358;
17'h12471:	data_out=16'h8a00;
17'h12472:	data_out=16'ha00;
17'h12473:	data_out=16'h9fe;
17'h12474:	data_out=16'h8a00;
17'h12475:	data_out=16'h89ff;
17'h12476:	data_out=16'h9fe;
17'h12477:	data_out=16'h9fa;
17'h12478:	data_out=16'h211;
17'h12479:	data_out=16'h8120;
17'h1247a:	data_out=16'h9ee;
17'h1247b:	data_out=16'h2d5;
17'h1247c:	data_out=16'h557;
17'h1247d:	data_out=16'h9ff;
17'h1247e:	data_out=16'h9e6;
17'h1247f:	data_out=16'ha00;
17'h12480:	data_out=16'ha00;
17'h12481:	data_out=16'h28b;
17'h12482:	data_out=16'h8524;
17'h12483:	data_out=16'ha00;
17'h12484:	data_out=16'h9d5;
17'h12485:	data_out=16'h9a8;
17'h12486:	data_out=16'h916;
17'h12487:	data_out=16'h6ec;
17'h12488:	data_out=16'h8979;
17'h12489:	data_out=16'h9ff;
17'h1248a:	data_out=16'h32d;
17'h1248b:	data_out=16'h857c;
17'h1248c:	data_out=16'h8a00;
17'h1248d:	data_out=16'h6a9;
17'h1248e:	data_out=16'hfb;
17'h1248f:	data_out=16'h82c8;
17'h12490:	data_out=16'ha00;
17'h12491:	data_out=16'h3dc;
17'h12492:	data_out=16'h8201;
17'h12493:	data_out=16'ha00;
17'h12494:	data_out=16'ha00;
17'h12495:	data_out=16'ha00;
17'h12496:	data_out=16'ha00;
17'h12497:	data_out=16'h69d;
17'h12498:	data_out=16'h2eb;
17'h12499:	data_out=16'h379;
17'h1249a:	data_out=16'h770;
17'h1249b:	data_out=16'h8150;
17'h1249c:	data_out=16'ha00;
17'h1249d:	data_out=16'h6d1;
17'h1249e:	data_out=16'ha00;
17'h1249f:	data_out=16'h9fe;
17'h124a0:	data_out=16'ha00;
17'h124a1:	data_out=16'hf1;
17'h124a2:	data_out=16'h9fe;
17'h124a3:	data_out=16'h86a9;
17'h124a4:	data_out=16'h86a8;
17'h124a5:	data_out=16'ha00;
17'h124a6:	data_out=16'h7e5;
17'h124a7:	data_out=16'h855;
17'h124a8:	data_out=16'hf0;
17'h124a9:	data_out=16'h9f7;
17'h124aa:	data_out=16'h847a;
17'h124ab:	data_out=16'ha00;
17'h124ac:	data_out=16'ha00;
17'h124ad:	data_out=16'h5da;
17'h124ae:	data_out=16'h81ba;
17'h124af:	data_out=16'ha00;
17'h124b0:	data_out=16'h8817;
17'h124b1:	data_out=16'h47e;
17'h124b2:	data_out=16'h878c;
17'h124b3:	data_out=16'ha00;
17'h124b4:	data_out=16'h8fe;
17'h124b5:	data_out=16'h84cc;
17'h124b6:	data_out=16'h8044;
17'h124b7:	data_out=16'h8531;
17'h124b8:	data_out=16'ha00;
17'h124b9:	data_out=16'ha00;
17'h124ba:	data_out=16'ha00;
17'h124bb:	data_out=16'h6e8;
17'h124bc:	data_out=16'h8911;
17'h124bd:	data_out=16'ha00;
17'h124be:	data_out=16'hf0;
17'h124bf:	data_out=16'h9ad;
17'h124c0:	data_out=16'h9fe;
17'h124c1:	data_out=16'h83c4;
17'h124c2:	data_out=16'h87b2;
17'h124c3:	data_out=16'h921;
17'h124c4:	data_out=16'ha00;
17'h124c5:	data_out=16'ha00;
17'h124c6:	data_out=16'h82a5;
17'h124c7:	data_out=16'ha00;
17'h124c8:	data_out=16'h419;
17'h124c9:	data_out=16'ha00;
17'h124ca:	data_out=16'h179;
17'h124cb:	data_out=16'h8a00;
17'h124cc:	data_out=16'h6d9;
17'h124cd:	data_out=16'h9fe;
17'h124ce:	data_out=16'h8720;
17'h124cf:	data_out=16'h9fd;
17'h124d0:	data_out=16'ha00;
17'h124d1:	data_out=16'h589;
17'h124d2:	data_out=16'h8388;
17'h124d3:	data_out=16'h838f;
17'h124d4:	data_out=16'ha00;
17'h124d5:	data_out=16'h8213;
17'h124d6:	data_out=16'h9fd;
17'h124d7:	data_out=16'ha00;
17'h124d8:	data_out=16'h8736;
17'h124d9:	data_out=16'ha00;
17'h124da:	data_out=16'h8a00;
17'h124db:	data_out=16'h621;
17'h124dc:	data_out=16'h191;
17'h124dd:	data_out=16'h71f;
17'h124de:	data_out=16'ha00;
17'h124df:	data_out=16'h3ff;
17'h124e0:	data_out=16'h8234;
17'h124e1:	data_out=16'h9df;
17'h124e2:	data_out=16'h86cd;
17'h124e3:	data_out=16'ha00;
17'h124e4:	data_out=16'ha00;
17'h124e5:	data_out=16'h90e;
17'h124e6:	data_out=16'h48f;
17'h124e7:	data_out=16'h79e;
17'h124e8:	data_out=16'hf2;
17'h124e9:	data_out=16'h89cf;
17'h124ea:	data_out=16'h102;
17'h124eb:	data_out=16'ha00;
17'h124ec:	data_out=16'h577;
17'h124ed:	data_out=16'ha00;
17'h124ee:	data_out=16'h101;
17'h124ef:	data_out=16'h879;
17'h124f0:	data_out=16'hfc;
17'h124f1:	data_out=16'h89f6;
17'h124f2:	data_out=16'ha00;
17'h124f3:	data_out=16'ha00;
17'h124f4:	data_out=16'h8890;
17'h124f5:	data_out=16'h8a00;
17'h124f6:	data_out=16'ha00;
17'h124f7:	data_out=16'h9fe;
17'h124f8:	data_out=16'h748;
17'h124f9:	data_out=16'h8540;
17'h124fa:	data_out=16'h9ff;
17'h124fb:	data_out=16'hef;
17'h124fc:	data_out=16'h176;
17'h124fd:	data_out=16'h72c;
17'h124fe:	data_out=16'ha00;
17'h124ff:	data_out=16'ha00;
17'h12500:	data_out=16'h60f;
17'h12501:	data_out=16'h30d;
17'h12502:	data_out=16'h59;
17'h12503:	data_out=16'h45b;
17'h12504:	data_out=16'h2c9;
17'h12505:	data_out=16'h36d;
17'h12506:	data_out=16'h1bf;
17'h12507:	data_out=16'h418;
17'h12508:	data_out=16'h80c8;
17'h12509:	data_out=16'h645;
17'h1250a:	data_out=16'h2e5;
17'h1250b:	data_out=16'h11a;
17'h1250c:	data_out=16'h8202;
17'h1250d:	data_out=16'h229;
17'h1250e:	data_out=16'h82;
17'h1250f:	data_out=16'h1e7;
17'h12510:	data_out=16'h397;
17'h12511:	data_out=16'h3bc;
17'h12512:	data_out=16'h211;
17'h12513:	data_out=16'h44a;
17'h12514:	data_out=16'h302;
17'h12515:	data_out=16'h298;
17'h12516:	data_out=16'h260;
17'h12517:	data_out=16'h25d;
17'h12518:	data_out=16'h129;
17'h12519:	data_out=16'h191;
17'h1251a:	data_out=16'h270;
17'h1251b:	data_out=16'h2f5;
17'h1251c:	data_out=16'h51e;
17'h1251d:	data_out=16'h435;
17'h1251e:	data_out=16'h361;
17'h1251f:	data_out=16'h40e;
17'h12520:	data_out=16'h87c;
17'h12521:	data_out=16'h8c;
17'h12522:	data_out=16'h5e7;
17'h12523:	data_out=16'h8224;
17'h12524:	data_out=16'h8224;
17'h12525:	data_out=16'h3e7;
17'h12526:	data_out=16'h329;
17'h12527:	data_out=16'h409;
17'h12528:	data_out=16'hb3;
17'h12529:	data_out=16'h377;
17'h1252a:	data_out=16'h1db;
17'h1252b:	data_out=16'h483;
17'h1252c:	data_out=16'h2a5;
17'h1252d:	data_out=16'h113;
17'h1252e:	data_out=16'h1c9;
17'h1252f:	data_out=16'h4ff;
17'h12530:	data_out=16'h8a;
17'h12531:	data_out=16'h563;
17'h12532:	data_out=16'hc5;
17'h12533:	data_out=16'h3bb;
17'h12534:	data_out=16'h509;
17'h12535:	data_out=16'h8009;
17'h12536:	data_out=16'h27;
17'h12537:	data_out=16'hee;
17'h12538:	data_out=16'h632;
17'h12539:	data_out=16'h3a4;
17'h1253a:	data_out=16'h4dd;
17'h1253b:	data_out=16'h2dc;
17'h1253c:	data_out=16'h8190;
17'h1253d:	data_out=16'h8c7;
17'h1253e:	data_out=16'haf;
17'h1253f:	data_out=16'h354;
17'h12540:	data_out=16'h44b;
17'h12541:	data_out=16'h808b;
17'h12542:	data_out=16'h80cf;
17'h12543:	data_out=16'h1b9;
17'h12544:	data_out=16'h458;
17'h12545:	data_out=16'h2a0;
17'h12546:	data_out=16'h9b;
17'h12547:	data_out=16'h47d;
17'h12548:	data_out=16'h37c;
17'h12549:	data_out=16'h42c;
17'h1254a:	data_out=16'h1d6;
17'h1254b:	data_out=16'h834b;
17'h1254c:	data_out=16'h201;
17'h1254d:	data_out=16'h5e6;
17'h1254e:	data_out=16'h1cc;
17'h1254f:	data_out=16'h238;
17'h12550:	data_out=16'h41b;
17'h12551:	data_out=16'h64;
17'h12552:	data_out=16'h80af;
17'h12553:	data_out=16'h482;
17'h12554:	data_out=16'h5a6;
17'h12555:	data_out=16'h820c;
17'h12556:	data_out=16'h49c;
17'h12557:	data_out=16'h486;
17'h12558:	data_out=16'h828e;
17'h12559:	data_out=16'h405;
17'h1255a:	data_out=16'h803c;
17'h1255b:	data_out=16'h215;
17'h1255c:	data_out=16'h21e;
17'h1255d:	data_out=16'h2e9;
17'h1255e:	data_out=16'h504;
17'h1255f:	data_out=16'h1d0;
17'h12560:	data_out=16'h22f;
17'h12561:	data_out=16'h49f;
17'h12562:	data_out=16'h804a;
17'h12563:	data_out=16'h397;
17'h12564:	data_out=16'h68a;
17'h12565:	data_out=16'h3de;
17'h12566:	data_out=16'h1fb;
17'h12567:	data_out=16'h2fc;
17'h12568:	data_out=16'h9d;
17'h12569:	data_out=16'h813a;
17'h1256a:	data_out=16'h6b;
17'h1256b:	data_out=16'h4e3;
17'h1256c:	data_out=16'h1c3;
17'h1256d:	data_out=16'h3ad;
17'h1256e:	data_out=16'h61;
17'h1256f:	data_out=16'h331;
17'h12570:	data_out=16'h85;
17'h12571:	data_out=16'h125;
17'h12572:	data_out=16'h49e;
17'h12573:	data_out=16'h643;
17'h12574:	data_out=16'h68;
17'h12575:	data_out=16'h822a;
17'h12576:	data_out=16'h3a2;
17'h12577:	data_out=16'h464;
17'h12578:	data_out=16'h208;
17'h12579:	data_out=16'h174;
17'h1257a:	data_out=16'h33d;
17'h1257b:	data_out=16'hbb;
17'h1257c:	data_out=16'h104;
17'h1257d:	data_out=16'h253;
17'h1257e:	data_out=16'h6a8;
17'h1257f:	data_out=16'h398;
17'h12580:	data_out=16'hf;
17'h12581:	data_out=16'ha;
17'h12582:	data_out=16'ha;
17'h12583:	data_out=16'h19;
17'h12584:	data_out=16'h1d;
17'h12585:	data_out=16'h11;
17'h12586:	data_out=16'h9;
17'h12587:	data_out=16'h1a;
17'h12588:	data_out=16'h5;
17'h12589:	data_out=16'h13;
17'h1258a:	data_out=16'hb;
17'h1258b:	data_out=16'h11;
17'h1258c:	data_out=16'h18;
17'h1258d:	data_out=16'he;
17'h1258e:	data_out=16'h2;
17'h1258f:	data_out=16'hd;
17'h12590:	data_out=16'hb;
17'h12591:	data_out=16'h13;
17'h12592:	data_out=16'h19;
17'h12593:	data_out=16'hf;
17'h12594:	data_out=16'h18;
17'h12595:	data_out=16'he;
17'h12596:	data_out=16'h1b;
17'h12597:	data_out=16'hf;
17'h12598:	data_out=16'h8;
17'h12599:	data_out=16'h5;
17'h1259a:	data_out=16'h10;
17'h1259b:	data_out=16'h1a;
17'h1259c:	data_out=16'h5;
17'h1259d:	data_out=16'hb;
17'h1259e:	data_out=16'h14;
17'h1259f:	data_out=16'h19;
17'h125a0:	data_out=16'hc;
17'h125a1:	data_out=16'hb;
17'h125a2:	data_out=16'h12;
17'h125a3:	data_out=16'h0;
17'h125a4:	data_out=16'h3;
17'h125a5:	data_out=16'h1e;
17'h125a6:	data_out=16'h17;
17'h125a7:	data_out=16'h10;
17'h125a8:	data_out=16'hc;
17'h125a9:	data_out=16'hb;
17'h125aa:	data_out=16'h19;
17'h125ab:	data_out=16'h9;
17'h125ac:	data_out=16'h13;
17'h125ad:	data_out=16'h1e;
17'h125ae:	data_out=16'h20;
17'h125af:	data_out=16'h19;
17'h125b0:	data_out=16'h14;
17'h125b1:	data_out=16'h11;
17'h125b2:	data_out=16'hc;
17'h125b3:	data_out=16'hf;
17'h125b4:	data_out=16'he;
17'h125b5:	data_out=16'h24;
17'h125b6:	data_out=16'h11;
17'h125b7:	data_out=16'h13;
17'h125b8:	data_out=16'h2;
17'h125b9:	data_out=16'h12;
17'h125ba:	data_out=16'h11;
17'h125bb:	data_out=16'h12;
17'h125bc:	data_out=16'h15;
17'h125bd:	data_out=16'ha;
17'h125be:	data_out=16'h4;
17'h125bf:	data_out=16'h1d;
17'h125c0:	data_out=16'h20;
17'h125c1:	data_out=16'h1c;
17'h125c2:	data_out=16'h12;
17'h125c3:	data_out=16'h8;
17'h125c4:	data_out=16'h1f;
17'h125c5:	data_out=16'h8;
17'h125c6:	data_out=16'hd;
17'h125c7:	data_out=16'h1a;
17'h125c8:	data_out=16'he;
17'h125c9:	data_out=16'hf;
17'h125ca:	data_out=16'h15;
17'h125cb:	data_out=16'h1f;
17'h125cc:	data_out=16'h14;
17'h125cd:	data_out=16'h8;
17'h125ce:	data_out=16'h16;
17'h125cf:	data_out=16'h1e;
17'h125d0:	data_out=16'h1e;
17'h125d1:	data_out=16'hf;
17'h125d2:	data_out=16'h8002;
17'h125d3:	data_out=16'h10;
17'h125d4:	data_out=16'h12;
17'h125d5:	data_out=16'h14;
17'h125d6:	data_out=16'h19;
17'h125d7:	data_out=16'ha;
17'h125d8:	data_out=16'he;
17'h125d9:	data_out=16'hf;
17'h125da:	data_out=16'h12;
17'h125db:	data_out=16'h10;
17'h125dc:	data_out=16'hd;
17'h125dd:	data_out=16'h19;
17'h125de:	data_out=16'h1b;
17'h125df:	data_out=16'h8;
17'h125e0:	data_out=16'h1b;
17'h125e1:	data_out=16'h9;
17'h125e2:	data_out=16'hd;
17'h125e3:	data_out=16'h19;
17'h125e4:	data_out=16'h8;
17'h125e5:	data_out=16'h1d;
17'h125e6:	data_out=16'hb;
17'h125e7:	data_out=16'he;
17'h125e8:	data_out=16'h2;
17'h125e9:	data_out=16'h16;
17'h125ea:	data_out=16'hb;
17'h125eb:	data_out=16'h12;
17'h125ec:	data_out=16'h1a;
17'h125ed:	data_out=16'hf;
17'h125ee:	data_out=16'h1;
17'h125ef:	data_out=16'h15;
17'h125f0:	data_out=16'hd;
17'h125f1:	data_out=16'h11;
17'h125f2:	data_out=16'h1d;
17'h125f3:	data_out=16'h12;
17'h125f4:	data_out=16'h1a;
17'h125f5:	data_out=16'h12;
17'h125f6:	data_out=16'hb;
17'h125f7:	data_out=16'h17;
17'h125f8:	data_out=16'h12;
17'h125f9:	data_out=16'h10;
17'h125fa:	data_out=16'hc;
17'h125fb:	data_out=16'h1;
17'h125fc:	data_out=16'h13;
17'h125fd:	data_out=16'h14;
17'h125fe:	data_out=16'he;
17'h125ff:	data_out=16'h1f;
17'h12600:	data_out=16'he;
17'h12601:	data_out=16'ha;
17'h12602:	data_out=16'hc;
17'h12603:	data_out=16'h11;
17'h12604:	data_out=16'hd;
17'h12605:	data_out=16'h2;
17'h12606:	data_out=16'h8002;
17'h12607:	data_out=16'h1;
17'h12608:	data_out=16'h10;
17'h12609:	data_out=16'hf;
17'h1260a:	data_out=16'h7;
17'h1260b:	data_out=16'hf;
17'h1260c:	data_out=16'h4;
17'h1260d:	data_out=16'hd;
17'h1260e:	data_out=16'h4;
17'h1260f:	data_out=16'h0;
17'h12610:	data_out=16'h8000;
17'h12611:	data_out=16'h8;
17'h12612:	data_out=16'ha;
17'h12613:	data_out=16'h8002;
17'h12614:	data_out=16'h3;
17'h12615:	data_out=16'h8004;
17'h12616:	data_out=16'h1;
17'h12617:	data_out=16'h1;
17'h12618:	data_out=16'h8002;
17'h12619:	data_out=16'h8004;
17'h1261a:	data_out=16'h4;
17'h1261b:	data_out=16'h8001;
17'h1261c:	data_out=16'h1;
17'h1261d:	data_out=16'hc;
17'h1261e:	data_out=16'h10;
17'h1261f:	data_out=16'h2;
17'h12620:	data_out=16'h9;
17'h12621:	data_out=16'h5;
17'h12622:	data_out=16'h1;
17'h12623:	data_out=16'h0;
17'h12624:	data_out=16'h9;
17'h12625:	data_out=16'h5;
17'h12626:	data_out=16'h7;
17'h12627:	data_out=16'hf;
17'h12628:	data_out=16'h8001;
17'h12629:	data_out=16'h8002;
17'h1262a:	data_out=16'hf;
17'h1262b:	data_out=16'h6;
17'h1262c:	data_out=16'hf;
17'h1262d:	data_out=16'h4;
17'h1262e:	data_out=16'h10;
17'h1262f:	data_out=16'h10;
17'h12630:	data_out=16'h10;
17'h12631:	data_out=16'h3;
17'h12632:	data_out=16'h10;
17'h12633:	data_out=16'h3;
17'h12634:	data_out=16'h5;
17'h12635:	data_out=16'h4;
17'h12636:	data_out=16'h5;
17'h12637:	data_out=16'h9;
17'h12638:	data_out=16'h8002;
17'h12639:	data_out=16'hb;
17'h1263a:	data_out=16'hb;
17'h1263b:	data_out=16'h9;
17'h1263c:	data_out=16'h7;
17'h1263d:	data_out=16'h8;
17'h1263e:	data_out=16'h8;
17'h1263f:	data_out=16'h8001;
17'h12640:	data_out=16'h4;
17'h12641:	data_out=16'h8001;
17'h12642:	data_out=16'h9;
17'h12643:	data_out=16'h8002;
17'h12644:	data_out=16'h7;
17'h12645:	data_out=16'h8004;
17'h12646:	data_out=16'h8006;
17'h12647:	data_out=16'hd;
17'h12648:	data_out=16'h0;
17'h12649:	data_out=16'hd;
17'h1264a:	data_out=16'h8;
17'h1264b:	data_out=16'h12;
17'h1264c:	data_out=16'h3;
17'h1264d:	data_out=16'h8001;
17'h1264e:	data_out=16'h11;
17'h1264f:	data_out=16'h3;
17'h12650:	data_out=16'ha;
17'h12651:	data_out=16'hd;
17'h12652:	data_out=16'h0;
17'h12653:	data_out=16'h1;
17'h12654:	data_out=16'h8002;
17'h12655:	data_out=16'he;
17'h12656:	data_out=16'hb;
17'h12657:	data_out=16'h6;
17'h12658:	data_out=16'ha;
17'h12659:	data_out=16'h5;
17'h1265a:	data_out=16'h8001;
17'h1265b:	data_out=16'h8004;
17'h1265c:	data_out=16'he;
17'h1265d:	data_out=16'hf;
17'h1265e:	data_out=16'h2;
17'h1265f:	data_out=16'h8001;
17'h12660:	data_out=16'h10;
17'h12661:	data_out=16'hb;
17'h12662:	data_out=16'h2;
17'h12663:	data_out=16'h4;
17'h12664:	data_out=16'ha;
17'h12665:	data_out=16'h4;
17'h12666:	data_out=16'h8005;
17'h12667:	data_out=16'he;
17'h12668:	data_out=16'h8005;
17'h12669:	data_out=16'h6;
17'h1266a:	data_out=16'h6;
17'h1266b:	data_out=16'h3;
17'h1266c:	data_out=16'ha;
17'h1266d:	data_out=16'ha;
17'h1266e:	data_out=16'h1;
17'h1266f:	data_out=16'h8001;
17'h12670:	data_out=16'h3;
17'h12671:	data_out=16'hf;
17'h12672:	data_out=16'h3;
17'h12673:	data_out=16'h7;
17'h12674:	data_out=16'ha;
17'h12675:	data_out=16'hd;
17'h12676:	data_out=16'h8002;
17'h12677:	data_out=16'h6;
17'h12678:	data_out=16'h1;
17'h12679:	data_out=16'h5;
17'h1267a:	data_out=16'h6;
17'h1267b:	data_out=16'h8002;
17'h1267c:	data_out=16'h8005;
17'h1267d:	data_out=16'h7;
17'h1267e:	data_out=16'h6;
17'h1267f:	data_out=16'h12;
17'h12680:	data_out=16'h8002;
17'h12681:	data_out=16'h62;
17'h12682:	data_out=16'h84;
17'h12683:	data_out=16'h85;
17'h12684:	data_out=16'h6a;
17'h12685:	data_out=16'h95;
17'h12686:	data_out=16'h80;
17'h12687:	data_out=16'h87;
17'h12688:	data_out=16'h58;
17'h12689:	data_out=16'h51;
17'h1268a:	data_out=16'h56;
17'h1268b:	data_out=16'h6d;
17'h1268c:	data_out=16'h6a;
17'h1268d:	data_out=16'h71;
17'h1268e:	data_out=16'h32;
17'h1268f:	data_out=16'h8c;
17'h12690:	data_out=16'h8f;
17'h12691:	data_out=16'h76;
17'h12692:	data_out=16'hb5;
17'h12693:	data_out=16'h95;
17'h12694:	data_out=16'hba;
17'h12695:	data_out=16'h47;
17'h12696:	data_out=16'h6b;
17'h12697:	data_out=16'hb0;
17'h12698:	data_out=16'h57;
17'h12699:	data_out=16'h30;
17'h1269a:	data_out=16'h6d;
17'h1269b:	data_out=16'h80;
17'h1269c:	data_out=16'h88;
17'h1269d:	data_out=16'h68;
17'h1269e:	data_out=16'h9b;
17'h1269f:	data_out=16'h9d;
17'h126a0:	data_out=16'h76;
17'h126a1:	data_out=16'h3c;
17'h126a2:	data_out=16'h79;
17'h126a3:	data_out=16'h20;
17'h126a4:	data_out=16'h19;
17'h126a5:	data_out=16'h97;
17'h126a6:	data_out=16'h53;
17'h126a7:	data_out=16'h6c;
17'h126a8:	data_out=16'h36;
17'h126a9:	data_out=16'h80;
17'h126aa:	data_out=16'ha4;
17'h126ab:	data_out=16'h45;
17'h126ac:	data_out=16'h6c;
17'h126ad:	data_out=16'h5b;
17'h126ae:	data_out=16'hd3;
17'h126af:	data_out=16'h96;
17'h126b0:	data_out=16'haf;
17'h126b1:	data_out=16'h4b;
17'h126b2:	data_out=16'hb0;
17'h126b3:	data_out=16'ha9;
17'h126b4:	data_out=16'h51;
17'h126b5:	data_out=16'h91;
17'h126b6:	data_out=16'h73;
17'h126b7:	data_out=16'h94;
17'h126b8:	data_out=16'h5a;
17'h126b9:	data_out=16'h84;
17'h126ba:	data_out=16'h78;
17'h126bb:	data_out=16'h50;
17'h126bc:	data_out=16'h81;
17'h126bd:	data_out=16'h5b;
17'h126be:	data_out=16'h3e;
17'h126bf:	data_out=16'h9c;
17'h126c0:	data_out=16'h9a;
17'h126c1:	data_out=16'h7f;
17'h126c2:	data_out=16'h5c;
17'h126c3:	data_out=16'h77;
17'h126c4:	data_out=16'h79;
17'h126c5:	data_out=16'h5b;
17'h126c6:	data_out=16'h4d;
17'h126c7:	data_out=16'h89;
17'h126c8:	data_out=16'hbb;
17'h126c9:	data_out=16'h8a;
17'h126ca:	data_out=16'hb0;
17'h126cb:	data_out=16'h74;
17'h126cc:	data_out=16'hbf;
17'h126cd:	data_out=16'h6e;
17'h126ce:	data_out=16'ha0;
17'h126cf:	data_out=16'haf;
17'h126d0:	data_out=16'h8d;
17'h126d1:	data_out=16'h6b;
17'h126d2:	data_out=16'h1c;
17'h126d3:	data_out=16'h68;
17'h126d4:	data_out=16'h99;
17'h126d5:	data_out=16'h85;
17'h126d6:	data_out=16'haf;
17'h126d7:	data_out=16'h9e;
17'h126d8:	data_out=16'h84;
17'h126d9:	data_out=16'ha7;
17'h126da:	data_out=16'h85;
17'h126db:	data_out=16'h74;
17'h126dc:	data_out=16'h62;
17'h126dd:	data_out=16'h95;
17'h126de:	data_out=16'ha3;
17'h126df:	data_out=16'h5e;
17'h126e0:	data_out=16'h75;
17'h126e1:	data_out=16'h81;
17'h126e2:	data_out=16'h6f;
17'h126e3:	data_out=16'hb7;
17'h126e4:	data_out=16'h72;
17'h126e5:	data_out=16'h8b;
17'h126e6:	data_out=16'h50;
17'h126e7:	data_out=16'h98;
17'h126e8:	data_out=16'h33;
17'h126e9:	data_out=16'h7b;
17'h126ea:	data_out=16'h2f;
17'h126eb:	data_out=16'h78;
17'h126ec:	data_out=16'h59;
17'h126ed:	data_out=16'hb7;
17'h126ee:	data_out=16'h32;
17'h126ef:	data_out=16'h96;
17'h126f0:	data_out=16'h30;
17'h126f1:	data_out=16'hbe;
17'h126f2:	data_out=16'hbe;
17'h126f3:	data_out=16'h81;
17'h126f4:	data_out=16'hac;
17'h126f5:	data_out=16'h5d;
17'h126f6:	data_out=16'h3c;
17'h126f7:	data_out=16'hab;
17'h126f8:	data_out=16'h6a;
17'h126f9:	data_out=16'he0;
17'h126fa:	data_out=16'hbe;
17'h126fb:	data_out=16'h38;
17'h126fc:	data_out=16'h52;
17'h126fd:	data_out=16'h8d;
17'h126fe:	data_out=16'h62;
17'h126ff:	data_out=16'h9b;
17'h12700:	data_out=16'h877f;
17'h12701:	data_out=16'h25a;
17'h12702:	data_out=16'h140;
17'h12703:	data_out=16'h1ba;
17'h12704:	data_out=16'h3a5;
17'h12705:	data_out=16'h93b;
17'h12706:	data_out=16'h771;
17'h12707:	data_out=16'h2a3;
17'h12708:	data_out=16'h8088;
17'h12709:	data_out=16'h5c;
17'h1270a:	data_out=16'h8a;
17'h1270b:	data_out=16'h72c;
17'h1270c:	data_out=16'h490;
17'h1270d:	data_out=16'h801c;
17'h1270e:	data_out=16'h159;
17'h1270f:	data_out=16'h2df;
17'h12710:	data_out=16'h129;
17'h12711:	data_out=16'h648;
17'h12712:	data_out=16'h3ba;
17'h12713:	data_out=16'h353;
17'h12714:	data_out=16'h56c;
17'h12715:	data_out=16'h80fb;
17'h12716:	data_out=16'h80a8;
17'h12717:	data_out=16'h53f;
17'h12718:	data_out=16'h14;
17'h12719:	data_out=16'h64f;
17'h1271a:	data_out=16'h46a;
17'h1271b:	data_out=16'h7ae;
17'h1271c:	data_out=16'h6a5;
17'h1271d:	data_out=16'h479;
17'h1271e:	data_out=16'h4a4;
17'h1271f:	data_out=16'h519;
17'h12720:	data_out=16'h7fa;
17'h12721:	data_out=16'h167;
17'h12722:	data_out=16'h253;
17'h12723:	data_out=16'h82ea;
17'h12724:	data_out=16'h82ea;
17'h12725:	data_out=16'h313;
17'h12726:	data_out=16'h8230;
17'h12727:	data_out=16'h5d2;
17'h12728:	data_out=16'h18c;
17'h12729:	data_out=16'h824b;
17'h1272a:	data_out=16'h8025;
17'h1272b:	data_out=16'ha00;
17'h1272c:	data_out=16'h807f;
17'h1272d:	data_out=16'h8550;
17'h1272e:	data_out=16'h38e;
17'h1272f:	data_out=16'h796;
17'h12730:	data_out=16'h371;
17'h12731:	data_out=16'h3ff;
17'h12732:	data_out=16'h3c4;
17'h12733:	data_out=16'h56f;
17'h12734:	data_out=16'h314;
17'h12735:	data_out=16'h9d3;
17'h12736:	data_out=16'h1a3;
17'h12737:	data_out=16'h26a;
17'h12738:	data_out=16'h657;
17'h12739:	data_out=16'h54a;
17'h1273a:	data_out=16'h81b1;
17'h1273b:	data_out=16'h26e;
17'h1273c:	data_out=16'h3e0;
17'h1273d:	data_out=16'h478;
17'h1273e:	data_out=16'h18d;
17'h1273f:	data_out=16'h93a;
17'h12740:	data_out=16'h3f0;
17'h12741:	data_out=16'h4d2;
17'h12742:	data_out=16'h8466;
17'h12743:	data_out=16'h588;
17'h12744:	data_out=16'h363;
17'h12745:	data_out=16'h8149;
17'h12746:	data_out=16'h228;
17'h12747:	data_out=16'h80ff;
17'h12748:	data_out=16'h5da;
17'h12749:	data_out=16'h347;
17'h1274a:	data_out=16'h29d;
17'h1274b:	data_out=16'h119;
17'h1274c:	data_out=16'h800e;
17'h1274d:	data_out=16'h26e;
17'h1274e:	data_out=16'h32e;
17'h1274f:	data_out=16'h8001;
17'h12750:	data_out=16'h116;
17'h12751:	data_out=16'h445;
17'h12752:	data_out=16'h8466;
17'h12753:	data_out=16'h879;
17'h12754:	data_out=16'h66f;
17'h12755:	data_out=16'h3c4;
17'h12756:	data_out=16'hc7;
17'h12757:	data_out=16'h98;
17'h12758:	data_out=16'hef;
17'h12759:	data_out=16'h306;
17'h1275a:	data_out=16'h609;
17'h1275b:	data_out=16'h636;
17'h1275c:	data_out=16'h75f;
17'h1275d:	data_out=16'h64;
17'h1275e:	data_out=16'h752;
17'h1275f:	data_out=16'h17;
17'h12760:	data_out=16'h835b;
17'h12761:	data_out=16'h5aa;
17'h12762:	data_out=16'h3c8;
17'h12763:	data_out=16'h5c4;
17'h12764:	data_out=16'h4a4;
17'h12765:	data_out=16'h62b;
17'h12766:	data_out=16'h8e2;
17'h12767:	data_out=16'h3dd;
17'h12768:	data_out=16'h173;
17'h12769:	data_out=16'h8094;
17'h1276a:	data_out=16'h150;
17'h1276b:	data_out=16'h646;
17'h1276c:	data_out=16'h8a00;
17'h1276d:	data_out=16'h5ab;
17'h1276e:	data_out=16'h150;
17'h1276f:	data_out=16'h41e;
17'h12770:	data_out=16'h155;
17'h12771:	data_out=16'h2d1;
17'h12772:	data_out=16'h39c;
17'h12773:	data_out=16'h69c;
17'h12774:	data_out=16'h360;
17'h12775:	data_out=16'h5cb;
17'h12776:	data_out=16'h8a9;
17'h12777:	data_out=16'h132;
17'h12778:	data_out=16'h554;
17'h12779:	data_out=16'h2e6;
17'h1277a:	data_out=16'h5cf;
17'h1277b:	data_out=16'h18e;
17'h1277c:	data_out=16'h32;
17'h1277d:	data_out=16'h843;
17'h1277e:	data_out=16'h321;
17'h1277f:	data_out=16'h95;
17'h12780:	data_out=16'h8a00;
17'h12781:	data_out=16'ha00;
17'h12782:	data_out=16'h9fb;
17'h12783:	data_out=16'h86b;
17'h12784:	data_out=16'ha00;
17'h12785:	data_out=16'ha00;
17'h12786:	data_out=16'h9f9;
17'h12787:	data_out=16'h2a1;
17'h12788:	data_out=16'h8561;
17'h12789:	data_out=16'h89fe;
17'h1278a:	data_out=16'h81b6;
17'h1278b:	data_out=16'h9df;
17'h1278c:	data_out=16'h598;
17'h1278d:	data_out=16'h7ed;
17'h1278e:	data_out=16'h365;
17'h1278f:	data_out=16'h9ce;
17'h12790:	data_out=16'h80fa;
17'h12791:	data_out=16'ha00;
17'h12792:	data_out=16'h907;
17'h12793:	data_out=16'h8fb;
17'h12794:	data_out=16'ha00;
17'h12795:	data_out=16'h510;
17'h12796:	data_out=16'hef;
17'h12797:	data_out=16'ha00;
17'h12798:	data_out=16'h78;
17'h12799:	data_out=16'ha00;
17'h1279a:	data_out=16'ha00;
17'h1279b:	data_out=16'ha00;
17'h1279c:	data_out=16'h9fe;
17'h1279d:	data_out=16'h9fd;
17'h1279e:	data_out=16'h9f9;
17'h1279f:	data_out=16'ha00;
17'h127a0:	data_out=16'ha00;
17'h127a1:	data_out=16'h3ab;
17'h127a2:	data_out=16'h8584;
17'h127a3:	data_out=16'h8a00;
17'h127a4:	data_out=16'h8a00;
17'h127a5:	data_out=16'h8444;
17'h127a6:	data_out=16'h8a00;
17'h127a7:	data_out=16'ha00;
17'h127a8:	data_out=16'h46c;
17'h127a9:	data_out=16'h85f5;
17'h127aa:	data_out=16'h89f8;
17'h127ab:	data_out=16'ha00;
17'h127ac:	data_out=16'h3ec;
17'h127ad:	data_out=16'h8a00;
17'h127ae:	data_out=16'h880;
17'h127af:	data_out=16'ha00;
17'h127b0:	data_out=16'h617;
17'h127b1:	data_out=16'ha00;
17'h127b2:	data_out=16'h77c;
17'h127b3:	data_out=16'ha00;
17'h127b4:	data_out=16'h5c0;
17'h127b5:	data_out=16'ha00;
17'h127b6:	data_out=16'h59c;
17'h127b7:	data_out=16'h9f9;
17'h127b8:	data_out=16'ha00;
17'h127b9:	data_out=16'ha00;
17'h127ba:	data_out=16'h89d3;
17'h127bb:	data_out=16'ha00;
17'h127bc:	data_out=16'ha00;
17'h127bd:	data_out=16'h9f3;
17'h127be:	data_out=16'h473;
17'h127bf:	data_out=16'ha00;
17'h127c0:	data_out=16'ha00;
17'h127c1:	data_out=16'h9ff;
17'h127c2:	data_out=16'h8a00;
17'h127c3:	data_out=16'ha00;
17'h127c4:	data_out=16'ha00;
17'h127c5:	data_out=16'h510;
17'h127c6:	data_out=16'h85f5;
17'h127c7:	data_out=16'h8a00;
17'h127c8:	data_out=16'h9fc;
17'h127c9:	data_out=16'h81b1;
17'h127ca:	data_out=16'ha00;
17'h127cb:	data_out=16'h8a00;
17'h127cc:	data_out=16'h8a00;
17'h127cd:	data_out=16'h843c;
17'h127ce:	data_out=16'h5e5;
17'h127cf:	data_out=16'h8a00;
17'h127d0:	data_out=16'h9f4;
17'h127d1:	data_out=16'h9fd;
17'h127d2:	data_out=16'h8a00;
17'h127d3:	data_out=16'ha00;
17'h127d4:	data_out=16'ha00;
17'h127d5:	data_out=16'h9f5;
17'h127d6:	data_out=16'h843e;
17'h127d7:	data_out=16'h856e;
17'h127d8:	data_out=16'ha00;
17'h127d9:	data_out=16'h69f;
17'h127da:	data_out=16'ha00;
17'h127db:	data_out=16'ha00;
17'h127dc:	data_out=16'ha00;
17'h127dd:	data_out=16'h83d3;
17'h127de:	data_out=16'ha00;
17'h127df:	data_out=16'h812a;
17'h127e0:	data_out=16'h8a00;
17'h127e1:	data_out=16'ha00;
17'h127e2:	data_out=16'h9f4;
17'h127e3:	data_out=16'ha00;
17'h127e4:	data_out=16'h6fd;
17'h127e5:	data_out=16'ha00;
17'h127e6:	data_out=16'ha00;
17'h127e7:	data_out=16'h2f9;
17'h127e8:	data_out=16'h3e8;
17'h127e9:	data_out=16'h8937;
17'h127ea:	data_out=16'h338;
17'h127eb:	data_out=16'ha00;
17'h127ec:	data_out=16'h8a00;
17'h127ed:	data_out=16'ha00;
17'h127ee:	data_out=16'h338;
17'h127ef:	data_out=16'ha00;
17'h127f0:	data_out=16'h352;
17'h127f1:	data_out=16'h9fc;
17'h127f2:	data_out=16'h9fb;
17'h127f3:	data_out=16'h9fd;
17'h127f4:	data_out=16'h55f;
17'h127f5:	data_out=16'ha00;
17'h127f6:	data_out=16'ha00;
17'h127f7:	data_out=16'h885;
17'h127f8:	data_out=16'h9f9;
17'h127f9:	data_out=16'h6b8;
17'h127fa:	data_out=16'ha00;
17'h127fb:	data_out=16'h475;
17'h127fc:	data_out=16'h3f8;
17'h127fd:	data_out=16'ha00;
17'h127fe:	data_out=16'h803a;
17'h127ff:	data_out=16'h7de;
17'h12800:	data_out=16'h888d;
17'h12801:	data_out=16'ha00;
17'h12802:	data_out=16'h9ef;
17'h12803:	data_out=16'h83e7;
17'h12804:	data_out=16'ha00;
17'h12805:	data_out=16'h9fd;
17'h12806:	data_out=16'h267;
17'h12807:	data_out=16'h8a00;
17'h12808:	data_out=16'h4ff;
17'h12809:	data_out=16'h8a00;
17'h1280a:	data_out=16'h897;
17'h1280b:	data_out=16'h388;
17'h1280c:	data_out=16'h8a00;
17'h1280d:	data_out=16'h878e;
17'h1280e:	data_out=16'h921;
17'h1280f:	data_out=16'h707;
17'h12810:	data_out=16'h89fe;
17'h12811:	data_out=16'ha00;
17'h12812:	data_out=16'h5b2;
17'h12813:	data_out=16'h9d;
17'h12814:	data_out=16'h9ef;
17'h12815:	data_out=16'h9ff;
17'h12816:	data_out=16'h822f;
17'h12817:	data_out=16'h649;
17'h12818:	data_out=16'h2a5;
17'h12819:	data_out=16'ha00;
17'h1281a:	data_out=16'h9fa;
17'h1281b:	data_out=16'h9f5;
17'h1281c:	data_out=16'h9f3;
17'h1281d:	data_out=16'h9fa;
17'h1281e:	data_out=16'h9f0;
17'h1281f:	data_out=16'h9fc;
17'h12820:	data_out=16'ha00;
17'h12821:	data_out=16'h962;
17'h12822:	data_out=16'h8a00;
17'h12823:	data_out=16'h87c0;
17'h12824:	data_out=16'h87b4;
17'h12825:	data_out=16'h89fb;
17'h12826:	data_out=16'h89fc;
17'h12827:	data_out=16'ha00;
17'h12828:	data_out=16'ha00;
17'h12829:	data_out=16'h89f9;
17'h1282a:	data_out=16'h89fc;
17'h1282b:	data_out=16'ha00;
17'h1282c:	data_out=16'h615;
17'h1282d:	data_out=16'h8a00;
17'h1282e:	data_out=16'h369;
17'h1282f:	data_out=16'h9fc;
17'h12830:	data_out=16'h900;
17'h12831:	data_out=16'ha00;
17'h12832:	data_out=16'ha00;
17'h12833:	data_out=16'h9fb;
17'h12834:	data_out=16'h8b2;
17'h12835:	data_out=16'h9ff;
17'h12836:	data_out=16'h9f9;
17'h12837:	data_out=16'h9ec;
17'h12838:	data_out=16'h9fa;
17'h12839:	data_out=16'h9fb;
17'h1283a:	data_out=16'h89fe;
17'h1283b:	data_out=16'ha00;
17'h1283c:	data_out=16'h9fe;
17'h1283d:	data_out=16'h9f9;
17'h1283e:	data_out=16'ha00;
17'h1283f:	data_out=16'h9fd;
17'h12840:	data_out=16'h721;
17'h12841:	data_out=16'h9ee;
17'h12842:	data_out=16'h8a00;
17'h12843:	data_out=16'h9f6;
17'h12844:	data_out=16'ha00;
17'h12845:	data_out=16'h9ff;
17'h12846:	data_out=16'h801e;
17'h12847:	data_out=16'h89ff;
17'h12848:	data_out=16'h8b3;
17'h12849:	data_out=16'h89fb;
17'h1284a:	data_out=16'h917;
17'h1284b:	data_out=16'h8a00;
17'h1284c:	data_out=16'h8a00;
17'h1284d:	data_out=16'h8a00;
17'h1284e:	data_out=16'h5a5;
17'h1284f:	data_out=16'h8a00;
17'h12850:	data_out=16'h83d;
17'h12851:	data_out=16'h9e2;
17'h12852:	data_out=16'h89ff;
17'h12853:	data_out=16'ha00;
17'h12854:	data_out=16'ha00;
17'h12855:	data_out=16'h59e;
17'h12856:	data_out=16'h52d;
17'h12857:	data_out=16'h811d;
17'h12858:	data_out=16'h9f7;
17'h12859:	data_out=16'h8089;
17'h1285a:	data_out=16'h9e9;
17'h1285b:	data_out=16'ha00;
17'h1285c:	data_out=16'h9fe;
17'h1285d:	data_out=16'h89a9;
17'h1285e:	data_out=16'h9f9;
17'h1285f:	data_out=16'h817b;
17'h12860:	data_out=16'h8a00;
17'h12861:	data_out=16'h9fe;
17'h12862:	data_out=16'hd2;
17'h12863:	data_out=16'h9fc;
17'h12864:	data_out=16'h469;
17'h12865:	data_out=16'h9ef;
17'h12866:	data_out=16'ha00;
17'h12867:	data_out=16'h8075;
17'h12868:	data_out=16'h9b3;
17'h12869:	data_out=16'h8811;
17'h1286a:	data_out=16'h8f2;
17'h1286b:	data_out=16'h9fa;
17'h1286c:	data_out=16'h89c4;
17'h1286d:	data_out=16'h9fc;
17'h1286e:	data_out=16'h8f1;
17'h1286f:	data_out=16'h901;
17'h12870:	data_out=16'h90e;
17'h12871:	data_out=16'h9e3;
17'h12872:	data_out=16'h9ff;
17'h12873:	data_out=16'h9ff;
17'h12874:	data_out=16'h85f;
17'h12875:	data_out=16'h9dd;
17'h12876:	data_out=16'ha00;
17'h12877:	data_out=16'h84dd;
17'h12878:	data_out=16'h7a6;
17'h12879:	data_out=16'h424;
17'h1287a:	data_out=16'h9f8;
17'h1287b:	data_out=16'ha00;
17'h1287c:	data_out=16'ha00;
17'h1287d:	data_out=16'ha00;
17'h1287e:	data_out=16'h8a00;
17'h1287f:	data_out=16'h9f5;
17'h12880:	data_out=16'h873c;
17'h12881:	data_out=16'ha00;
17'h12882:	data_out=16'h6a3;
17'h12883:	data_out=16'h89e7;
17'h12884:	data_out=16'h9f0;
17'h12885:	data_out=16'h9f7;
17'h12886:	data_out=16'h7fe;
17'h12887:	data_out=16'h8a00;
17'h12888:	data_out=16'h335;
17'h12889:	data_out=16'h89fe;
17'h1288a:	data_out=16'h9fe;
17'h1288b:	data_out=16'h28c;
17'h1288c:	data_out=16'h8a00;
17'h1288d:	data_out=16'h89ff;
17'h1288e:	data_out=16'h9fc;
17'h1288f:	data_out=16'h8903;
17'h12890:	data_out=16'h89fc;
17'h12891:	data_out=16'ha00;
17'h12892:	data_out=16'h814;
17'h12893:	data_out=16'ha00;
17'h12894:	data_out=16'h9fe;
17'h12895:	data_out=16'h8b4;
17'h12896:	data_out=16'h89d9;
17'h12897:	data_out=16'h75c;
17'h12898:	data_out=16'h89dc;
17'h12899:	data_out=16'ha00;
17'h1289a:	data_out=16'h9f2;
17'h1289b:	data_out=16'h73f;
17'h1289c:	data_out=16'ha00;
17'h1289d:	data_out=16'ha00;
17'h1289e:	data_out=16'h68d;
17'h1289f:	data_out=16'ha00;
17'h128a0:	data_out=16'ha00;
17'h128a1:	data_out=16'h9fc;
17'h128a2:	data_out=16'h8a00;
17'h128a3:	data_out=16'h9eb;
17'h128a4:	data_out=16'h9ed;
17'h128a5:	data_out=16'h89fc;
17'h128a6:	data_out=16'h89e3;
17'h128a7:	data_out=16'ha00;
17'h128a8:	data_out=16'h9fc;
17'h128a9:	data_out=16'h89e1;
17'h128aa:	data_out=16'h89ef;
17'h128ab:	data_out=16'ha00;
17'h128ac:	data_out=16'h8434;
17'h128ad:	data_out=16'h89eb;
17'h128ae:	data_out=16'h8891;
17'h128af:	data_out=16'ha00;
17'h128b0:	data_out=16'h8a8;
17'h128b1:	data_out=16'ha00;
17'h128b2:	data_out=16'ha00;
17'h128b3:	data_out=16'h9fb;
17'h128b4:	data_out=16'ha00;
17'h128b5:	data_out=16'h9ff;
17'h128b6:	data_out=16'h88fd;
17'h128b7:	data_out=16'h8c6;
17'h128b8:	data_out=16'h9fe;
17'h128b9:	data_out=16'h9f6;
17'h128ba:	data_out=16'h89fd;
17'h128bb:	data_out=16'h7ce;
17'h128bc:	data_out=16'ha00;
17'h128bd:	data_out=16'h9e7;
17'h128be:	data_out=16'h9fc;
17'h128bf:	data_out=16'h9f6;
17'h128c0:	data_out=16'h81cb;
17'h128c1:	data_out=16'h82f5;
17'h128c2:	data_out=16'h8a00;
17'h128c3:	data_out=16'h9f8;
17'h128c4:	data_out=16'ha00;
17'h128c5:	data_out=16'h861;
17'h128c6:	data_out=16'h99c;
17'h128c7:	data_out=16'h89ff;
17'h128c8:	data_out=16'h89ec;
17'h128c9:	data_out=16'h89fd;
17'h128ca:	data_out=16'h8745;
17'h128cb:	data_out=16'h8a00;
17'h128cc:	data_out=16'h8a00;
17'h128cd:	data_out=16'h8a00;
17'h128ce:	data_out=16'h850e;
17'h128cf:	data_out=16'h8a00;
17'h128d0:	data_out=16'h89d9;
17'h128d1:	data_out=16'h3ad;
17'h128d2:	data_out=16'h88b1;
17'h128d3:	data_out=16'ha00;
17'h128d4:	data_out=16'ha00;
17'h128d5:	data_out=16'h40c;
17'h128d6:	data_out=16'h939;
17'h128d7:	data_out=16'h6f2;
17'h128d8:	data_out=16'h9f7;
17'h128d9:	data_out=16'h82a4;
17'h128da:	data_out=16'h9fe;
17'h128db:	data_out=16'ha00;
17'h128dc:	data_out=16'h9fd;
17'h128dd:	data_out=16'h8986;
17'h128de:	data_out=16'ha00;
17'h128df:	data_out=16'h89c6;
17'h128e0:	data_out=16'h89d1;
17'h128e1:	data_out=16'ha00;
17'h128e2:	data_out=16'h23b;
17'h128e3:	data_out=16'h9ff;
17'h128e4:	data_out=16'ha00;
17'h128e5:	data_out=16'h9fe;
17'h128e6:	data_out=16'ha00;
17'h128e7:	data_out=16'h886b;
17'h128e8:	data_out=16'h9fc;
17'h128e9:	data_out=16'h89fb;
17'h128ea:	data_out=16'h9fd;
17'h128eb:	data_out=16'h9f3;
17'h128ec:	data_out=16'h899b;
17'h128ed:	data_out=16'h9ff;
17'h128ee:	data_out=16'h9fd;
17'h128ef:	data_out=16'h8fc;
17'h128f0:	data_out=16'h9fc;
17'h128f1:	data_out=16'h80f6;
17'h128f2:	data_out=16'h9f8;
17'h128f3:	data_out=16'ha00;
17'h128f4:	data_out=16'h83b;
17'h128f5:	data_out=16'h9de;
17'h128f6:	data_out=16'h9ff;
17'h128f7:	data_out=16'h89ff;
17'h128f8:	data_out=16'h9f9;
17'h128f9:	data_out=16'h8a00;
17'h128fa:	data_out=16'ha00;
17'h128fb:	data_out=16'h9fc;
17'h128fc:	data_out=16'h872d;
17'h128fd:	data_out=16'h9ed;
17'h128fe:	data_out=16'h8531;
17'h128ff:	data_out=16'h899e;
17'h12900:	data_out=16'h88ee;
17'h12901:	data_out=16'ha00;
17'h12902:	data_out=16'h8333;
17'h12903:	data_out=16'h89fd;
17'h12904:	data_out=16'h9e3;
17'h12905:	data_out=16'h9f3;
17'h12906:	data_out=16'h8a7;
17'h12907:	data_out=16'h8a00;
17'h12908:	data_out=16'h89ad;
17'h12909:	data_out=16'h8a00;
17'h1290a:	data_out=16'ha00;
17'h1290b:	data_out=16'h89bd;
17'h1290c:	data_out=16'h8a00;
17'h1290d:	data_out=16'h8a00;
17'h1290e:	data_out=16'h9f7;
17'h1290f:	data_out=16'h89ff;
17'h12910:	data_out=16'h89fe;
17'h12911:	data_out=16'ha00;
17'h12912:	data_out=16'h85fe;
17'h12913:	data_out=16'ha00;
17'h12914:	data_out=16'h1f6;
17'h12915:	data_out=16'h553;
17'h12916:	data_out=16'h89ec;
17'h12917:	data_out=16'h8139;
17'h12918:	data_out=16'h89ff;
17'h12919:	data_out=16'h9ff;
17'h1291a:	data_out=16'h9f1;
17'h1291b:	data_out=16'h85ca;
17'h1291c:	data_out=16'h9f1;
17'h1291d:	data_out=16'ha00;
17'h1291e:	data_out=16'h898e;
17'h1291f:	data_out=16'h467;
17'h12920:	data_out=16'h9fc;
17'h12921:	data_out=16'h9f6;
17'h12922:	data_out=16'h8a00;
17'h12923:	data_out=16'h9ed;
17'h12924:	data_out=16'h9ee;
17'h12925:	data_out=16'h89fd;
17'h12926:	data_out=16'h89ef;
17'h12927:	data_out=16'ha00;
17'h12928:	data_out=16'h9f7;
17'h12929:	data_out=16'h89d2;
17'h1292a:	data_out=16'h89ff;
17'h1292b:	data_out=16'ha00;
17'h1292c:	data_out=16'h89dd;
17'h1292d:	data_out=16'h255;
17'h1292e:	data_out=16'h88a8;
17'h1292f:	data_out=16'h6da;
17'h12930:	data_out=16'h904;
17'h12931:	data_out=16'ha00;
17'h12932:	data_out=16'ha00;
17'h12933:	data_out=16'h74a;
17'h12934:	data_out=16'ha00;
17'h12935:	data_out=16'h9da;
17'h12936:	data_out=16'h8991;
17'h12937:	data_out=16'h439;
17'h12938:	data_out=16'ha00;
17'h12939:	data_out=16'h370;
17'h1293a:	data_out=16'h89ff;
17'h1293b:	data_out=16'h782;
17'h1293c:	data_out=16'ha00;
17'h1293d:	data_out=16'h9c0;
17'h1293e:	data_out=16'h9f7;
17'h1293f:	data_out=16'h9f1;
17'h12940:	data_out=16'h9e0;
17'h12941:	data_out=16'h8a00;
17'h12942:	data_out=16'h8a00;
17'h12943:	data_out=16'h3db;
17'h12944:	data_out=16'ha00;
17'h12945:	data_out=16'h4c0;
17'h12946:	data_out=16'h9e0;
17'h12947:	data_out=16'h8a00;
17'h12948:	data_out=16'h89fd;
17'h12949:	data_out=16'h89fc;
17'h1294a:	data_out=16'h8987;
17'h1294b:	data_out=16'h8a00;
17'h1294c:	data_out=16'h8a00;
17'h1294d:	data_out=16'h8a00;
17'h1294e:	data_out=16'h89d4;
17'h1294f:	data_out=16'h8a00;
17'h12950:	data_out=16'h89fa;
17'h12951:	data_out=16'h89fe;
17'h12952:	data_out=16'h8a00;
17'h12953:	data_out=16'ha00;
17'h12954:	data_out=16'h9f5;
17'h12955:	data_out=16'h86bc;
17'h12956:	data_out=16'h7a1;
17'h12957:	data_out=16'h9a2;
17'h12958:	data_out=16'h8370;
17'h12959:	data_out=16'h9d2;
17'h1295a:	data_out=16'h9f1;
17'h1295b:	data_out=16'ha00;
17'h1295c:	data_out=16'h9f9;
17'h1295d:	data_out=16'h895b;
17'h1295e:	data_out=16'h8189;
17'h1295f:	data_out=16'h89e5;
17'h12960:	data_out=16'h89cf;
17'h12961:	data_out=16'ha00;
17'h12962:	data_out=16'h88ec;
17'h12963:	data_out=16'h9b7;
17'h12964:	data_out=16'ha00;
17'h12965:	data_out=16'h9fe;
17'h12966:	data_out=16'h9fd;
17'h12967:	data_out=16'h8997;
17'h12968:	data_out=16'h9f6;
17'h12969:	data_out=16'h8a00;
17'h1296a:	data_out=16'h9f7;
17'h1296b:	data_out=16'h9ea;
17'h1296c:	data_out=16'h899f;
17'h1296d:	data_out=16'h944;
17'h1296e:	data_out=16'h9f7;
17'h1296f:	data_out=16'h9ea;
17'h12970:	data_out=16'h9f7;
17'h12971:	data_out=16'h89f0;
17'h12972:	data_out=16'h9f1;
17'h12973:	data_out=16'ha00;
17'h12974:	data_out=16'h8dd;
17'h12975:	data_out=16'h9f3;
17'h12976:	data_out=16'h9fc;
17'h12977:	data_out=16'h8a00;
17'h12978:	data_out=16'h9ee;
17'h12979:	data_out=16'h8a00;
17'h1297a:	data_out=16'h693;
17'h1297b:	data_out=16'h9f7;
17'h1297c:	data_out=16'h89f4;
17'h1297d:	data_out=16'h9d6;
17'h1297e:	data_out=16'h1dd;
17'h1297f:	data_out=16'h89da;
17'h12980:	data_out=16'h8789;
17'h12981:	data_out=16'ha00;
17'h12982:	data_out=16'h8a00;
17'h12983:	data_out=16'h89fa;
17'h12984:	data_out=16'h9f2;
17'h12985:	data_out=16'h9e8;
17'h12986:	data_out=16'h81e;
17'h12987:	data_out=16'h8a00;
17'h12988:	data_out=16'h89b9;
17'h12989:	data_out=16'h8a00;
17'h1298a:	data_out=16'ha00;
17'h1298b:	data_out=16'h89c7;
17'h1298c:	data_out=16'h8a00;
17'h1298d:	data_out=16'h8a00;
17'h1298e:	data_out=16'h9f8;
17'h1298f:	data_out=16'h8a00;
17'h12990:	data_out=16'h89fb;
17'h12991:	data_out=16'ha00;
17'h12992:	data_out=16'h8a00;
17'h12993:	data_out=16'ha00;
17'h12994:	data_out=16'h8966;
17'h12995:	data_out=16'h239;
17'h12996:	data_out=16'h89ab;
17'h12997:	data_out=16'h8962;
17'h12998:	data_out=16'h8a00;
17'h12999:	data_out=16'h9ff;
17'h1299a:	data_out=16'h9f6;
17'h1299b:	data_out=16'h89c8;
17'h1299c:	data_out=16'h6f3;
17'h1299d:	data_out=16'ha00;
17'h1299e:	data_out=16'h89bc;
17'h1299f:	data_out=16'h875c;
17'h129a0:	data_out=16'h9f7;
17'h129a1:	data_out=16'h9f7;
17'h129a2:	data_out=16'h89fb;
17'h129a3:	data_out=16'h9fd;
17'h129a4:	data_out=16'h9fc;
17'h129a5:	data_out=16'h89fa;
17'h129a6:	data_out=16'h89cb;
17'h129a7:	data_out=16'h9ff;
17'h129a8:	data_out=16'h9f6;
17'h129a9:	data_out=16'h89e3;
17'h129aa:	data_out=16'h8994;
17'h129ab:	data_out=16'h9ea;
17'h129ac:	data_out=16'h898e;
17'h129ad:	data_out=16'h4f0;
17'h129ae:	data_out=16'h8828;
17'h129af:	data_out=16'h24;
17'h129b0:	data_out=16'h8f4;
17'h129b1:	data_out=16'ha00;
17'h129b2:	data_out=16'ha00;
17'h129b3:	data_out=16'h89e4;
17'h129b4:	data_out=16'ha00;
17'h129b5:	data_out=16'h96a;
17'h129b6:	data_out=16'h8981;
17'h129b7:	data_out=16'h19b;
17'h129b8:	data_out=16'ha00;
17'h129b9:	data_out=16'h89fd;
17'h129ba:	data_out=16'h8a00;
17'h129bb:	data_out=16'h8f3;
17'h129bc:	data_out=16'ha00;
17'h129bd:	data_out=16'h526;
17'h129be:	data_out=16'h9f6;
17'h129bf:	data_out=16'h9e5;
17'h129c0:	data_out=16'h9f5;
17'h129c1:	data_out=16'h8a00;
17'h129c2:	data_out=16'h8a00;
17'h129c3:	data_out=16'h9f1;
17'h129c4:	data_out=16'ha00;
17'h129c5:	data_out=16'h188;
17'h129c6:	data_out=16'h9f0;
17'h129c7:	data_out=16'h8a00;
17'h129c8:	data_out=16'h89fd;
17'h129c9:	data_out=16'h89f9;
17'h129ca:	data_out=16'h8998;
17'h129cb:	data_out=16'h8a00;
17'h129cc:	data_out=16'h8a00;
17'h129cd:	data_out=16'h89f9;
17'h129ce:	data_out=16'h89eb;
17'h129cf:	data_out=16'h8a00;
17'h129d0:	data_out=16'h89f6;
17'h129d1:	data_out=16'h8a00;
17'h129d2:	data_out=16'h8640;
17'h129d3:	data_out=16'h9fd;
17'h129d4:	data_out=16'h9f8;
17'h129d5:	data_out=16'h89e9;
17'h129d6:	data_out=16'h935;
17'h129d7:	data_out=16'h4fc;
17'h129d8:	data_out=16'h8a00;
17'h129d9:	data_out=16'h9f0;
17'h129da:	data_out=16'h64c;
17'h129db:	data_out=16'ha00;
17'h129dc:	data_out=16'h9f1;
17'h129dd:	data_out=16'h87be;
17'h129de:	data_out=16'h83b3;
17'h129df:	data_out=16'h89d9;
17'h129e0:	data_out=16'h89cc;
17'h129e1:	data_out=16'ha00;
17'h129e2:	data_out=16'h87d4;
17'h129e3:	data_out=16'h899f;
17'h129e4:	data_out=16'ha00;
17'h129e5:	data_out=16'ha00;
17'h129e6:	data_out=16'h9df;
17'h129e7:	data_out=16'h89b9;
17'h129e8:	data_out=16'h9f7;
17'h129e9:	data_out=16'h8a00;
17'h129ea:	data_out=16'h9f8;
17'h129eb:	data_out=16'h9e8;
17'h129ec:	data_out=16'h87d7;
17'h129ed:	data_out=16'h89a7;
17'h129ee:	data_out=16'h9f8;
17'h129ef:	data_out=16'ha00;
17'h129f0:	data_out=16'h9f8;
17'h129f1:	data_out=16'h89cc;
17'h129f2:	data_out=16'ha00;
17'h129f3:	data_out=16'ha00;
17'h129f4:	data_out=16'h8cf;
17'h129f5:	data_out=16'h9e7;
17'h129f6:	data_out=16'h9f2;
17'h129f7:	data_out=16'h8a00;
17'h129f8:	data_out=16'h9d4;
17'h129f9:	data_out=16'h8a00;
17'h129fa:	data_out=16'h896e;
17'h129fb:	data_out=16'h9f6;
17'h129fc:	data_out=16'h8a00;
17'h129fd:	data_out=16'h8933;
17'h129fe:	data_out=16'h85b;
17'h129ff:	data_out=16'h89f9;
17'h12a00:	data_out=16'h943;
17'h12a01:	data_out=16'ha00;
17'h12a02:	data_out=16'h89c2;
17'h12a03:	data_out=16'h89e7;
17'h12a04:	data_out=16'h9f6;
17'h12a05:	data_out=16'h9e3;
17'h12a06:	data_out=16'h50f;
17'h12a07:	data_out=16'h8a00;
17'h12a08:	data_out=16'h8998;
17'h12a09:	data_out=16'h8a00;
17'h12a0a:	data_out=16'ha00;
17'h12a0b:	data_out=16'h89c2;
17'h12a0c:	data_out=16'h8a00;
17'h12a0d:	data_out=16'h8a00;
17'h12a0e:	data_out=16'h9fe;
17'h12a0f:	data_out=16'h89e0;
17'h12a10:	data_out=16'h89f5;
17'h12a11:	data_out=16'ha00;
17'h12a12:	data_out=16'h8a00;
17'h12a13:	data_out=16'ha00;
17'h12a14:	data_out=16'h89fc;
17'h12a15:	data_out=16'h287;
17'h12a16:	data_out=16'h897e;
17'h12a17:	data_out=16'h89ef;
17'h12a18:	data_out=16'h8a00;
17'h12a19:	data_out=16'h9f7;
17'h12a1a:	data_out=16'h9f0;
17'h12a1b:	data_out=16'h89e0;
17'h12a1c:	data_out=16'h354;
17'h12a1d:	data_out=16'ha00;
17'h12a1e:	data_out=16'h89e2;
17'h12a1f:	data_out=16'h89e0;
17'h12a20:	data_out=16'h9f0;
17'h12a21:	data_out=16'h9fd;
17'h12a22:	data_out=16'h89e1;
17'h12a23:	data_out=16'ha00;
17'h12a24:	data_out=16'ha00;
17'h12a25:	data_out=16'h89e1;
17'h12a26:	data_out=16'h896b;
17'h12a27:	data_out=16'h9fc;
17'h12a28:	data_out=16'h9fc;
17'h12a29:	data_out=16'h89f0;
17'h12a2a:	data_out=16'h8931;
17'h12a2b:	data_out=16'h9e3;
17'h12a2c:	data_out=16'h8987;
17'h12a2d:	data_out=16'h897e;
17'h12a2e:	data_out=16'h88f7;
17'h12a2f:	data_out=16'h7bf;
17'h12a30:	data_out=16'h7a9;
17'h12a31:	data_out=16'ha00;
17'h12a32:	data_out=16'ha00;
17'h12a33:	data_out=16'h8a00;
17'h12a34:	data_out=16'ha00;
17'h12a35:	data_out=16'h825;
17'h12a36:	data_out=16'h88d5;
17'h12a37:	data_out=16'h899c;
17'h12a38:	data_out=16'ha00;
17'h12a39:	data_out=16'h8a00;
17'h12a3a:	data_out=16'h89fd;
17'h12a3b:	data_out=16'h73c;
17'h12a3c:	data_out=16'ha00;
17'h12a3d:	data_out=16'h390;
17'h12a3e:	data_out=16'h9fc;
17'h12a3f:	data_out=16'h9e2;
17'h12a40:	data_out=16'ha00;
17'h12a41:	data_out=16'h89f3;
17'h12a42:	data_out=16'h89dc;
17'h12a43:	data_out=16'h53e;
17'h12a44:	data_out=16'h9f9;
17'h12a45:	data_out=16'h1ef;
17'h12a46:	data_out=16'h9f1;
17'h12a47:	data_out=16'h8a00;
17'h12a48:	data_out=16'h89fa;
17'h12a49:	data_out=16'h89d5;
17'h12a4a:	data_out=16'h8944;
17'h12a4b:	data_out=16'h8a00;
17'h12a4c:	data_out=16'h89ef;
17'h12a4d:	data_out=16'h89dc;
17'h12a4e:	data_out=16'h8562;
17'h12a4f:	data_out=16'h89f4;
17'h12a50:	data_out=16'h89f8;
17'h12a51:	data_out=16'h8a00;
17'h12a52:	data_out=16'h848b;
17'h12a53:	data_out=16'h9f5;
17'h12a54:	data_out=16'h9ff;
17'h12a55:	data_out=16'h8a00;
17'h12a56:	data_out=16'h881d;
17'h12a57:	data_out=16'h896a;
17'h12a58:	data_out=16'h8a00;
17'h12a59:	data_out=16'h9f2;
17'h12a5a:	data_out=16'h82d8;
17'h12a5b:	data_out=16'ha00;
17'h12a5c:	data_out=16'h9eb;
17'h12a5d:	data_out=16'h444;
17'h12a5e:	data_out=16'h96c;
17'h12a5f:	data_out=16'h89d9;
17'h12a60:	data_out=16'h899a;
17'h12a61:	data_out=16'ha00;
17'h12a62:	data_out=16'h87fa;
17'h12a63:	data_out=16'h8a00;
17'h12a64:	data_out=16'ha00;
17'h12a65:	data_out=16'ha00;
17'h12a66:	data_out=16'h895c;
17'h12a67:	data_out=16'h89e8;
17'h12a68:	data_out=16'h9fd;
17'h12a69:	data_out=16'h8a00;
17'h12a6a:	data_out=16'h9fe;
17'h12a6b:	data_out=16'h881;
17'h12a6c:	data_out=16'ha00;
17'h12a6d:	data_out=16'h8a00;
17'h12a6e:	data_out=16'h9fe;
17'h12a6f:	data_out=16'ha00;
17'h12a70:	data_out=16'h9fe;
17'h12a71:	data_out=16'h89df;
17'h12a72:	data_out=16'ha00;
17'h12a73:	data_out=16'ha00;
17'h12a74:	data_out=16'h7d7;
17'h12a75:	data_out=16'h9e1;
17'h12a76:	data_out=16'h846a;
17'h12a77:	data_out=16'h8a00;
17'h12a78:	data_out=16'h9d2;
17'h12a79:	data_out=16'h8a00;
17'h12a7a:	data_out=16'h89fe;
17'h12a7b:	data_out=16'h9fc;
17'h12a7c:	data_out=16'h8a00;
17'h12a7d:	data_out=16'h89fe;
17'h12a7e:	data_out=16'h47d;
17'h12a7f:	data_out=16'h89fa;
17'h12a80:	data_out=16'h9f6;
17'h12a81:	data_out=16'ha00;
17'h12a82:	data_out=16'h89a2;
17'h12a83:	data_out=16'h8961;
17'h12a84:	data_out=16'h9f7;
17'h12a85:	data_out=16'h9cb;
17'h12a86:	data_out=16'h81c5;
17'h12a87:	data_out=16'h8a00;
17'h12a88:	data_out=16'h896a;
17'h12a89:	data_out=16'h89b3;
17'h12a8a:	data_out=16'ha00;
17'h12a8b:	data_out=16'h8864;
17'h12a8c:	data_out=16'h89de;
17'h12a8d:	data_out=16'h8a00;
17'h12a8e:	data_out=16'h856f;
17'h12a8f:	data_out=16'h89ac;
17'h12a90:	data_out=16'h893f;
17'h12a91:	data_out=16'ha00;
17'h12a92:	data_out=16'h8a00;
17'h12a93:	data_out=16'ha00;
17'h12a94:	data_out=16'h89b0;
17'h12a95:	data_out=16'h7a4;
17'h12a96:	data_out=16'h81d6;
17'h12a97:	data_out=16'h89a0;
17'h12a98:	data_out=16'h8a00;
17'h12a99:	data_out=16'h9f5;
17'h12a9a:	data_out=16'h9e4;
17'h12a9b:	data_out=16'h8975;
17'h12a9c:	data_out=16'h24;
17'h12a9d:	data_out=16'ha00;
17'h12a9e:	data_out=16'h89a9;
17'h12a9f:	data_out=16'h89ef;
17'h12aa0:	data_out=16'h9f0;
17'h12aa1:	data_out=16'h874b;
17'h12aa2:	data_out=16'h897d;
17'h12aa3:	data_out=16'ha00;
17'h12aa4:	data_out=16'ha00;
17'h12aa5:	data_out=16'h8969;
17'h12aa6:	data_out=16'h890f;
17'h12aa7:	data_out=16'h9fc;
17'h12aa8:	data_out=16'h8941;
17'h12aa9:	data_out=16'h89e7;
17'h12aaa:	data_out=16'h878c;
17'h12aab:	data_out=16'h9e8;
17'h12aac:	data_out=16'h8059;
17'h12aad:	data_out=16'h897c;
17'h12aae:	data_out=16'h87ea;
17'h12aaf:	data_out=16'h9fe;
17'h12ab0:	data_out=16'h604;
17'h12ab1:	data_out=16'ha00;
17'h12ab2:	data_out=16'ha00;
17'h12ab3:	data_out=16'h89fc;
17'h12ab4:	data_out=16'ha00;
17'h12ab5:	data_out=16'h9ff;
17'h12ab6:	data_out=16'h867d;
17'h12ab7:	data_out=16'h897d;
17'h12ab8:	data_out=16'ha00;
17'h12ab9:	data_out=16'h89fd;
17'h12aba:	data_out=16'h89e8;
17'h12abb:	data_out=16'h945;
17'h12abc:	data_out=16'ha00;
17'h12abd:	data_out=16'h9e0;
17'h12abe:	data_out=16'h8947;
17'h12abf:	data_out=16'h9ca;
17'h12ac0:	data_out=16'ha00;
17'h12ac1:	data_out=16'h89b4;
17'h12ac2:	data_out=16'h897c;
17'h12ac3:	data_out=16'h510;
17'h12ac4:	data_out=16'h9e2;
17'h12ac5:	data_out=16'h758;
17'h12ac6:	data_out=16'h9f2;
17'h12ac7:	data_out=16'h89fd;
17'h12ac8:	data_out=16'h887f;
17'h12ac9:	data_out=16'h88a1;
17'h12aca:	data_out=16'hee;
17'h12acb:	data_out=16'h89af;
17'h12acc:	data_out=16'h89d0;
17'h12acd:	data_out=16'h8985;
17'h12ace:	data_out=16'h81c3;
17'h12acf:	data_out=16'h89c4;
17'h12ad0:	data_out=16'h890b;
17'h12ad1:	data_out=16'h8a00;
17'h12ad2:	data_out=16'h24b;
17'h12ad3:	data_out=16'h9f9;
17'h12ad4:	data_out=16'h9fc;
17'h12ad5:	data_out=16'h89c4;
17'h12ad6:	data_out=16'h86c0;
17'h12ad7:	data_out=16'h897b;
17'h12ad8:	data_out=16'h89ff;
17'h12ad9:	data_out=16'ha00;
17'h12ada:	data_out=16'h89fe;
17'h12adb:	data_out=16'ha00;
17'h12adc:	data_out=16'h9e8;
17'h12add:	data_out=16'ha00;
17'h12ade:	data_out=16'ha00;
17'h12adf:	data_out=16'h89ce;
17'h12ae0:	data_out=16'h8921;
17'h12ae1:	data_out=16'ha00;
17'h12ae2:	data_out=16'h85f3;
17'h12ae3:	data_out=16'h89e0;
17'h12ae4:	data_out=16'ha00;
17'h12ae5:	data_out=16'ha00;
17'h12ae6:	data_out=16'h8766;
17'h12ae7:	data_out=16'h89d9;
17'h12ae8:	data_out=16'h884e;
17'h12ae9:	data_out=16'h89d3;
17'h12aea:	data_out=16'h84a7;
17'h12aeb:	data_out=16'ha00;
17'h12aec:	data_out=16'h9ff;
17'h12aed:	data_out=16'h89e1;
17'h12aee:	data_out=16'h84a8;
17'h12aef:	data_out=16'ha00;
17'h12af0:	data_out=16'h8504;
17'h12af1:	data_out=16'h89d2;
17'h12af2:	data_out=16'ha00;
17'h12af3:	data_out=16'ha00;
17'h12af4:	data_out=16'h632;
17'h12af5:	data_out=16'h9db;
17'h12af6:	data_out=16'h8735;
17'h12af7:	data_out=16'h89b0;
17'h12af8:	data_out=16'ha00;
17'h12af9:	data_out=16'h8a00;
17'h12afa:	data_out=16'h89b8;
17'h12afb:	data_out=16'h894c;
17'h12afc:	data_out=16'h8a00;
17'h12afd:	data_out=16'h89f5;
17'h12afe:	data_out=16'h18d;
17'h12aff:	data_out=16'h89fa;
17'h12b00:	data_out=16'h9d9;
17'h12b01:	data_out=16'ha00;
17'h12b02:	data_out=16'h898c;
17'h12b03:	data_out=16'h87fc;
17'h12b04:	data_out=16'ha00;
17'h12b05:	data_out=16'h9e8;
17'h12b06:	data_out=16'h89c5;
17'h12b07:	data_out=16'h89f0;
17'h12b08:	data_out=16'h8933;
17'h12b09:	data_out=16'h8993;
17'h12b0a:	data_out=16'ha00;
17'h12b0b:	data_out=16'h87c7;
17'h12b0c:	data_out=16'h80c4;
17'h12b0d:	data_out=16'h8a00;
17'h12b0e:	data_out=16'h89e5;
17'h12b0f:	data_out=16'h89a5;
17'h12b10:	data_out=16'h8619;
17'h12b11:	data_out=16'ha00;
17'h12b12:	data_out=16'h8a00;
17'h12b13:	data_out=16'h890;
17'h12b14:	data_out=16'h898e;
17'h12b15:	data_out=16'h5dd;
17'h12b16:	data_out=16'h9f1;
17'h12b17:	data_out=16'h8964;
17'h12b18:	data_out=16'h8a00;
17'h12b19:	data_out=16'h761;
17'h12b1a:	data_out=16'ha00;
17'h12b1b:	data_out=16'h8923;
17'h12b1c:	data_out=16'h8964;
17'h12b1d:	data_out=16'ha00;
17'h12b1e:	data_out=16'h8989;
17'h12b1f:	data_out=16'h89e8;
17'h12b20:	data_out=16'h9fc;
17'h12b21:	data_out=16'h89e8;
17'h12b22:	data_out=16'h897a;
17'h12b23:	data_out=16'h839;
17'h12b24:	data_out=16'h80f;
17'h12b25:	data_out=16'h8949;
17'h12b26:	data_out=16'h88f7;
17'h12b27:	data_out=16'ha00;
17'h12b28:	data_out=16'h89e8;
17'h12b29:	data_out=16'h89eb;
17'h12b2a:	data_out=16'h859c;
17'h12b2b:	data_out=16'h81c;
17'h12b2c:	data_out=16'h9ea;
17'h12b2d:	data_out=16'h89e2;
17'h12b2e:	data_out=16'h8848;
17'h12b2f:	data_out=16'ha00;
17'h12b30:	data_out=16'h3da;
17'h12b31:	data_out=16'ha00;
17'h12b32:	data_out=16'ha00;
17'h12b33:	data_out=16'h89f5;
17'h12b34:	data_out=16'ha00;
17'h12b35:	data_out=16'ha00;
17'h12b36:	data_out=16'h857a;
17'h12b37:	data_out=16'h8977;
17'h12b38:	data_out=16'h9fe;
17'h12b39:	data_out=16'h89fb;
17'h12b3a:	data_out=16'h89d2;
17'h12b3b:	data_out=16'h9d2;
17'h12b3c:	data_out=16'h800a;
17'h12b3d:	data_out=16'h9d5;
17'h12b3e:	data_out=16'h89e7;
17'h12b3f:	data_out=16'h9e7;
17'h12b40:	data_out=16'ha00;
17'h12b41:	data_out=16'h88d2;
17'h12b42:	data_out=16'h920;
17'h12b43:	data_out=16'h1e1;
17'h12b44:	data_out=16'ha00;
17'h12b45:	data_out=16'h7e0;
17'h12b46:	data_out=16'h8586;
17'h12b47:	data_out=16'h89ff;
17'h12b48:	data_out=16'h8650;
17'h12b49:	data_out=16'h889a;
17'h12b4a:	data_out=16'h9f3;
17'h12b4b:	data_out=16'h8e6;
17'h12b4c:	data_out=16'h89f3;
17'h12b4d:	data_out=16'h897f;
17'h12b4e:	data_out=16'h85a8;
17'h12b4f:	data_out=16'h89d0;
17'h12b50:	data_out=16'h8364;
17'h12b51:	data_out=16'h8a00;
17'h12b52:	data_out=16'h8247;
17'h12b53:	data_out=16'h9fa;
17'h12b54:	data_out=16'h9fc;
17'h12b55:	data_out=16'h8997;
17'h12b56:	data_out=16'h88db;
17'h12b57:	data_out=16'h89b4;
17'h12b58:	data_out=16'h89ed;
17'h12b59:	data_out=16'ha00;
17'h12b5a:	data_out=16'h89ff;
17'h12b5b:	data_out=16'ha00;
17'h12b5c:	data_out=16'h4c2;
17'h12b5d:	data_out=16'ha00;
17'h12b5e:	data_out=16'ha00;
17'h12b5f:	data_out=16'h89b4;
17'h12b60:	data_out=16'h88b4;
17'h12b61:	data_out=16'ha00;
17'h12b62:	data_out=16'h86da;
17'h12b63:	data_out=16'h89d1;
17'h12b64:	data_out=16'h9f2;
17'h12b65:	data_out=16'ha00;
17'h12b66:	data_out=16'h8564;
17'h12b67:	data_out=16'h89ff;
17'h12b68:	data_out=16'h89e9;
17'h12b69:	data_out=16'h89ce;
17'h12b6a:	data_out=16'h89e2;
17'h12b6b:	data_out=16'ha00;
17'h12b6c:	data_out=16'h9f0;
17'h12b6d:	data_out=16'h89d4;
17'h12b6e:	data_out=16'h89e2;
17'h12b6f:	data_out=16'ha00;
17'h12b70:	data_out=16'h89e4;
17'h12b71:	data_out=16'h89dd;
17'h12b72:	data_out=16'ha00;
17'h12b73:	data_out=16'ha00;
17'h12b74:	data_out=16'h40f;
17'h12b75:	data_out=16'h8154;
17'h12b76:	data_out=16'h8986;
17'h12b77:	data_out=16'h8954;
17'h12b78:	data_out=16'ha00;
17'h12b79:	data_out=16'h89e7;
17'h12b7a:	data_out=16'h8997;
17'h12b7b:	data_out=16'h89e7;
17'h12b7c:	data_out=16'h8a00;
17'h12b7d:	data_out=16'h89ec;
17'h12b7e:	data_out=16'h89b2;
17'h12b7f:	data_out=16'h89f5;
17'h12b80:	data_out=16'h9ea;
17'h12b81:	data_out=16'ha00;
17'h12b82:	data_out=16'h8960;
17'h12b83:	data_out=16'h893b;
17'h12b84:	data_out=16'ha00;
17'h12b85:	data_out=16'h9ff;
17'h12b86:	data_out=16'h89bf;
17'h12b87:	data_out=16'ha00;
17'h12b88:	data_out=16'h86f7;
17'h12b89:	data_out=16'h88db;
17'h12b8a:	data_out=16'ha00;
17'h12b8b:	data_out=16'h8957;
17'h12b8c:	data_out=16'ha00;
17'h12b8d:	data_out=16'h8a00;
17'h12b8e:	data_out=16'h89ed;
17'h12b8f:	data_out=16'h8954;
17'h12b90:	data_out=16'h831a;
17'h12b91:	data_out=16'ha00;
17'h12b92:	data_out=16'h8a00;
17'h12b93:	data_out=16'h85ee;
17'h12b94:	data_out=16'h89c8;
17'h12b95:	data_out=16'h80d4;
17'h12b96:	data_out=16'ha00;
17'h12b97:	data_out=16'h89a0;
17'h12b98:	data_out=16'h8a00;
17'h12b99:	data_out=16'h8924;
17'h12b9a:	data_out=16'ha00;
17'h12b9b:	data_out=16'h8950;
17'h12b9c:	data_out=16'h89d1;
17'h12b9d:	data_out=16'ha00;
17'h12b9e:	data_out=16'h8986;
17'h12b9f:	data_out=16'h89e8;
17'h12ba0:	data_out=16'h9ff;
17'h12ba1:	data_out=16'h89ee;
17'h12ba2:	data_out=16'h897f;
17'h12ba3:	data_out=16'h506;
17'h12ba4:	data_out=16'h4fc;
17'h12ba5:	data_out=16'h88bc;
17'h12ba6:	data_out=16'h88da;
17'h12ba7:	data_out=16'ha00;
17'h12ba8:	data_out=16'h89ed;
17'h12ba9:	data_out=16'h89b1;
17'h12baa:	data_out=16'h808f;
17'h12bab:	data_out=16'h81fc;
17'h12bac:	data_out=16'ha00;
17'h12bad:	data_out=16'h89e7;
17'h12bae:	data_out=16'h88d2;
17'h12baf:	data_out=16'ha00;
17'h12bb0:	data_out=16'h42f;
17'h12bb1:	data_out=16'ha00;
17'h12bb2:	data_out=16'ha00;
17'h12bb3:	data_out=16'h89fe;
17'h12bb4:	data_out=16'ha00;
17'h12bb5:	data_out=16'ha00;
17'h12bb6:	data_out=16'h8288;
17'h12bb7:	data_out=16'h895f;
17'h12bb8:	data_out=16'h9f7;
17'h12bb9:	data_out=16'h89ff;
17'h12bba:	data_out=16'h8706;
17'h12bbb:	data_out=16'h9fd;
17'h12bbc:	data_out=16'h8861;
17'h12bbd:	data_out=16'h9f9;
17'h12bbe:	data_out=16'h89ec;
17'h12bbf:	data_out=16'h9ff;
17'h12bc0:	data_out=16'ha00;
17'h12bc1:	data_out=16'h852e;
17'h12bc2:	data_out=16'h9fb;
17'h12bc3:	data_out=16'h88c6;
17'h12bc4:	data_out=16'ha00;
17'h12bc5:	data_out=16'h12d;
17'h12bc6:	data_out=16'h8681;
17'h12bc7:	data_out=16'h89f1;
17'h12bc8:	data_out=16'h17e;
17'h12bc9:	data_out=16'h86a7;
17'h12bca:	data_out=16'ha00;
17'h12bcb:	data_out=16'h9e8;
17'h12bcc:	data_out=16'h89f6;
17'h12bcd:	data_out=16'h889d;
17'h12bce:	data_out=16'h8374;
17'h12bcf:	data_out=16'h223;
17'h12bd0:	data_out=16'h8350;
17'h12bd1:	data_out=16'h8a00;
17'h12bd2:	data_out=16'h3ad;
17'h12bd3:	data_out=16'h9fb;
17'h12bd4:	data_out=16'h9fc;
17'h12bd5:	data_out=16'h89a4;
17'h12bd6:	data_out=16'h887e;
17'h12bd7:	data_out=16'h89b6;
17'h12bd8:	data_out=16'h89fb;
17'h12bd9:	data_out=16'ha00;
17'h12bda:	data_out=16'h8a00;
17'h12bdb:	data_out=16'h48e;
17'h12bdc:	data_out=16'h8976;
17'h12bdd:	data_out=16'ha00;
17'h12bde:	data_out=16'ha00;
17'h12bdf:	data_out=16'h862f;
17'h12be0:	data_out=16'h887d;
17'h12be1:	data_out=16'ha00;
17'h12be2:	data_out=16'h8924;
17'h12be3:	data_out=16'h89e4;
17'h12be4:	data_out=16'h9e6;
17'h12be5:	data_out=16'ha00;
17'h12be6:	data_out=16'h88ba;
17'h12be7:	data_out=16'h8a00;
17'h12be8:	data_out=16'h89ee;
17'h12be9:	data_out=16'h89c8;
17'h12bea:	data_out=16'h89ec;
17'h12beb:	data_out=16'ha00;
17'h12bec:	data_out=16'ha00;
17'h12bed:	data_out=16'h89e7;
17'h12bee:	data_out=16'h89ec;
17'h12bef:	data_out=16'ha00;
17'h12bf0:	data_out=16'h89ec;
17'h12bf1:	data_out=16'h8978;
17'h12bf2:	data_out=16'ha00;
17'h12bf3:	data_out=16'h9ff;
17'h12bf4:	data_out=16'h434;
17'h12bf5:	data_out=16'h88c1;
17'h12bf6:	data_out=16'h89b8;
17'h12bf7:	data_out=16'h8661;
17'h12bf8:	data_out=16'ha00;
17'h12bf9:	data_out=16'h896e;
17'h12bfa:	data_out=16'h89ba;
17'h12bfb:	data_out=16'h89ec;
17'h12bfc:	data_out=16'h8a00;
17'h12bfd:	data_out=16'h89d2;
17'h12bfe:	data_out=16'h89be;
17'h12bff:	data_out=16'h89ec;
17'h12c00:	data_out=16'h9aa;
17'h12c01:	data_out=16'h9ff;
17'h12c02:	data_out=16'h8996;
17'h12c03:	data_out=16'h89ca;
17'h12c04:	data_out=16'h9fc;
17'h12c05:	data_out=16'h9fe;
17'h12c06:	data_out=16'h89d0;
17'h12c07:	data_out=16'ha00;
17'h12c08:	data_out=16'h85fe;
17'h12c09:	data_out=16'h86ed;
17'h12c0a:	data_out=16'ha00;
17'h12c0b:	data_out=16'h89b2;
17'h12c0c:	data_out=16'ha00;
17'h12c0d:	data_out=16'h8a00;
17'h12c0e:	data_out=16'h89f1;
17'h12c0f:	data_out=16'h884a;
17'h12c10:	data_out=16'h81cb;
17'h12c11:	data_out=16'ha00;
17'h12c12:	data_out=16'h8a00;
17'h12c13:	data_out=16'h8740;
17'h12c14:	data_out=16'h89f7;
17'h12c15:	data_out=16'h86a4;
17'h12c16:	data_out=16'h9f4;
17'h12c17:	data_out=16'h89e0;
17'h12c18:	data_out=16'h8a00;
17'h12c19:	data_out=16'h8487;
17'h12c1a:	data_out=16'h9fb;
17'h12c1b:	data_out=16'h89c8;
17'h12c1c:	data_out=16'h8a00;
17'h12c1d:	data_out=16'ha00;
17'h12c1e:	data_out=16'h89de;
17'h12c1f:	data_out=16'h89f1;
17'h12c20:	data_out=16'h9de;
17'h12c21:	data_out=16'h89f2;
17'h12c22:	data_out=16'h88b0;
17'h12c23:	data_out=16'h6f2;
17'h12c24:	data_out=16'h70a;
17'h12c25:	data_out=16'h8745;
17'h12c26:	data_out=16'h897a;
17'h12c27:	data_out=16'h9fd;
17'h12c28:	data_out=16'h89ef;
17'h12c29:	data_out=16'h895f;
17'h12c2a:	data_out=16'h9ea;
17'h12c2b:	data_out=16'h88eb;
17'h12c2c:	data_out=16'h9f2;
17'h12c2d:	data_out=16'h89f9;
17'h12c2e:	data_out=16'h8972;
17'h12c2f:	data_out=16'h9ff;
17'h12c30:	data_out=16'h9ec;
17'h12c31:	data_out=16'ha00;
17'h12c32:	data_out=16'ha00;
17'h12c33:	data_out=16'h8a00;
17'h12c34:	data_out=16'ha00;
17'h12c35:	data_out=16'h9fc;
17'h12c36:	data_out=16'h81a2;
17'h12c37:	data_out=16'h8997;
17'h12c38:	data_out=16'h9dd;
17'h12c39:	data_out=16'h8a00;
17'h12c3a:	data_out=16'h85a1;
17'h12c3b:	data_out=16'h9f9;
17'h12c3c:	data_out=16'h8977;
17'h12c3d:	data_out=16'h8720;
17'h12c3e:	data_out=16'h89ee;
17'h12c3f:	data_out=16'h9fe;
17'h12c40:	data_out=16'ha00;
17'h12c41:	data_out=16'h9ec;
17'h12c42:	data_out=16'h9f9;
17'h12c43:	data_out=16'h853c;
17'h12c44:	data_out=16'h88d;
17'h12c45:	data_out=16'h85fa;
17'h12c46:	data_out=16'h3fd;
17'h12c47:	data_out=16'h89db;
17'h12c48:	data_out=16'h5bf;
17'h12c49:	data_out=16'h286;
17'h12c4a:	data_out=16'ha00;
17'h12c4b:	data_out=16'h9f4;
17'h12c4c:	data_out=16'h8250;
17'h12c4d:	data_out=16'h861e;
17'h12c4e:	data_out=16'hcc;
17'h12c4f:	data_out=16'h9c8;
17'h12c50:	data_out=16'h855e;
17'h12c51:	data_out=16'h8a00;
17'h12c52:	data_out=16'h9b4;
17'h12c53:	data_out=16'h9fc;
17'h12c54:	data_out=16'h9f4;
17'h12c55:	data_out=16'h89e3;
17'h12c56:	data_out=16'h88f1;
17'h12c57:	data_out=16'h89f3;
17'h12c58:	data_out=16'h8a00;
17'h12c59:	data_out=16'ha00;
17'h12c5a:	data_out=16'h8a00;
17'h12c5b:	data_out=16'h85c1;
17'h12c5c:	data_out=16'h89e3;
17'h12c5d:	data_out=16'ha00;
17'h12c5e:	data_out=16'ha00;
17'h12c5f:	data_out=16'h86b0;
17'h12c60:	data_out=16'h8926;
17'h12c61:	data_out=16'h9fe;
17'h12c62:	data_out=16'h899a;
17'h12c63:	data_out=16'h89f1;
17'h12c64:	data_out=16'h9bf;
17'h12c65:	data_out=16'ha00;
17'h12c66:	data_out=16'h9e6;
17'h12c67:	data_out=16'h89fb;
17'h12c68:	data_out=16'h89f2;
17'h12c69:	data_out=16'h89f4;
17'h12c6a:	data_out=16'h89f2;
17'h12c6b:	data_out=16'ha00;
17'h12c6c:	data_out=16'h9d9;
17'h12c6d:	data_out=16'h89f4;
17'h12c6e:	data_out=16'h89f2;
17'h12c6f:	data_out=16'ha00;
17'h12c70:	data_out=16'h89f1;
17'h12c71:	data_out=16'h8922;
17'h12c72:	data_out=16'ha00;
17'h12c73:	data_out=16'h9fb;
17'h12c74:	data_out=16'h9e5;
17'h12c75:	data_out=16'h88e9;
17'h12c76:	data_out=16'h89ac;
17'h12c77:	data_out=16'h8297;
17'h12c78:	data_out=16'ha00;
17'h12c79:	data_out=16'h8331;
17'h12c7a:	data_out=16'h89e6;
17'h12c7b:	data_out=16'h89ee;
17'h12c7c:	data_out=16'h8a00;
17'h12c7d:	data_out=16'h89d0;
17'h12c7e:	data_out=16'h89f8;
17'h12c7f:	data_out=16'h89ff;
17'h12c80:	data_out=16'h89a7;
17'h12c81:	data_out=16'h9d5;
17'h12c82:	data_out=16'h89cb;
17'h12c83:	data_out=16'h89ff;
17'h12c84:	data_out=16'h9e6;
17'h12c85:	data_out=16'h9df;
17'h12c86:	data_out=16'h89f4;
17'h12c87:	data_out=16'h9ff;
17'h12c88:	data_out=16'h892b;
17'h12c89:	data_out=16'h87d6;
17'h12c8a:	data_out=16'h9d1;
17'h12c8b:	data_out=16'h89e5;
17'h12c8c:	data_out=16'ha00;
17'h12c8d:	data_out=16'h8a00;
17'h12c8e:	data_out=16'h88e2;
17'h12c8f:	data_out=16'h89aa;
17'h12c90:	data_out=16'h8329;
17'h12c91:	data_out=16'ha00;
17'h12c92:	data_out=16'h8a00;
17'h12c93:	data_out=16'h8877;
17'h12c94:	data_out=16'h89ff;
17'h12c95:	data_out=16'h88fd;
17'h12c96:	data_out=16'h8117;
17'h12c97:	data_out=16'h89ff;
17'h12c98:	data_out=16'h8a00;
17'h12c99:	data_out=16'ha00;
17'h12c9a:	data_out=16'h9d1;
17'h12c9b:	data_out=16'h89ff;
17'h12c9c:	data_out=16'h8a00;
17'h12c9d:	data_out=16'h9e8;
17'h12c9e:	data_out=16'h89f8;
17'h12c9f:	data_out=16'h89f4;
17'h12ca0:	data_out=16'h89e9;
17'h12ca1:	data_out=16'h8885;
17'h12ca2:	data_out=16'h88c1;
17'h12ca3:	data_out=16'h8530;
17'h12ca4:	data_out=16'h84c3;
17'h12ca5:	data_out=16'h8764;
17'h12ca6:	data_out=16'h89d4;
17'h12ca7:	data_out=16'h89d1;
17'h12ca8:	data_out=16'h8750;
17'h12ca9:	data_out=16'h8080;
17'h12caa:	data_out=16'h1bd;
17'h12cab:	data_out=16'h8953;
17'h12cac:	data_out=16'h8674;
17'h12cad:	data_out=16'h89ff;
17'h12cae:	data_out=16'h89f0;
17'h12caf:	data_out=16'h9bf;
17'h12cb0:	data_out=16'ha00;
17'h12cb1:	data_out=16'h87a6;
17'h12cb2:	data_out=16'ha00;
17'h12cb3:	data_out=16'h8a00;
17'h12cb4:	data_out=16'h9e1;
17'h12cb5:	data_out=16'h70c;
17'h12cb6:	data_out=16'h8620;
17'h12cb7:	data_out=16'h89ca;
17'h12cb8:	data_out=16'h88b2;
17'h12cb9:	data_out=16'h8a00;
17'h12cba:	data_out=16'h8661;
17'h12cbb:	data_out=16'h9e8;
17'h12cbc:	data_out=16'h89ff;
17'h12cbd:	data_out=16'h89ef;
17'h12cbe:	data_out=16'h873d;
17'h12cbf:	data_out=16'h9dd;
17'h12cc0:	data_out=16'ha00;
17'h12cc1:	data_out=16'h4a1;
17'h12cc2:	data_out=16'h9dd;
17'h12cc3:	data_out=16'h9fe;
17'h12cc4:	data_out=16'h89d9;
17'h12cc5:	data_out=16'h888e;
17'h12cc6:	data_out=16'h9eb;
17'h12cc7:	data_out=16'h89f2;
17'h12cc8:	data_out=16'h8452;
17'h12cc9:	data_out=16'h83e0;
17'h12cca:	data_out=16'h9fe;
17'h12ccb:	data_out=16'h9e4;
17'h12ccc:	data_out=16'h3a7;
17'h12ccd:	data_out=16'h8775;
17'h12cce:	data_out=16'h8281;
17'h12ccf:	data_out=16'h9dc;
17'h12cd0:	data_out=16'h8857;
17'h12cd1:	data_out=16'h8a00;
17'h12cd2:	data_out=16'h9e0;
17'h12cd3:	data_out=16'h2ae;
17'h12cd4:	data_out=16'h8946;
17'h12cd5:	data_out=16'h89c7;
17'h12cd6:	data_out=16'h89a3;
17'h12cd7:	data_out=16'h89fb;
17'h12cd8:	data_out=16'h8a00;
17'h12cd9:	data_out=16'h9d0;
17'h12cda:	data_out=16'h8a00;
17'h12cdb:	data_out=16'h89ba;
17'h12cdc:	data_out=16'h89f6;
17'h12cdd:	data_out=16'h9fc;
17'h12cde:	data_out=16'ha00;
17'h12cdf:	data_out=16'h89da;
17'h12ce0:	data_out=16'h89e0;
17'h12ce1:	data_out=16'h9cb;
17'h12ce2:	data_out=16'h89f1;
17'h12ce3:	data_out=16'h89fe;
17'h12ce4:	data_out=16'h721;
17'h12ce5:	data_out=16'ha00;
17'h12ce6:	data_out=16'h9fb;
17'h12ce7:	data_out=16'h89f7;
17'h12ce8:	data_out=16'h8852;
17'h12ce9:	data_out=16'h8a00;
17'h12cea:	data_out=16'h8960;
17'h12ceb:	data_out=16'h9fe;
17'h12cec:	data_out=16'h677;
17'h12ced:	data_out=16'h89fe;
17'h12cee:	data_out=16'h8959;
17'h12cef:	data_out=16'ha00;
17'h12cf0:	data_out=16'h8906;
17'h12cf1:	data_out=16'h89f0;
17'h12cf2:	data_out=16'h9d2;
17'h12cf3:	data_out=16'h9cb;
17'h12cf4:	data_out=16'ha00;
17'h12cf5:	data_out=16'h8618;
17'h12cf6:	data_out=16'h8997;
17'h12cf7:	data_out=16'h8342;
17'h12cf8:	data_out=16'ha00;
17'h12cf9:	data_out=16'h89ad;
17'h12cfa:	data_out=16'h89fc;
17'h12cfb:	data_out=16'h872f;
17'h12cfc:	data_out=16'h8a00;
17'h12cfd:	data_out=16'h89d7;
17'h12cfe:	data_out=16'h89fc;
17'h12cff:	data_out=16'h8a00;
17'h12d00:	data_out=16'h89e7;
17'h12d01:	data_out=16'h4b8;
17'h12d02:	data_out=16'h899a;
17'h12d03:	data_out=16'h89eb;
17'h12d04:	data_out=16'h6b4;
17'h12d05:	data_out=16'h9ce;
17'h12d06:	data_out=16'h89fe;
17'h12d07:	data_out=16'ha00;
17'h12d08:	data_out=16'h8971;
17'h12d09:	data_out=16'h8878;
17'h12d0a:	data_out=16'h75b;
17'h12d0b:	data_out=16'h89e3;
17'h12d0c:	data_out=16'h9ff;
17'h12d0d:	data_out=16'h89d1;
17'h12d0e:	data_out=16'h8aa;
17'h12d0f:	data_out=16'h81f2;
17'h12d10:	data_out=16'h89aa;
17'h12d11:	data_out=16'h8a00;
17'h12d12:	data_out=16'h89fc;
17'h12d13:	data_out=16'h87bd;
17'h12d14:	data_out=16'h89e5;
17'h12d15:	data_out=16'h84b8;
17'h12d16:	data_out=16'h9e6;
17'h12d17:	data_out=16'h89be;
17'h12d18:	data_out=16'h89fa;
17'h12d19:	data_out=16'h9bf;
17'h12d1a:	data_out=16'h956;
17'h12d1b:	data_out=16'h89f7;
17'h12d1c:	data_out=16'h8a00;
17'h12d1d:	data_out=16'h89f7;
17'h12d1e:	data_out=16'h89f3;
17'h12d1f:	data_out=16'h898b;
17'h12d20:	data_out=16'h89f5;
17'h12d21:	data_out=16'h8e2;
17'h12d22:	data_out=16'h89fb;
17'h12d23:	data_out=16'h89da;
17'h12d24:	data_out=16'h89da;
17'h12d25:	data_out=16'h8923;
17'h12d26:	data_out=16'h89fd;
17'h12d27:	data_out=16'h89fa;
17'h12d28:	data_out=16'h95d;
17'h12d29:	data_out=16'h9ec;
17'h12d2a:	data_out=16'h3b5;
17'h12d2b:	data_out=16'h89b7;
17'h12d2c:	data_out=16'h9d9;
17'h12d2d:	data_out=16'h89ff;
17'h12d2e:	data_out=16'h89e7;
17'h12d2f:	data_out=16'h435;
17'h12d30:	data_out=16'ha00;
17'h12d31:	data_out=16'h89fe;
17'h12d32:	data_out=16'h9aa;
17'h12d33:	data_out=16'h89f6;
17'h12d34:	data_out=16'h8032;
17'h12d35:	data_out=16'h8017;
17'h12d36:	data_out=16'h863b;
17'h12d37:	data_out=16'h89bf;
17'h12d38:	data_out=16'h8a00;
17'h12d39:	data_out=16'h89f7;
17'h12d3a:	data_out=16'h87af;
17'h12d3b:	data_out=16'h381;
17'h12d3c:	data_out=16'h8a00;
17'h12d3d:	data_out=16'h89f8;
17'h12d3e:	data_out=16'h962;
17'h12d3f:	data_out=16'h9cd;
17'h12d40:	data_out=16'h9cd;
17'h12d41:	data_out=16'hf8;
17'h12d42:	data_out=16'h9a8;
17'h12d43:	data_out=16'ha00;
17'h12d44:	data_out=16'h8a00;
17'h12d45:	data_out=16'h83e7;
17'h12d46:	data_out=16'h872c;
17'h12d47:	data_out=16'h89e3;
17'h12d48:	data_out=16'h88c9;
17'h12d49:	data_out=16'h87cc;
17'h12d4a:	data_out=16'h9fc;
17'h12d4b:	data_out=16'h986;
17'h12d4c:	data_out=16'h89f3;
17'h12d4d:	data_out=16'h89f7;
17'h12d4e:	data_out=16'h314;
17'h12d4f:	data_out=16'h86eb;
17'h12d50:	data_out=16'h860e;
17'h12d51:	data_out=16'h89ad;
17'h12d52:	data_out=16'h87c8;
17'h12d53:	data_out=16'h82c9;
17'h12d54:	data_out=16'h89f0;
17'h12d55:	data_out=16'h85e9;
17'h12d56:	data_out=16'h89fe;
17'h12d57:	data_out=16'h89fd;
17'h12d58:	data_out=16'h89f9;
17'h12d59:	data_out=16'h877;
17'h12d5a:	data_out=16'h89e8;
17'h12d5b:	data_out=16'h8a00;
17'h12d5c:	data_out=16'h89e7;
17'h12d5d:	data_out=16'h9ca;
17'h12d5e:	data_out=16'ha00;
17'h12d5f:	data_out=16'h89fc;
17'h12d60:	data_out=16'h89fe;
17'h12d61:	data_out=16'h8ea;
17'h12d62:	data_out=16'h87e0;
17'h12d63:	data_out=16'h89f4;
17'h12d64:	data_out=16'h89f4;
17'h12d65:	data_out=16'h95d;
17'h12d66:	data_out=16'h9ef;
17'h12d67:	data_out=16'h89f2;
17'h12d68:	data_out=16'h90d;
17'h12d69:	data_out=16'h89f7;
17'h12d6a:	data_out=16'h86e;
17'h12d6b:	data_out=16'h9db;
17'h12d6c:	data_out=16'h83e4;
17'h12d6d:	data_out=16'h89f4;
17'h12d6e:	data_out=16'h871;
17'h12d6f:	data_out=16'h9f7;
17'h12d70:	data_out=16'h897;
17'h12d71:	data_out=16'h8561;
17'h12d72:	data_out=16'h960;
17'h12d73:	data_out=16'h9a2;
17'h12d74:	data_out=16'ha00;
17'h12d75:	data_out=16'h5af;
17'h12d76:	data_out=16'h89f5;
17'h12d77:	data_out=16'h860a;
17'h12d78:	data_out=16'h9fb;
17'h12d79:	data_out=16'h89ed;
17'h12d7a:	data_out=16'h89f0;
17'h12d7b:	data_out=16'h966;
17'h12d7c:	data_out=16'h89f6;
17'h12d7d:	data_out=16'h8971;
17'h12d7e:	data_out=16'h89fa;
17'h12d7f:	data_out=16'h8a00;
17'h12d80:	data_out=16'h8732;
17'h12d81:	data_out=16'h8676;
17'h12d82:	data_out=16'h88ab;
17'h12d83:	data_out=16'h8950;
17'h12d84:	data_out=16'h634;
17'h12d85:	data_out=16'h9ca;
17'h12d86:	data_out=16'h8a00;
17'h12d87:	data_out=16'ha00;
17'h12d88:	data_out=16'h887f;
17'h12d89:	data_out=16'h8996;
17'h12d8a:	data_out=16'h1b9;
17'h12d8b:	data_out=16'h89d6;
17'h12d8c:	data_out=16'h9ff;
17'h12d8d:	data_out=16'h8160;
17'h12d8e:	data_out=16'h8e8;
17'h12d8f:	data_out=16'h17;
17'h12d90:	data_out=16'h89ed;
17'h12d91:	data_out=16'h8a00;
17'h12d92:	data_out=16'h89b9;
17'h12d93:	data_out=16'h89b3;
17'h12d94:	data_out=16'h89bd;
17'h12d95:	data_out=16'h4f0;
17'h12d96:	data_out=16'h9f1;
17'h12d97:	data_out=16'h87d9;
17'h12d98:	data_out=16'h89ed;
17'h12d99:	data_out=16'h992;
17'h12d9a:	data_out=16'h984;
17'h12d9b:	data_out=16'h850d;
17'h12d9c:	data_out=16'h89fd;
17'h12d9d:	data_out=16'h89fe;
17'h12d9e:	data_out=16'h8848;
17'h12d9f:	data_out=16'h88b2;
17'h12da0:	data_out=16'h89e3;
17'h12da1:	data_out=16'h90c;
17'h12da2:	data_out=16'h8a00;
17'h12da3:	data_out=16'h89ef;
17'h12da4:	data_out=16'h89f0;
17'h12da5:	data_out=16'h89df;
17'h12da6:	data_out=16'h89f2;
17'h12da7:	data_out=16'h89f0;
17'h12da8:	data_out=16'h95f;
17'h12da9:	data_out=16'h9f1;
17'h12daa:	data_out=16'h1c7;
17'h12dab:	data_out=16'h89ab;
17'h12dac:	data_out=16'h9f0;
17'h12dad:	data_out=16'h89ff;
17'h12dae:	data_out=16'h899b;
17'h12daf:	data_out=16'h8340;
17'h12db0:	data_out=16'ha00;
17'h12db1:	data_out=16'h4bb;
17'h12db2:	data_out=16'h5f3;
17'h12db3:	data_out=16'h89eb;
17'h12db4:	data_out=16'h82c4;
17'h12db5:	data_out=16'hab;
17'h12db6:	data_out=16'h856c;
17'h12db7:	data_out=16'h89af;
17'h12db8:	data_out=16'h8a00;
17'h12db9:	data_out=16'h89f9;
17'h12dba:	data_out=16'h87ea;
17'h12dbb:	data_out=16'h1b0;
17'h12dbc:	data_out=16'h8a00;
17'h12dbd:	data_out=16'h89f4;
17'h12dbe:	data_out=16'h965;
17'h12dbf:	data_out=16'h9ca;
17'h12dc0:	data_out=16'h97d;
17'h12dc1:	data_out=16'h9d7;
17'h12dc2:	data_out=16'h4c;
17'h12dc3:	data_out=16'ha00;
17'h12dc4:	data_out=16'h38f;
17'h12dc5:	data_out=16'h69c;
17'h12dc6:	data_out=16'h8a00;
17'h12dc7:	data_out=16'h89bf;
17'h12dc8:	data_out=16'h89b0;
17'h12dc9:	data_out=16'h89e1;
17'h12dca:	data_out=16'h9fe;
17'h12dcb:	data_out=16'h875;
17'h12dcc:	data_out=16'h89ff;
17'h12dcd:	data_out=16'h8a00;
17'h12dce:	data_out=16'h38d;
17'h12dcf:	data_out=16'h88a7;
17'h12dd0:	data_out=16'h85b4;
17'h12dd1:	data_out=16'h80cd;
17'h12dd2:	data_out=16'h8653;
17'h12dd3:	data_out=16'h8477;
17'h12dd4:	data_out=16'h89d8;
17'h12dd5:	data_out=16'h8037;
17'h12dd6:	data_out=16'h89ff;
17'h12dd7:	data_out=16'h8a00;
17'h12dd8:	data_out=16'h85cf;
17'h12dd9:	data_out=16'h82e7;
17'h12dda:	data_out=16'h8873;
17'h12ddb:	data_out=16'h89fd;
17'h12ddc:	data_out=16'h86a4;
17'h12ddd:	data_out=16'h9e1;
17'h12dde:	data_out=16'h38a;
17'h12ddf:	data_out=16'h89ef;
17'h12de0:	data_out=16'h89ff;
17'h12de1:	data_out=16'h5d3;
17'h12de2:	data_out=16'h87c1;
17'h12de3:	data_out=16'h89d6;
17'h12de4:	data_out=16'h89f7;
17'h12de5:	data_out=16'h2f0;
17'h12de6:	data_out=16'ha00;
17'h12de7:	data_out=16'h9e8;
17'h12de8:	data_out=16'h927;
17'h12de9:	data_out=16'h89eb;
17'h12dea:	data_out=16'h8be;
17'h12deb:	data_out=16'h9d4;
17'h12dec:	data_out=16'h57f;
17'h12ded:	data_out=16'h89db;
17'h12dee:	data_out=16'h8c0;
17'h12def:	data_out=16'h9ee;
17'h12df0:	data_out=16'h8dc;
17'h12df1:	data_out=16'h576;
17'h12df2:	data_out=16'h80c4;
17'h12df3:	data_out=16'h86b;
17'h12df4:	data_out=16'ha00;
17'h12df5:	data_out=16'h7c3;
17'h12df6:	data_out=16'h89f3;
17'h12df7:	data_out=16'h89a2;
17'h12df8:	data_out=16'h9a9;
17'h12df9:	data_out=16'h856a;
17'h12dfa:	data_out=16'h89c6;
17'h12dfb:	data_out=16'h968;
17'h12dfc:	data_out=16'h89ed;
17'h12dfd:	data_out=16'h83b0;
17'h12dfe:	data_out=16'h88a4;
17'h12dff:	data_out=16'h8a00;
17'h12e00:	data_out=16'h8453;
17'h12e01:	data_out=16'h86d5;
17'h12e02:	data_out=16'h89ca;
17'h12e03:	data_out=16'h8920;
17'h12e04:	data_out=16'h9d4;
17'h12e05:	data_out=16'h9ef;
17'h12e06:	data_out=16'h8a00;
17'h12e07:	data_out=16'h9ff;
17'h12e08:	data_out=16'h8978;
17'h12e09:	data_out=16'h89af;
17'h12e0a:	data_out=16'h80f6;
17'h12e0b:	data_out=16'h89e4;
17'h12e0c:	data_out=16'h9fb;
17'h12e0d:	data_out=16'h822d;
17'h12e0e:	data_out=16'h623;
17'h12e0f:	data_out=16'h8995;
17'h12e10:	data_out=16'h89ea;
17'h12e11:	data_out=16'h8a00;
17'h12e12:	data_out=16'h89dc;
17'h12e13:	data_out=16'h89c8;
17'h12e14:	data_out=16'h899c;
17'h12e15:	data_out=16'h602;
17'h12e16:	data_out=16'h9f6;
17'h12e17:	data_out=16'h8771;
17'h12e18:	data_out=16'h89f5;
17'h12e19:	data_out=16'h9e5;
17'h12e1a:	data_out=16'h9e8;
17'h12e1b:	data_out=16'h899f;
17'h12e1c:	data_out=16'h89af;
17'h12e1d:	data_out=16'h89ca;
17'h12e1e:	data_out=16'h8982;
17'h12e1f:	data_out=16'h89a0;
17'h12e20:	data_out=16'h8962;
17'h12e21:	data_out=16'h663;
17'h12e22:	data_out=16'h8a00;
17'h12e23:	data_out=16'h89fd;
17'h12e24:	data_out=16'h89fc;
17'h12e25:	data_out=16'h8a00;
17'h12e26:	data_out=16'h8a00;
17'h12e27:	data_out=16'h3e1;
17'h12e28:	data_out=16'h6ee;
17'h12e29:	data_out=16'h9f5;
17'h12e2a:	data_out=16'h889b;
17'h12e2b:	data_out=16'h89bc;
17'h12e2c:	data_out=16'h9f8;
17'h12e2d:	data_out=16'h8a00;
17'h12e2e:	data_out=16'h89c5;
17'h12e2f:	data_out=16'h831e;
17'h12e30:	data_out=16'ha00;
17'h12e31:	data_out=16'h9de;
17'h12e32:	data_out=16'h613;
17'h12e33:	data_out=16'h89c7;
17'h12e34:	data_out=16'h8791;
17'h12e35:	data_out=16'hd4;
17'h12e36:	data_out=16'h8919;
17'h12e37:	data_out=16'h89ca;
17'h12e38:	data_out=16'h8a00;
17'h12e39:	data_out=16'h89e3;
17'h12e3a:	data_out=16'h89d6;
17'h12e3b:	data_out=16'h858;
17'h12e3c:	data_out=16'h89e3;
17'h12e3d:	data_out=16'h8970;
17'h12e3e:	data_out=16'h6ff;
17'h12e3f:	data_out=16'h9ef;
17'h12e40:	data_out=16'h9d3;
17'h12e41:	data_out=16'h9df;
17'h12e42:	data_out=16'h89be;
17'h12e43:	data_out=16'ha00;
17'h12e44:	data_out=16'h9d8;
17'h12e45:	data_out=16'h76e;
17'h12e46:	data_out=16'h8a00;
17'h12e47:	data_out=16'h89ff;
17'h12e48:	data_out=16'h89b9;
17'h12e49:	data_out=16'h89f4;
17'h12e4a:	data_out=16'ha00;
17'h12e4b:	data_out=16'h89a6;
17'h12e4c:	data_out=16'h8a00;
17'h12e4d:	data_out=16'h8a00;
17'h12e4e:	data_out=16'h8341;
17'h12e4f:	data_out=16'h8a00;
17'h12e50:	data_out=16'h2b5;
17'h12e51:	data_out=16'h8132;
17'h12e52:	data_out=16'h89f8;
17'h12e53:	data_out=16'h88b1;
17'h12e54:	data_out=16'h899b;
17'h12e55:	data_out=16'h8679;
17'h12e56:	data_out=16'h8a00;
17'h12e57:	data_out=16'h8a00;
17'h12e58:	data_out=16'h8718;
17'h12e59:	data_out=16'h89c3;
17'h12e5a:	data_out=16'h8905;
17'h12e5b:	data_out=16'h235;
17'h12e5c:	data_out=16'h82c3;
17'h12e5d:	data_out=16'h2ce;
17'h12e5e:	data_out=16'h1ec;
17'h12e5f:	data_out=16'h89f0;
17'h12e60:	data_out=16'h8a00;
17'h12e61:	data_out=16'h7be;
17'h12e62:	data_out=16'h8956;
17'h12e63:	data_out=16'h89aa;
17'h12e64:	data_out=16'h89fe;
17'h12e65:	data_out=16'h2a0;
17'h12e66:	data_out=16'ha00;
17'h12e67:	data_out=16'ha00;
17'h12e68:	data_out=16'h66d;
17'h12e69:	data_out=16'h89fa;
17'h12e6a:	data_out=16'h5e5;
17'h12e6b:	data_out=16'h9eb;
17'h12e6c:	data_out=16'h426;
17'h12e6d:	data_out=16'h89b1;
17'h12e6e:	data_out=16'h5ea;
17'h12e6f:	data_out=16'ha00;
17'h12e70:	data_out=16'h617;
17'h12e71:	data_out=16'h87d1;
17'h12e72:	data_out=16'h8949;
17'h12e73:	data_out=16'h8273;
17'h12e74:	data_out=16'ha00;
17'h12e75:	data_out=16'h936;
17'h12e76:	data_out=16'h89e8;
17'h12e77:	data_out=16'h89ab;
17'h12e78:	data_out=16'h442;
17'h12e79:	data_out=16'h89f2;
17'h12e7a:	data_out=16'h8998;
17'h12e7b:	data_out=16'h70a;
17'h12e7c:	data_out=16'h89f4;
17'h12e7d:	data_out=16'h80aa;
17'h12e7e:	data_out=16'h89f0;
17'h12e7f:	data_out=16'h88a0;
17'h12e80:	data_out=16'h874f;
17'h12e81:	data_out=16'h85b8;
17'h12e82:	data_out=16'h89c8;
17'h12e83:	data_out=16'h8969;
17'h12e84:	data_out=16'h9f8;
17'h12e85:	data_out=16'ha00;
17'h12e86:	data_out=16'h89f6;
17'h12e87:	data_out=16'h9ed;
17'h12e88:	data_out=16'h89c5;
17'h12e89:	data_out=16'h89e4;
17'h12e8a:	data_out=16'h874;
17'h12e8b:	data_out=16'h89f9;
17'h12e8c:	data_out=16'h654;
17'h12e8d:	data_out=16'h87ec;
17'h12e8e:	data_out=16'h967;
17'h12e8f:	data_out=16'h89b6;
17'h12e90:	data_out=16'h89d7;
17'h12e91:	data_out=16'h8a00;
17'h12e92:	data_out=16'h89f7;
17'h12e93:	data_out=16'h89cb;
17'h12e94:	data_out=16'h89ad;
17'h12e95:	data_out=16'h9f8;
17'h12e96:	data_out=16'h9fb;
17'h12e97:	data_out=16'h8969;
17'h12e98:	data_out=16'h89e5;
17'h12e99:	data_out=16'ha00;
17'h12e9a:	data_out=16'ha00;
17'h12e9b:	data_out=16'h89a4;
17'h12e9c:	data_out=16'h8984;
17'h12e9d:	data_out=16'h89cc;
17'h12e9e:	data_out=16'h89a3;
17'h12e9f:	data_out=16'h89cb;
17'h12ea0:	data_out=16'h86de;
17'h12ea1:	data_out=16'h984;
17'h12ea2:	data_out=16'h89fe;
17'h12ea3:	data_out=16'h8073;
17'h12ea4:	data_out=16'h8066;
17'h12ea5:	data_out=16'h89ff;
17'h12ea6:	data_out=16'h89fd;
17'h12ea7:	data_out=16'h89d0;
17'h12ea8:	data_out=16'h9a7;
17'h12ea9:	data_out=16'h9f9;
17'h12eaa:	data_out=16'h88fd;
17'h12eab:	data_out=16'h89dd;
17'h12eac:	data_out=16'h9fe;
17'h12ead:	data_out=16'h8a00;
17'h12eae:	data_out=16'h89f5;
17'h12eaf:	data_out=16'h8214;
17'h12eb0:	data_out=16'ha00;
17'h12eb1:	data_out=16'h9f6;
17'h12eb2:	data_out=16'h9f5;
17'h12eb3:	data_out=16'h89db;
17'h12eb4:	data_out=16'h8917;
17'h12eb5:	data_out=16'h8b7;
17'h12eb6:	data_out=16'h892a;
17'h12eb7:	data_out=16'h89d6;
17'h12eb8:	data_out=16'h8a00;
17'h12eb9:	data_out=16'h89ed;
17'h12eba:	data_out=16'h89e4;
17'h12ebb:	data_out=16'h9fc;
17'h12ebc:	data_out=16'h8962;
17'h12ebd:	data_out=16'h8379;
17'h12ebe:	data_out=16'h9b1;
17'h12ebf:	data_out=16'ha00;
17'h12ec0:	data_out=16'h9fd;
17'h12ec1:	data_out=16'h87d3;
17'h12ec2:	data_out=16'h89d6;
17'h12ec3:	data_out=16'h9fc;
17'h12ec4:	data_out=16'h9ed;
17'h12ec5:	data_out=16'h9f8;
17'h12ec6:	data_out=16'h89f4;
17'h12ec7:	data_out=16'h8a00;
17'h12ec8:	data_out=16'h89f1;
17'h12ec9:	data_out=16'h8928;
17'h12eca:	data_out=16'ha00;
17'h12ecb:	data_out=16'h89cf;
17'h12ecc:	data_out=16'h89ff;
17'h12ecd:	data_out=16'h89f3;
17'h12ece:	data_out=16'h89f6;
17'h12ecf:	data_out=16'h89ff;
17'h12ed0:	data_out=16'h9fd;
17'h12ed1:	data_out=16'h547;
17'h12ed2:	data_out=16'h5aa;
17'h12ed3:	data_out=16'h88ba;
17'h12ed4:	data_out=16'h8921;
17'h12ed5:	data_out=16'h88a2;
17'h12ed6:	data_out=16'h89fa;
17'h12ed7:	data_out=16'h89fe;
17'h12ed8:	data_out=16'h87a8;
17'h12ed9:	data_out=16'h9b9;
17'h12eda:	data_out=16'h89ba;
17'h12edb:	data_out=16'h9cf;
17'h12edc:	data_out=16'h324;
17'h12edd:	data_out=16'h5bb;
17'h12ede:	data_out=16'h18c;
17'h12edf:	data_out=16'h89e4;
17'h12ee0:	data_out=16'h89e7;
17'h12ee1:	data_out=16'h9f8;
17'h12ee2:	data_out=16'h898b;
17'h12ee3:	data_out=16'h89cf;
17'h12ee4:	data_out=16'h8a00;
17'h12ee5:	data_out=16'h9f3;
17'h12ee6:	data_out=16'ha00;
17'h12ee7:	data_out=16'ha00;
17'h12ee8:	data_out=16'h96c;
17'h12ee9:	data_out=16'h89fc;
17'h12eea:	data_out=16'h953;
17'h12eeb:	data_out=16'ha00;
17'h12eec:	data_out=16'h32b;
17'h12eed:	data_out=16'h89d3;
17'h12eee:	data_out=16'h957;
17'h12eef:	data_out=16'ha00;
17'h12ef0:	data_out=16'h968;
17'h12ef1:	data_out=16'h865d;
17'h12ef2:	data_out=16'h37b;
17'h12ef3:	data_out=16'h9fe;
17'h12ef4:	data_out=16'ha00;
17'h12ef5:	data_out=16'h9fe;
17'h12ef6:	data_out=16'h8224;
17'h12ef7:	data_out=16'h89d6;
17'h12ef8:	data_out=16'h216;
17'h12ef9:	data_out=16'h89e8;
17'h12efa:	data_out=16'h89b0;
17'h12efb:	data_out=16'h9b9;
17'h12efc:	data_out=16'h899b;
17'h12efd:	data_out=16'h930;
17'h12efe:	data_out=16'h89e6;
17'h12eff:	data_out=16'h86a;
17'h12f00:	data_out=16'h8960;
17'h12f01:	data_out=16'h89cc;
17'h12f02:	data_out=16'h89e2;
17'h12f03:	data_out=16'h896f;
17'h12f04:	data_out=16'ha00;
17'h12f05:	data_out=16'ha00;
17'h12f06:	data_out=16'h89ca;
17'h12f07:	data_out=16'h89a4;
17'h12f08:	data_out=16'h89ea;
17'h12f09:	data_out=16'h89ba;
17'h12f0a:	data_out=16'h856;
17'h12f0b:	data_out=16'h89dc;
17'h12f0c:	data_out=16'h89e6;
17'h12f0d:	data_out=16'h88be;
17'h12f0e:	data_out=16'h2b3;
17'h12f0f:	data_out=16'h89ce;
17'h12f10:	data_out=16'h89c3;
17'h12f11:	data_out=16'h8a00;
17'h12f12:	data_out=16'h89f4;
17'h12f13:	data_out=16'h89a4;
17'h12f14:	data_out=16'h8979;
17'h12f15:	data_out=16'ha00;
17'h12f16:	data_out=16'h9fe;
17'h12f17:	data_out=16'h8940;
17'h12f18:	data_out=16'h89d6;
17'h12f19:	data_out=16'ha00;
17'h12f1a:	data_out=16'ha00;
17'h12f1b:	data_out=16'h89a9;
17'h12f1c:	data_out=16'h892e;
17'h12f1d:	data_out=16'h89fb;
17'h12f1e:	data_out=16'h897d;
17'h12f1f:	data_out=16'h8904;
17'h12f20:	data_out=16'h8728;
17'h12f21:	data_out=16'h27a;
17'h12f22:	data_out=16'h89ed;
17'h12f23:	data_out=16'h8392;
17'h12f24:	data_out=16'h838c;
17'h12f25:	data_out=16'h89e5;
17'h12f26:	data_out=16'h8a00;
17'h12f27:	data_out=16'h89da;
17'h12f28:	data_out=16'h21b;
17'h12f29:	data_out=16'h9f7;
17'h12f2a:	data_out=16'h89c7;
17'h12f2b:	data_out=16'h408;
17'h12f2c:	data_out=16'h9ff;
17'h12f2d:	data_out=16'h8a00;
17'h12f2e:	data_out=16'h89da;
17'h12f2f:	data_out=16'h86c9;
17'h12f30:	data_out=16'ha00;
17'h12f31:	data_out=16'h9f9;
17'h12f32:	data_out=16'h9d5;
17'h12f33:	data_out=16'h899b;
17'h12f34:	data_out=16'h89da;
17'h12f35:	data_out=16'h950;
17'h12f36:	data_out=16'h89cd;
17'h12f37:	data_out=16'h89f2;
17'h12f38:	data_out=16'h8a00;
17'h12f39:	data_out=16'h89ad;
17'h12f3a:	data_out=16'h89db;
17'h12f3b:	data_out=16'h9e6;
17'h12f3c:	data_out=16'h8892;
17'h12f3d:	data_out=16'h85ef;
17'h12f3e:	data_out=16'h21b;
17'h12f3f:	data_out=16'ha00;
17'h12f40:	data_out=16'ha00;
17'h12f41:	data_out=16'h895c;
17'h12f42:	data_out=16'h8a00;
17'h12f43:	data_out=16'h9e1;
17'h12f44:	data_out=16'h9fe;
17'h12f45:	data_out=16'h9ff;
17'h12f46:	data_out=16'h8a00;
17'h12f47:	data_out=16'h8a00;
17'h12f48:	data_out=16'h89d8;
17'h12f49:	data_out=16'h8969;
17'h12f4a:	data_out=16'h8567;
17'h12f4b:	data_out=16'h89fe;
17'h12f4c:	data_out=16'h8a00;
17'h12f4d:	data_out=16'h89b7;
17'h12f4e:	data_out=16'h8a00;
17'h12f4f:	data_out=16'h8a00;
17'h12f50:	data_out=16'h9ff;
17'h12f51:	data_out=16'h9d3;
17'h12f52:	data_out=16'h8a;
17'h12f53:	data_out=16'h89a3;
17'h12f54:	data_out=16'h8982;
17'h12f55:	data_out=16'h896b;
17'h12f56:	data_out=16'h89fe;
17'h12f57:	data_out=16'h89b2;
17'h12f58:	data_out=16'h813c;
17'h12f59:	data_out=16'h87d9;
17'h12f5a:	data_out=16'h89ac;
17'h12f5b:	data_out=16'h9df;
17'h12f5c:	data_out=16'h37;
17'h12f5d:	data_out=16'h82f8;
17'h12f5e:	data_out=16'h85d4;
17'h12f5f:	data_out=16'h89f3;
17'h12f60:	data_out=16'h8a00;
17'h12f61:	data_out=16'ha00;
17'h12f62:	data_out=16'h89ab;
17'h12f63:	data_out=16'h8996;
17'h12f64:	data_out=16'h8a00;
17'h12f65:	data_out=16'h807d;
17'h12f66:	data_out=16'ha00;
17'h12f67:	data_out=16'ha00;
17'h12f68:	data_out=16'h24b;
17'h12f69:	data_out=16'h8a00;
17'h12f6a:	data_out=16'h2f8;
17'h12f6b:	data_out=16'h9ff;
17'h12f6c:	data_out=16'h83c8;
17'h12f6d:	data_out=16'h8999;
17'h12f6e:	data_out=16'h2f9;
17'h12f6f:	data_out=16'ha00;
17'h12f70:	data_out=16'h2d3;
17'h12f71:	data_out=16'h8928;
17'h12f72:	data_out=16'h8840;
17'h12f73:	data_out=16'h9fd;
17'h12f74:	data_out=16'ha00;
17'h12f75:	data_out=16'ha00;
17'h12f76:	data_out=16'ha00;
17'h12f77:	data_out=16'h89d2;
17'h12f78:	data_out=16'h272;
17'h12f79:	data_out=16'h89f9;
17'h12f7a:	data_out=16'h898a;
17'h12f7b:	data_out=16'h21d;
17'h12f7c:	data_out=16'h89cc;
17'h12f7d:	data_out=16'h8ea;
17'h12f7e:	data_out=16'h89e8;
17'h12f7f:	data_out=16'h9f3;
17'h12f80:	data_out=16'h89ac;
17'h12f81:	data_out=16'h89dd;
17'h12f82:	data_out=16'h89f0;
17'h12f83:	data_out=16'h89b0;
17'h12f84:	data_out=16'ha00;
17'h12f85:	data_out=16'ha00;
17'h12f86:	data_out=16'h89e3;
17'h12f87:	data_out=16'h89fa;
17'h12f88:	data_out=16'h89f4;
17'h12f89:	data_out=16'h89e9;
17'h12f8a:	data_out=16'h9b8;
17'h12f8b:	data_out=16'h89e2;
17'h12f8c:	data_out=16'h8a00;
17'h12f8d:	data_out=16'h89c0;
17'h12f8e:	data_out=16'h9fe;
17'h12f8f:	data_out=16'h89f0;
17'h12f90:	data_out=16'h89d9;
17'h12f91:	data_out=16'h89f3;
17'h12f92:	data_out=16'h89f6;
17'h12f93:	data_out=16'h89c5;
17'h12f94:	data_out=16'h897b;
17'h12f95:	data_out=16'ha00;
17'h12f96:	data_out=16'h854c;
17'h12f97:	data_out=16'h8993;
17'h12f98:	data_out=16'h89db;
17'h12f99:	data_out=16'h9fb;
17'h12f9a:	data_out=16'ha00;
17'h12f9b:	data_out=16'h89c2;
17'h12f9c:	data_out=16'h89ae;
17'h12f9d:	data_out=16'h89f9;
17'h12f9e:	data_out=16'h8983;
17'h12f9f:	data_out=16'h8795;
17'h12fa0:	data_out=16'h867a;
17'h12fa1:	data_out=16'h989;
17'h12fa2:	data_out=16'h89a2;
17'h12fa3:	data_out=16'h36d;
17'h12fa4:	data_out=16'h382;
17'h12fa5:	data_out=16'h89c7;
17'h12fa6:	data_out=16'h8a00;
17'h12fa7:	data_out=16'h8929;
17'h12fa8:	data_out=16'h8b6;
17'h12fa9:	data_out=16'h9f3;
17'h12faa:	data_out=16'h89f5;
17'h12fab:	data_out=16'h9ff;
17'h12fac:	data_out=16'h539;
17'h12fad:	data_out=16'h8a00;
17'h12fae:	data_out=16'h89e1;
17'h12faf:	data_out=16'h8923;
17'h12fb0:	data_out=16'ha00;
17'h12fb1:	data_out=16'h9fb;
17'h12fb2:	data_out=16'h9bd;
17'h12fb3:	data_out=16'h89a7;
17'h12fb4:	data_out=16'h8a00;
17'h12fb5:	data_out=16'h9fb;
17'h12fb6:	data_out=16'h89ee;
17'h12fb7:	data_out=16'h89f0;
17'h12fb8:	data_out=16'h89fb;
17'h12fb9:	data_out=16'h89b3;
17'h12fba:	data_out=16'h89c2;
17'h12fbb:	data_out=16'h9eb;
17'h12fbc:	data_out=16'h86e9;
17'h12fbd:	data_out=16'h859f;
17'h12fbe:	data_out=16'h8af;
17'h12fbf:	data_out=16'ha00;
17'h12fc0:	data_out=16'h2c8;
17'h12fc1:	data_out=16'h88ff;
17'h12fc2:	data_out=16'h8a00;
17'h12fc3:	data_out=16'ha00;
17'h12fc4:	data_out=16'ha00;
17'h12fc5:	data_out=16'ha00;
17'h12fc6:	data_out=16'h89f2;
17'h12fc7:	data_out=16'h89fd;
17'h12fc8:	data_out=16'h89f4;
17'h12fc9:	data_out=16'h86a1;
17'h12fca:	data_out=16'h88c6;
17'h12fcb:	data_out=16'h8a00;
17'h12fcc:	data_out=16'h8a00;
17'h12fcd:	data_out=16'h88f2;
17'h12fce:	data_out=16'h8a00;
17'h12fcf:	data_out=16'h8a00;
17'h12fd0:	data_out=16'h7dc;
17'h12fd1:	data_out=16'h8b7;
17'h12fd2:	data_out=16'h89e;
17'h12fd3:	data_out=16'h88a1;
17'h12fd4:	data_out=16'h8982;
17'h12fd5:	data_out=16'h898f;
17'h12fd6:	data_out=16'h78c;
17'h12fd7:	data_out=16'h8608;
17'h12fd8:	data_out=16'h8157;
17'h12fd9:	data_out=16'h462;
17'h12fda:	data_out=16'h89c0;
17'h12fdb:	data_out=16'ha00;
17'h12fdc:	data_out=16'h8459;
17'h12fdd:	data_out=16'h87ef;
17'h12fde:	data_out=16'h896d;
17'h12fdf:	data_out=16'h89f6;
17'h12fe0:	data_out=16'h8a00;
17'h12fe1:	data_out=16'ha00;
17'h12fe2:	data_out=16'h89d5;
17'h12fe3:	data_out=16'h899c;
17'h12fe4:	data_out=16'h8a00;
17'h12fe5:	data_out=16'h8260;
17'h12fe6:	data_out=16'ha00;
17'h12fe7:	data_out=16'ha00;
17'h12fe8:	data_out=16'h93b;
17'h12fe9:	data_out=16'h89ff;
17'h12fea:	data_out=16'h9fe;
17'h12feb:	data_out=16'h83e;
17'h12fec:	data_out=16'h88af;
17'h12fed:	data_out=16'h89a2;
17'h12fee:	data_out=16'h9fe;
17'h12fef:	data_out=16'ha00;
17'h12ff0:	data_out=16'h9fe;
17'h12ff1:	data_out=16'h8996;
17'h12ff2:	data_out=16'h80f1;
17'h12ff3:	data_out=16'h9ff;
17'h12ff4:	data_out=16'h9e5;
17'h12ff5:	data_out=16'ha00;
17'h12ff6:	data_out=16'ha00;
17'h12ff7:	data_out=16'h89f4;
17'h12ff8:	data_out=16'h918;
17'h12ff9:	data_out=16'h89f9;
17'h12ffa:	data_out=16'h898c;
17'h12ffb:	data_out=16'h8ab;
17'h12ffc:	data_out=16'h89d5;
17'h12ffd:	data_out=16'h745;
17'h12ffe:	data_out=16'h8a00;
17'h12fff:	data_out=16'ha00;
17'h13000:	data_out=16'h868a;
17'h13001:	data_out=16'h8991;
17'h13002:	data_out=16'h89dc;
17'h13003:	data_out=16'h89a4;
17'h13004:	data_out=16'ha00;
17'h13005:	data_out=16'ha00;
17'h13006:	data_out=16'h89fc;
17'h13007:	data_out=16'h89fa;
17'h13008:	data_out=16'h89f2;
17'h13009:	data_out=16'h89f4;
17'h1300a:	data_out=16'h9fa;
17'h1300b:	data_out=16'h89e9;
17'h1300c:	data_out=16'h89fb;
17'h1300d:	data_out=16'h89c9;
17'h1300e:	data_out=16'h9ff;
17'h1300f:	data_out=16'h89ec;
17'h13010:	data_out=16'h89e9;
17'h13011:	data_out=16'h86f3;
17'h13012:	data_out=16'h89f5;
17'h13013:	data_out=16'h89b7;
17'h13014:	data_out=16'h899a;
17'h13015:	data_out=16'ha00;
17'h13016:	data_out=16'h53a;
17'h13017:	data_out=16'h89be;
17'h13018:	data_out=16'h89ef;
17'h13019:	data_out=16'h9f0;
17'h1301a:	data_out=16'ha00;
17'h1301b:	data_out=16'h89cd;
17'h1301c:	data_out=16'h83b3;
17'h1301d:	data_out=16'h89fa;
17'h1301e:	data_out=16'h89ad;
17'h1301f:	data_out=16'h88a6;
17'h13020:	data_out=16'h8978;
17'h13021:	data_out=16'h9ff;
17'h13022:	data_out=16'h56c;
17'h13023:	data_out=16'h9d8;
17'h13024:	data_out=16'h9d9;
17'h13025:	data_out=16'h894d;
17'h13026:	data_out=16'h89b7;
17'h13027:	data_out=16'h89ad;
17'h13028:	data_out=16'h9ff;
17'h13029:	data_out=16'ha00;
17'h1302a:	data_out=16'h89ee;
17'h1302b:	data_out=16'h9f3;
17'h1302c:	data_out=16'ha00;
17'h1302d:	data_out=16'h8a00;
17'h1302e:	data_out=16'h89f2;
17'h1302f:	data_out=16'h89ec;
17'h13030:	data_out=16'ha00;
17'h13031:	data_out=16'h9e8;
17'h13032:	data_out=16'h9cd;
17'h13033:	data_out=16'h89e5;
17'h13034:	data_out=16'h89ff;
17'h13035:	data_out=16'h9f4;
17'h13036:	data_out=16'h89ec;
17'h13037:	data_out=16'h89dc;
17'h13038:	data_out=16'h89fb;
17'h13039:	data_out=16'h89ea;
17'h1303a:	data_out=16'h89d7;
17'h1303b:	data_out=16'h9eb;
17'h1303c:	data_out=16'h8458;
17'h1303d:	data_out=16'h4c5;
17'h1303e:	data_out=16'h9ff;
17'h1303f:	data_out=16'ha00;
17'h13040:	data_out=16'h8281;
17'h13041:	data_out=16'h890c;
17'h13042:	data_out=16'h89fe;
17'h13043:	data_out=16'h751;
17'h13044:	data_out=16'ha00;
17'h13045:	data_out=16'ha00;
17'h13046:	data_out=16'h839f;
17'h13047:	data_out=16'h89f8;
17'h13048:	data_out=16'h89f5;
17'h13049:	data_out=16'h82e9;
17'h1304a:	data_out=16'h89f3;
17'h1304b:	data_out=16'h89ff;
17'h1304c:	data_out=16'h89fb;
17'h1304d:	data_out=16'h9ef;
17'h1304e:	data_out=16'h89fe;
17'h1304f:	data_out=16'h89fe;
17'h13050:	data_out=16'h5a3;
17'h13051:	data_out=16'ha00;
17'h13052:	data_out=16'h9c3;
17'h13053:	data_out=16'h89c2;
17'h13054:	data_out=16'h89d9;
17'h13055:	data_out=16'h88fb;
17'h13056:	data_out=16'h9f0;
17'h13057:	data_out=16'h9fd;
17'h13058:	data_out=16'h9d;
17'h13059:	data_out=16'h984;
17'h1305a:	data_out=16'h89ed;
17'h1305b:	data_out=16'ha00;
17'h1305c:	data_out=16'h86f9;
17'h1305d:	data_out=16'h8933;
17'h1305e:	data_out=16'h89f3;
17'h1305f:	data_out=16'h89f6;
17'h13060:	data_out=16'h89fb;
17'h13061:	data_out=16'ha00;
17'h13062:	data_out=16'h89f0;
17'h13063:	data_out=16'h89e5;
17'h13064:	data_out=16'h8a00;
17'h13065:	data_out=16'h88b4;
17'h13066:	data_out=16'h9fa;
17'h13067:	data_out=16'ha00;
17'h13068:	data_out=16'h9ff;
17'h13069:	data_out=16'h89f6;
17'h1306a:	data_out=16'h9ff;
17'h1306b:	data_out=16'h756;
17'h1306c:	data_out=16'h8886;
17'h1306d:	data_out=16'h89e6;
17'h1306e:	data_out=16'h9ff;
17'h1306f:	data_out=16'ha00;
17'h13070:	data_out=16'h9ff;
17'h13071:	data_out=16'h89d9;
17'h13072:	data_out=16'h992;
17'h13073:	data_out=16'ha00;
17'h13074:	data_out=16'h9fc;
17'h13075:	data_out=16'ha00;
17'h13076:	data_out=16'ha00;
17'h13077:	data_out=16'h89f0;
17'h13078:	data_out=16'h765;
17'h13079:	data_out=16'h83c5;
17'h1307a:	data_out=16'h89dd;
17'h1307b:	data_out=16'h9ff;
17'h1307c:	data_out=16'h89f0;
17'h1307d:	data_out=16'h831b;
17'h1307e:	data_out=16'h89fe;
17'h1307f:	data_out=16'h9fd;
17'h13080:	data_out=16'h9ff;
17'h13081:	data_out=16'h88cb;
17'h13082:	data_out=16'h896d;
17'h13083:	data_out=16'h897e;
17'h13084:	data_out=16'ha00;
17'h13085:	data_out=16'ha00;
17'h13086:	data_out=16'h89fd;
17'h13087:	data_out=16'h89fb;
17'h13088:	data_out=16'h89ea;
17'h13089:	data_out=16'h89b8;
17'h1308a:	data_out=16'h9fc;
17'h1308b:	data_out=16'h89f5;
17'h1308c:	data_out=16'h89fb;
17'h1308d:	data_out=16'h8998;
17'h1308e:	data_out=16'ha00;
17'h1308f:	data_out=16'h89be;
17'h13090:	data_out=16'h89d0;
17'h13091:	data_out=16'h6a7;
17'h13092:	data_out=16'h89e9;
17'h13093:	data_out=16'h891d;
17'h13094:	data_out=16'h89a3;
17'h13095:	data_out=16'ha00;
17'h13096:	data_out=16'ha00;
17'h13097:	data_out=16'h89d5;
17'h13098:	data_out=16'h9f3;
17'h13099:	data_out=16'h9e1;
17'h1309a:	data_out=16'ha00;
17'h1309b:	data_out=16'h8992;
17'h1309c:	data_out=16'h9ff;
17'h1309d:	data_out=16'h86c6;
17'h1309e:	data_out=16'h895a;
17'h1309f:	data_out=16'h8065;
17'h130a0:	data_out=16'h9f4;
17'h130a1:	data_out=16'ha00;
17'h130a2:	data_out=16'ha00;
17'h130a3:	data_out=16'h9fe;
17'h130a4:	data_out=16'h9ff;
17'h130a5:	data_out=16'h77c;
17'h130a6:	data_out=16'h88d3;
17'h130a7:	data_out=16'h8998;
17'h130a8:	data_out=16'ha00;
17'h130a9:	data_out=16'ha00;
17'h130aa:	data_out=16'h89d7;
17'h130ab:	data_out=16'h9fe;
17'h130ac:	data_out=16'ha00;
17'h130ad:	data_out=16'h8a00;
17'h130ae:	data_out=16'h89fb;
17'h130af:	data_out=16'h89df;
17'h130b0:	data_out=16'h9ff;
17'h130b1:	data_out=16'h1c1;
17'h130b2:	data_out=16'h9d3;
17'h130b3:	data_out=16'h89d0;
17'h130b4:	data_out=16'h89fe;
17'h130b5:	data_out=16'ha00;
17'h130b6:	data_out=16'h89b3;
17'h130b7:	data_out=16'h8974;
17'h130b8:	data_out=16'h69;
17'h130b9:	data_out=16'h89bb;
17'h130ba:	data_out=16'h89bd;
17'h130bb:	data_out=16'h9ec;
17'h130bc:	data_out=16'h85c4;
17'h130bd:	data_out=16'ha00;
17'h130be:	data_out=16'ha00;
17'h130bf:	data_out=16'ha00;
17'h130c0:	data_out=16'ha00;
17'h130c1:	data_out=16'h88ea;
17'h130c2:	data_out=16'h89fd;
17'h130c3:	data_out=16'h82cd;
17'h130c4:	data_out=16'ha00;
17'h130c5:	data_out=16'ha00;
17'h130c6:	data_out=16'h80e1;
17'h130c7:	data_out=16'h89ed;
17'h130c8:	data_out=16'h89fa;
17'h130c9:	data_out=16'ha00;
17'h130ca:	data_out=16'h89f7;
17'h130cb:	data_out=16'h89fe;
17'h130cc:	data_out=16'h8983;
17'h130cd:	data_out=16'ha00;
17'h130ce:	data_out=16'h8500;
17'h130cf:	data_out=16'h81a5;
17'h130d0:	data_out=16'h9f1;
17'h130d1:	data_out=16'h94c;
17'h130d2:	data_out=16'h9fe;
17'h130d3:	data_out=16'h89a6;
17'h130d4:	data_out=16'h8965;
17'h130d5:	data_out=16'h8428;
17'h130d6:	data_out=16'ha00;
17'h130d7:	data_out=16'ha00;
17'h130d8:	data_out=16'h7e3;
17'h130d9:	data_out=16'h9fb;
17'h130da:	data_out=16'h89fb;
17'h130db:	data_out=16'ha00;
17'h130dc:	data_out=16'h88e4;
17'h130dd:	data_out=16'h86e2;
17'h130de:	data_out=16'h89f2;
17'h130df:	data_out=16'h87d2;
17'h130e0:	data_out=16'h89bb;
17'h130e1:	data_out=16'ha00;
17'h130e2:	data_out=16'h89ca;
17'h130e3:	data_out=16'h89e6;
17'h130e4:	data_out=16'h88fa;
17'h130e5:	data_out=16'h89fe;
17'h130e6:	data_out=16'h9f3;
17'h130e7:	data_out=16'ha00;
17'h130e8:	data_out=16'ha00;
17'h130e9:	data_out=16'h89f3;
17'h130ea:	data_out=16'ha00;
17'h130eb:	data_out=16'h9f7;
17'h130ec:	data_out=16'h9ff;
17'h130ed:	data_out=16'h89e2;
17'h130ee:	data_out=16'ha00;
17'h130ef:	data_out=16'h83f2;
17'h130f0:	data_out=16'ha00;
17'h130f1:	data_out=16'h89bf;
17'h130f2:	data_out=16'h9db;
17'h130f3:	data_out=16'ha00;
17'h130f4:	data_out=16'h9fa;
17'h130f5:	data_out=16'h9ff;
17'h130f6:	data_out=16'ha00;
17'h130f7:	data_out=16'h82e9;
17'h130f8:	data_out=16'h16;
17'h130f9:	data_out=16'hf4;
17'h130fa:	data_out=16'h89c9;
17'h130fb:	data_out=16'ha00;
17'h130fc:	data_out=16'h60a;
17'h130fd:	data_out=16'h204;
17'h130fe:	data_out=16'h89ff;
17'h130ff:	data_out=16'ha00;
17'h13100:	data_out=16'h9f4;
17'h13101:	data_out=16'hff;
17'h13102:	data_out=16'h89a4;
17'h13103:	data_out=16'h89ce;
17'h13104:	data_out=16'ha00;
17'h13105:	data_out=16'h871;
17'h13106:	data_out=16'h89fa;
17'h13107:	data_out=16'h89fe;
17'h13108:	data_out=16'h89e3;
17'h13109:	data_out=16'h715;
17'h1310a:	data_out=16'h9ff;
17'h1310b:	data_out=16'h89f0;
17'h1310c:	data_out=16'h89ff;
17'h1310d:	data_out=16'h89f0;
17'h1310e:	data_out=16'ha00;
17'h1310f:	data_out=16'h89d9;
17'h13110:	data_out=16'h9f4;
17'h13111:	data_out=16'h9e4;
17'h13112:	data_out=16'h89fa;
17'h13113:	data_out=16'h89b7;
17'h13114:	data_out=16'h89e0;
17'h13115:	data_out=16'ha00;
17'h13116:	data_out=16'h938;
17'h13117:	data_out=16'h89fd;
17'h13118:	data_out=16'ha00;
17'h13119:	data_out=16'h9f4;
17'h1311a:	data_out=16'h9fd;
17'h1311b:	data_out=16'h89c8;
17'h1311c:	data_out=16'h9da;
17'h1311d:	data_out=16'h3c9;
17'h1311e:	data_out=16'h88d2;
17'h1311f:	data_out=16'h810e;
17'h13120:	data_out=16'h9f1;
17'h13121:	data_out=16'ha00;
17'h13122:	data_out=16'ha00;
17'h13123:	data_out=16'ha00;
17'h13124:	data_out=16'ha00;
17'h13125:	data_out=16'ha00;
17'h13126:	data_out=16'h116;
17'h13127:	data_out=16'h4de;
17'h13128:	data_out=16'ha00;
17'h13129:	data_out=16'h8b8;
17'h1312a:	data_out=16'h89ea;
17'h1312b:	data_out=16'ha00;
17'h1312c:	data_out=16'h9fb;
17'h1312d:	data_out=16'h8341;
17'h1312e:	data_out=16'h89fe;
17'h1312f:	data_out=16'h89ea;
17'h13130:	data_out=16'h9fb;
17'h13131:	data_out=16'h886a;
17'h13132:	data_out=16'h9b5;
17'h13133:	data_out=16'h89d7;
17'h13134:	data_out=16'h89e8;
17'h13135:	data_out=16'ha00;
17'h13136:	data_out=16'h89a4;
17'h13137:	data_out=16'h89af;
17'h13138:	data_out=16'h9b4;
17'h13139:	data_out=16'h8981;
17'h1313a:	data_out=16'h9f8;
17'h1313b:	data_out=16'h9c6;
17'h1313c:	data_out=16'h88de;
17'h1313d:	data_out=16'ha00;
17'h1313e:	data_out=16'ha00;
17'h1313f:	data_out=16'h93e;
17'h13140:	data_out=16'ha00;
17'h13141:	data_out=16'h8978;
17'h13142:	data_out=16'h89ff;
17'h13143:	data_out=16'h897a;
17'h13144:	data_out=16'ha00;
17'h13145:	data_out=16'ha00;
17'h13146:	data_out=16'h9ad;
17'h13147:	data_out=16'h21a;
17'h13148:	data_out=16'h89fd;
17'h13149:	data_out=16'ha00;
17'h1314a:	data_out=16'h89fc;
17'h1314b:	data_out=16'h8a00;
17'h1314c:	data_out=16'h8200;
17'h1314d:	data_out=16'ha00;
17'h1314e:	data_out=16'h872b;
17'h1314f:	data_out=16'h9fe;
17'h13150:	data_out=16'h99b;
17'h13151:	data_out=16'h88ae;
17'h13152:	data_out=16'ha00;
17'h13153:	data_out=16'h89bd;
17'h13154:	data_out=16'h9e5;
17'h13155:	data_out=16'h898b;
17'h13156:	data_out=16'ha00;
17'h13157:	data_out=16'ha00;
17'h13158:	data_out=16'h5c9;
17'h13159:	data_out=16'ha00;
17'h1315a:	data_out=16'h89fd;
17'h1315b:	data_out=16'ha00;
17'h1315c:	data_out=16'h89eb;
17'h1315d:	data_out=16'h850b;
17'h1315e:	data_out=16'h89fc;
17'h1315f:	data_out=16'h7c9;
17'h13160:	data_out=16'h89c9;
17'h13161:	data_out=16'ha00;
17'h13162:	data_out=16'h89f5;
17'h13163:	data_out=16'h89f7;
17'h13164:	data_out=16'h6fc;
17'h13165:	data_out=16'h89f5;
17'h13166:	data_out=16'h252;
17'h13167:	data_out=16'ha00;
17'h13168:	data_out=16'ha00;
17'h13169:	data_out=16'h89f8;
17'h1316a:	data_out=16'ha00;
17'h1316b:	data_out=16'h9e8;
17'h1316c:	data_out=16'h9fb;
17'h1316d:	data_out=16'h89ef;
17'h1316e:	data_out=16'ha00;
17'h1316f:	data_out=16'h89e3;
17'h13170:	data_out=16'ha00;
17'h13171:	data_out=16'h89f9;
17'h13172:	data_out=16'h9fb;
17'h13173:	data_out=16'h9f9;
17'h13174:	data_out=16'h9fe;
17'h13175:	data_out=16'h467;
17'h13176:	data_out=16'ha00;
17'h13177:	data_out=16'h8c0;
17'h13178:	data_out=16'h8774;
17'h13179:	data_out=16'h8214;
17'h1317a:	data_out=16'h89f5;
17'h1317b:	data_out=16'ha00;
17'h1317c:	data_out=16'h9b2;
17'h1317d:	data_out=16'h8223;
17'h1317e:	data_out=16'h410;
17'h1317f:	data_out=16'ha00;
17'h13180:	data_out=16'ha00;
17'h13181:	data_out=16'h82e;
17'h13182:	data_out=16'h89df;
17'h13183:	data_out=16'h47c;
17'h13184:	data_out=16'ha00;
17'h13185:	data_out=16'h9f3;
17'h13186:	data_out=16'h8742;
17'h13187:	data_out=16'h845d;
17'h13188:	data_out=16'h89e0;
17'h13189:	data_out=16'h9b5;
17'h1318a:	data_out=16'h9fc;
17'h1318b:	data_out=16'h882b;
17'h1318c:	data_out=16'h8a00;
17'h1318d:	data_out=16'h89fa;
17'h1318e:	data_out=16'ha00;
17'h1318f:	data_out=16'h89b5;
17'h13190:	data_out=16'ha00;
17'h13191:	data_out=16'h9fb;
17'h13192:	data_out=16'h89fc;
17'h13193:	data_out=16'h507;
17'h13194:	data_out=16'h213;
17'h13195:	data_out=16'ha00;
17'h13196:	data_out=16'h9fa;
17'h13197:	data_out=16'h8a00;
17'h13198:	data_out=16'ha00;
17'h13199:	data_out=16'h591;
17'h1319a:	data_out=16'h9fa;
17'h1319b:	data_out=16'h89e8;
17'h1319c:	data_out=16'h9f5;
17'h1319d:	data_out=16'h908;
17'h1319e:	data_out=16'h19d;
17'h1319f:	data_out=16'h8c7;
17'h131a0:	data_out=16'h9ff;
17'h131a1:	data_out=16'ha00;
17'h131a2:	data_out=16'ha00;
17'h131a3:	data_out=16'ha00;
17'h131a4:	data_out=16'ha00;
17'h131a5:	data_out=16'ha00;
17'h131a6:	data_out=16'h866;
17'h131a7:	data_out=16'h9fd;
17'h131a8:	data_out=16'ha00;
17'h131a9:	data_out=16'h2d2;
17'h131aa:	data_out=16'h89f6;
17'h131ab:	data_out=16'ha00;
17'h131ac:	data_out=16'ha00;
17'h131ad:	data_out=16'h8105;
17'h131ae:	data_out=16'h8a00;
17'h131af:	data_out=16'h9cb;
17'h131b0:	data_out=16'h8999;
17'h131b1:	data_out=16'h87a2;
17'h131b2:	data_out=16'h8933;
17'h131b3:	data_out=16'h9ea;
17'h131b4:	data_out=16'h687;
17'h131b5:	data_out=16'h9fe;
17'h131b6:	data_out=16'h345;
17'h131b7:	data_out=16'h89e6;
17'h131b8:	data_out=16'h9ea;
17'h131b9:	data_out=16'h9f4;
17'h131ba:	data_out=16'ha00;
17'h131bb:	data_out=16'h93a;
17'h131bc:	data_out=16'h89dd;
17'h131bd:	data_out=16'ha00;
17'h131be:	data_out=16'ha00;
17'h131bf:	data_out=16'h9f4;
17'h131c0:	data_out=16'h9f9;
17'h131c1:	data_out=16'h8996;
17'h131c2:	data_out=16'h8a00;
17'h131c3:	data_out=16'h89f9;
17'h131c4:	data_out=16'h9fe;
17'h131c5:	data_out=16'ha00;
17'h131c6:	data_out=16'h57b;
17'h131c7:	data_out=16'h9f6;
17'h131c8:	data_out=16'h89ff;
17'h131c9:	data_out=16'ha00;
17'h131ca:	data_out=16'h89fe;
17'h131cb:	data_out=16'h8a00;
17'h131cc:	data_out=16'h81e2;
17'h131cd:	data_out=16'ha00;
17'h131ce:	data_out=16'h8818;
17'h131cf:	data_out=16'ha00;
17'h131d0:	data_out=16'h9f3;
17'h131d1:	data_out=16'h49;
17'h131d2:	data_out=16'ha00;
17'h131d3:	data_out=16'h89df;
17'h131d4:	data_out=16'h9fa;
17'h131d5:	data_out=16'h82fe;
17'h131d6:	data_out=16'ha00;
17'h131d7:	data_out=16'ha00;
17'h131d8:	data_out=16'h820d;
17'h131d9:	data_out=16'h9fe;
17'h131da:	data_out=16'h8a00;
17'h131db:	data_out=16'ha00;
17'h131dc:	data_out=16'h878a;
17'h131dd:	data_out=16'h9fa;
17'h131de:	data_out=16'h943;
17'h131df:	data_out=16'h9fe;
17'h131e0:	data_out=16'h8837;
17'h131e1:	data_out=16'h9f7;
17'h131e2:	data_out=16'h89fa;
17'h131e3:	data_out=16'h8ee;
17'h131e4:	data_out=16'ha00;
17'h131e5:	data_out=16'h81d2;
17'h131e6:	data_out=16'h557;
17'h131e7:	data_out=16'ha00;
17'h131e8:	data_out=16'ha00;
17'h131e9:	data_out=16'h89f6;
17'h131ea:	data_out=16'ha00;
17'h131eb:	data_out=16'h9f9;
17'h131ec:	data_out=16'ha00;
17'h131ed:	data_out=16'h964;
17'h131ee:	data_out=16'ha00;
17'h131ef:	data_out=16'h8a00;
17'h131f0:	data_out=16'ha00;
17'h131f1:	data_out=16'h89ff;
17'h131f2:	data_out=16'h9fe;
17'h131f3:	data_out=16'h9f8;
17'h131f4:	data_out=16'h89d6;
17'h131f5:	data_out=16'h89e9;
17'h131f6:	data_out=16'ha00;
17'h131f7:	data_out=16'h9f3;
17'h131f8:	data_out=16'h8941;
17'h131f9:	data_out=16'h861f;
17'h131fa:	data_out=16'h6d0;
17'h131fb:	data_out=16'ha00;
17'h131fc:	data_out=16'h9ff;
17'h131fd:	data_out=16'h4b3;
17'h131fe:	data_out=16'h8f4;
17'h131ff:	data_out=16'ha00;
17'h13200:	data_out=16'ha00;
17'h13201:	data_out=16'h3d7;
17'h13202:	data_out=16'h89b3;
17'h13203:	data_out=16'ha00;
17'h13204:	data_out=16'h9fc;
17'h13205:	data_out=16'h8d8;
17'h13206:	data_out=16'h87a;
17'h13207:	data_out=16'h2ec;
17'h13208:	data_out=16'h89ee;
17'h13209:	data_out=16'h9f9;
17'h1320a:	data_out=16'h68b;
17'h1320b:	data_out=16'h1b5;
17'h1320c:	data_out=16'h8a00;
17'h1320d:	data_out=16'h500;
17'h1320e:	data_out=16'h25a;
17'h1320f:	data_out=16'h8650;
17'h13210:	data_out=16'ha00;
17'h13211:	data_out=16'h5c5;
17'h13212:	data_out=16'h829c;
17'h13213:	data_out=16'ha00;
17'h13214:	data_out=16'h9fa;
17'h13215:	data_out=16'ha00;
17'h13216:	data_out=16'ha00;
17'h13217:	data_out=16'h9f3;
17'h13218:	data_out=16'h69c;
17'h13219:	data_out=16'he1;
17'h1321a:	data_out=16'h94b;
17'h1321b:	data_out=16'h898e;
17'h1321c:	data_out=16'h9ff;
17'h1321d:	data_out=16'h917;
17'h1321e:	data_out=16'ha00;
17'h1321f:	data_out=16'h978;
17'h13220:	data_out=16'ha00;
17'h13221:	data_out=16'h241;
17'h13222:	data_out=16'h9ff;
17'h13223:	data_out=16'h51;
17'h13224:	data_out=16'h56;
17'h13225:	data_out=16'ha00;
17'h13226:	data_out=16'h9f8;
17'h13227:	data_out=16'h9f8;
17'h13228:	data_out=16'h239;
17'h13229:	data_out=16'h9fe;
17'h1322a:	data_out=16'h8383;
17'h1322b:	data_out=16'h9fe;
17'h1322c:	data_out=16'ha00;
17'h1322d:	data_out=16'h9fe;
17'h1322e:	data_out=16'h80d5;
17'h1322f:	data_out=16'h9f9;
17'h13230:	data_out=16'h89fb;
17'h13231:	data_out=16'h80ca;
17'h13232:	data_out=16'h8a00;
17'h13233:	data_out=16'h9fd;
17'h13234:	data_out=16'h8c1;
17'h13235:	data_out=16'h81e1;
17'h13236:	data_out=16'h378;
17'h13237:	data_out=16'h89f2;
17'h13238:	data_out=16'h9ed;
17'h13239:	data_out=16'ha00;
17'h1323a:	data_out=16'h9ff;
17'h1323b:	data_out=16'h3c7;
17'h1323c:	data_out=16'h888e;
17'h1323d:	data_out=16'ha00;
17'h1323e:	data_out=16'h238;
17'h1323f:	data_out=16'h8ea;
17'h13240:	data_out=16'h9f6;
17'h13241:	data_out=16'h858e;
17'h13242:	data_out=16'h87fa;
17'h13243:	data_out=16'ha00;
17'h13244:	data_out=16'h9f7;
17'h13245:	data_out=16'ha00;
17'h13246:	data_out=16'hcc;
17'h13247:	data_out=16'h9fd;
17'h13248:	data_out=16'h310;
17'h13249:	data_out=16'ha00;
17'h1324a:	data_out=16'h8a00;
17'h1324b:	data_out=16'h89fe;
17'h1324c:	data_out=16'h9fc;
17'h1324d:	data_out=16'h9fe;
17'h1324e:	data_out=16'h8987;
17'h1324f:	data_out=16'h9fd;
17'h13250:	data_out=16'ha00;
17'h13251:	data_out=16'h9fe;
17'h13252:	data_out=16'h7c2;
17'h13253:	data_out=16'h8a00;
17'h13254:	data_out=16'h9fb;
17'h13255:	data_out=16'h2ae;
17'h13256:	data_out=16'h9fe;
17'h13257:	data_out=16'ha00;
17'h13258:	data_out=16'h869f;
17'h13259:	data_out=16'h9f9;
17'h1325a:	data_out=16'h89fe;
17'h1325b:	data_out=16'h9fb;
17'h1325c:	data_out=16'h8361;
17'h1325d:	data_out=16'h9fe;
17'h1325e:	data_out=16'h9f6;
17'h1325f:	data_out=16'h75a;
17'h13260:	data_out=16'h672;
17'h13261:	data_out=16'h976;
17'h13262:	data_out=16'h860c;
17'h13263:	data_out=16'h9f8;
17'h13264:	data_out=16'ha00;
17'h13265:	data_out=16'h89b;
17'h13266:	data_out=16'h284;
17'h13267:	data_out=16'h9fd;
17'h13268:	data_out=16'h246;
17'h13269:	data_out=16'h89e8;
17'h1326a:	data_out=16'h270;
17'h1326b:	data_out=16'ha00;
17'h1326c:	data_out=16'ha00;
17'h1326d:	data_out=16'h9f9;
17'h1326e:	data_out=16'h26f;
17'h1326f:	data_out=16'h3a7;
17'h13270:	data_out=16'h25f;
17'h13271:	data_out=16'h8a00;
17'h13272:	data_out=16'ha00;
17'h13273:	data_out=16'h9f5;
17'h13274:	data_out=16'h89fc;
17'h13275:	data_out=16'h8a00;
17'h13276:	data_out=16'h9ff;
17'h13277:	data_out=16'h9fa;
17'h13278:	data_out=16'h781;
17'h13279:	data_out=16'h86d3;
17'h1327a:	data_out=16'h9f7;
17'h1327b:	data_out=16'h235;
17'h1327c:	data_out=16'h1d3;
17'h1327d:	data_out=16'h9fc;
17'h1327e:	data_out=16'h9fd;
17'h1327f:	data_out=16'ha00;
17'h13280:	data_out=16'ha00;
17'h13281:	data_out=16'h5f1;
17'h13282:	data_out=16'h81d6;
17'h13283:	data_out=16'h9ff;
17'h13284:	data_out=16'h771;
17'h13285:	data_out=16'h9fa;
17'h13286:	data_out=16'hd0;
17'h13287:	data_out=16'h5e5;
17'h13288:	data_out=16'h80ec;
17'h13289:	data_out=16'ha00;
17'h1328a:	data_out=16'h7ac;
17'h1328b:	data_out=16'h8858;
17'h1328c:	data_out=16'h8a00;
17'h1328d:	data_out=16'h62f;
17'h1328e:	data_out=16'h10e;
17'h1328f:	data_out=16'h80f3;
17'h13290:	data_out=16'ha00;
17'h13291:	data_out=16'h1b6;
17'h13292:	data_out=16'h843e;
17'h13293:	data_out=16'ha00;
17'h13294:	data_out=16'h730;
17'h13295:	data_out=16'ha00;
17'h13296:	data_out=16'ha00;
17'h13297:	data_out=16'h2c9;
17'h13298:	data_out=16'h3a3;
17'h13299:	data_out=16'h808a;
17'h1329a:	data_out=16'h5a5;
17'h1329b:	data_out=16'h82f4;
17'h1329c:	data_out=16'ha00;
17'h1329d:	data_out=16'h71e;
17'h1329e:	data_out=16'h724;
17'h1329f:	data_out=16'h9d9;
17'h132a0:	data_out=16'ha00;
17'h132a1:	data_out=16'h103;
17'h132a2:	data_out=16'ha00;
17'h132a3:	data_out=16'h84ca;
17'h132a4:	data_out=16'h84c8;
17'h132a5:	data_out=16'h96f;
17'h132a6:	data_out=16'h5cd;
17'h132a7:	data_out=16'h749;
17'h132a8:	data_out=16'hf6;
17'h132a9:	data_out=16'h85a;
17'h132aa:	data_out=16'h8327;
17'h132ab:	data_out=16'h84d;
17'h132ac:	data_out=16'ha00;
17'h132ad:	data_out=16'haf;
17'h132ae:	data_out=16'h80a3;
17'h132af:	data_out=16'ha00;
17'h132b0:	data_out=16'h82c5;
17'h132b1:	data_out=16'h780;
17'h132b2:	data_out=16'h8307;
17'h132b3:	data_out=16'ha00;
17'h132b4:	data_out=16'h67d;
17'h132b5:	data_out=16'h12a;
17'h132b6:	data_out=16'h32f;
17'h132b7:	data_out=16'h82ac;
17'h132b8:	data_out=16'h8c2;
17'h132b9:	data_out=16'ha00;
17'h132ba:	data_out=16'ha00;
17'h132bb:	data_out=16'h96c;
17'h132bc:	data_out=16'h840c;
17'h132bd:	data_out=16'ha00;
17'h132be:	data_out=16'hf5;
17'h132bf:	data_out=16'h9fd;
17'h132c0:	data_out=16'ha00;
17'h132c1:	data_out=16'h76;
17'h132c2:	data_out=16'h8891;
17'h132c3:	data_out=16'h2eb;
17'h132c4:	data_out=16'ha00;
17'h132c5:	data_out=16'ha00;
17'h132c6:	data_out=16'h80bd;
17'h132c7:	data_out=16'ha00;
17'h132c8:	data_out=16'h28;
17'h132c9:	data_out=16'ha00;
17'h132ca:	data_out=16'h2f2;
17'h132cb:	data_out=16'h8a00;
17'h132cc:	data_out=16'h1ef;
17'h132cd:	data_out=16'ha00;
17'h132ce:	data_out=16'h837b;
17'h132cf:	data_out=16'h493;
17'h132d0:	data_out=16'ha00;
17'h132d1:	data_out=16'h6e8;
17'h132d2:	data_out=16'h829e;
17'h132d3:	data_out=16'h8197;
17'h132d4:	data_out=16'ha00;
17'h132d5:	data_out=16'h161;
17'h132d6:	data_out=16'h9fe;
17'h132d7:	data_out=16'ha00;
17'h132d8:	data_out=16'h805c;
17'h132d9:	data_out=16'ha00;
17'h132da:	data_out=16'h8a00;
17'h132db:	data_out=16'ha00;
17'h132dc:	data_out=16'h48d;
17'h132dd:	data_out=16'h6a9;
17'h132de:	data_out=16'h9ff;
17'h132df:	data_out=16'h3d4;
17'h132e0:	data_out=16'h8153;
17'h132e1:	data_out=16'h9ff;
17'h132e2:	data_out=16'h8681;
17'h132e3:	data_out=16'h962;
17'h132e4:	data_out=16'h983;
17'h132e5:	data_out=16'hee;
17'h132e6:	data_out=16'h39;
17'h132e7:	data_out=16'h34a;
17'h132e8:	data_out=16'h100;
17'h132e9:	data_out=16'h8274;
17'h132ea:	data_out=16'h115;
17'h132eb:	data_out=16'ha00;
17'h132ec:	data_out=16'h93f;
17'h132ed:	data_out=16'h9c5;
17'h132ee:	data_out=16'h115;
17'h132ef:	data_out=16'h6ee;
17'h132f0:	data_out=16'h110;
17'h132f1:	data_out=16'h837c;
17'h132f2:	data_out=16'ha00;
17'h132f3:	data_out=16'h9ff;
17'h132f4:	data_out=16'h82ed;
17'h132f5:	data_out=16'h8874;
17'h132f6:	data_out=16'h5cf;
17'h132f7:	data_out=16'ha00;
17'h132f8:	data_out=16'h176;
17'h132f9:	data_out=16'h80f9;
17'h132fa:	data_out=16'h7c7;
17'h132fb:	data_out=16'hf4;
17'h132fc:	data_out=16'h2ae;
17'h132fd:	data_out=16'he5;
17'h132fe:	data_out=16'ha00;
17'h132ff:	data_out=16'ha00;
17'h13300:	data_out=16'h440;
17'h13301:	data_out=16'h30a;
17'h13302:	data_out=16'h809f;
17'h13303:	data_out=16'hf9;
17'h13304:	data_out=16'h1d7;
17'h13305:	data_out=16'h4f;
17'h13306:	data_out=16'h8052;
17'h13307:	data_out=16'h350;
17'h13308:	data_out=16'h55;
17'h13309:	data_out=16'h3db;
17'h1330a:	data_out=16'h3e5;
17'h1330b:	data_out=16'h800f;
17'h1330c:	data_out=16'h28c;
17'h1330d:	data_out=16'h8032;
17'h1330e:	data_out=16'h8001;
17'h1330f:	data_out=16'h8038;
17'h13310:	data_out=16'h211;
17'h13311:	data_out=16'h33c;
17'h13312:	data_out=16'h83;
17'h13313:	data_out=16'h106;
17'h13314:	data_out=16'h8007;
17'h13315:	data_out=16'h19f;
17'h13316:	data_out=16'h14f;
17'h13317:	data_out=16'h8084;
17'h13318:	data_out=16'hab;
17'h13319:	data_out=16'h1ca;
17'h1331a:	data_out=16'h15d;
17'h1331b:	data_out=16'h8011;
17'h1331c:	data_out=16'h1b1;
17'h1331d:	data_out=16'h3a8;
17'h1331e:	data_out=16'h44;
17'h1331f:	data_out=16'h65;
17'h13320:	data_out=16'h360;
17'h13321:	data_out=16'h800b;
17'h13322:	data_out=16'h329;
17'h13323:	data_out=16'h1a1;
17'h13324:	data_out=16'h1a4;
17'h13325:	data_out=16'h2b5;
17'h13326:	data_out=16'h291;
17'h13327:	data_out=16'h339;
17'h13328:	data_out=16'h9;
17'h13329:	data_out=16'h8043;
17'h1332a:	data_out=16'h8c;
17'h1332b:	data_out=16'h303;
17'h1332c:	data_out=16'h170;
17'h1332d:	data_out=16'h1fd;
17'h1332e:	data_out=16'h808a;
17'h1332f:	data_out=16'h221;
17'h13330:	data_out=16'h96;
17'h13331:	data_out=16'h50f;
17'h13332:	data_out=16'ha4;
17'h13333:	data_out=16'h7c;
17'h13334:	data_out=16'h4b3;
17'h13335:	data_out=16'h247;
17'h13336:	data_out=16'h2c;
17'h13337:	data_out=16'h80a2;
17'h13338:	data_out=16'h236;
17'h13339:	data_out=16'h72;
17'h1333a:	data_out=16'h304;
17'h1333b:	data_out=16'h372;
17'h1333c:	data_out=16'h8127;
17'h1333d:	data_out=16'h477;
17'h1333e:	data_out=16'h8003;
17'h1333f:	data_out=16'h86;
17'h13340:	data_out=16'h19a;
17'h13341:	data_out=16'h80c2;
17'h13342:	data_out=16'hb9;
17'h13343:	data_out=16'h8100;
17'h13344:	data_out=16'h2fa;
17'h13345:	data_out=16'h1a1;
17'h13346:	data_out=16'h8029;
17'h13347:	data_out=16'h277;
17'h13348:	data_out=16'h99;
17'h13349:	data_out=16'h2be;
17'h1334a:	data_out=16'he3;
17'h1334b:	data_out=16'he6;
17'h1334c:	data_out=16'ha0;
17'h1334d:	data_out=16'h38a;
17'h1334e:	data_out=16'h800e;
17'h1334f:	data_out=16'h148;
17'h13350:	data_out=16'hd9;
17'h13351:	data_out=16'h807c;
17'h13352:	data_out=16'h201;
17'h13353:	data_out=16'h1d8;
17'h13354:	data_out=16'h241;
17'h13355:	data_out=16'h81bc;
17'h13356:	data_out=16'h1eb;
17'h13357:	data_out=16'h1fa;
17'h13358:	data_out=16'h81aa;
17'h13359:	data_out=16'h1bd;
17'h1335a:	data_out=16'h81df;
17'h1335b:	data_out=16'h8e;
17'h1335c:	data_out=16'h143;
17'h1335d:	data_out=16'he1;
17'h1335e:	data_out=16'h1a4;
17'h1335f:	data_out=16'h120;
17'h13360:	data_out=16'h308;
17'h13361:	data_out=16'h2a1;
17'h13362:	data_out=16'h8204;
17'h13363:	data_out=16'h65;
17'h13364:	data_out=16'h4da;
17'h13365:	data_out=16'h2b1;
17'h13366:	data_out=16'h200;
17'h13367:	data_out=16'hf8;
17'h13368:	data_out=16'h8001;
17'h13369:	data_out=16'h67;
17'h1336a:	data_out=16'h8013;
17'h1336b:	data_out=16'h1f7;
17'h1336c:	data_out=16'h30c;
17'h1336d:	data_out=16'h72;
17'h1336e:	data_out=16'h8023;
17'h1336f:	data_out=16'h55;
17'h13370:	data_out=16'h8000;
17'h13371:	data_out=16'h804c;
17'h13372:	data_out=16'h106;
17'h13373:	data_out=16'h21b;
17'h13374:	data_out=16'h8d;
17'h13375:	data_out=16'h829c;
17'h13376:	data_out=16'h2bc;
17'h13377:	data_out=16'h1e6;
17'h13378:	data_out=16'h8055;
17'h13379:	data_out=16'h80ca;
17'h1337a:	data_out=16'h10;
17'h1337b:	data_out=16'he;
17'h1337c:	data_out=16'h4d;
17'h1337d:	data_out=16'h80d2;
17'h1337e:	data_out=16'h3bd;
17'h1337f:	data_out=16'h124;
17'h13380:	data_out=16'h9;
17'h13381:	data_out=16'h8002;
17'h13382:	data_out=16'h11;
17'h13383:	data_out=16'he;
17'h13384:	data_out=16'ha;
17'h13385:	data_out=16'h5;
17'h13386:	data_out=16'h1;
17'h13387:	data_out=16'h6;
17'h13388:	data_out=16'h2;
17'h13389:	data_out=16'h8002;
17'h1338a:	data_out=16'h14;
17'h1338b:	data_out=16'h7;
17'h1338c:	data_out=16'h2;
17'h1338d:	data_out=16'h8002;
17'h1338e:	data_out=16'h6;
17'h1338f:	data_out=16'h8002;
17'h13390:	data_out=16'hf;
17'h13391:	data_out=16'h5;
17'h13392:	data_out=16'h13;
17'h13393:	data_out=16'h3;
17'h13394:	data_out=16'hc;
17'h13395:	data_out=16'h7;
17'h13396:	data_out=16'h2;
17'h13397:	data_out=16'h12;
17'h13398:	data_out=16'h5;
17'h13399:	data_out=16'h1;
17'h1339a:	data_out=16'h2;
17'h1339b:	data_out=16'h8;
17'h1339c:	data_out=16'h4;
17'h1339d:	data_out=16'h10;
17'h1339e:	data_out=16'he;
17'h1339f:	data_out=16'h8000;
17'h133a0:	data_out=16'he;
17'h133a1:	data_out=16'h3;
17'h133a2:	data_out=16'hf;
17'h133a3:	data_out=16'h6;
17'h133a4:	data_out=16'hc;
17'h133a5:	data_out=16'h5;
17'h133a6:	data_out=16'h11;
17'h133a7:	data_out=16'h14;
17'h133a8:	data_out=16'h8004;
17'h133a9:	data_out=16'he;
17'h133aa:	data_out=16'hc;
17'h133ab:	data_out=16'h8000;
17'h133ac:	data_out=16'hd;
17'h133ad:	data_out=16'h1;
17'h133ae:	data_out=16'ha;
17'h133af:	data_out=16'ha;
17'h133b0:	data_out=16'hc;
17'h133b1:	data_out=16'h8004;
17'h133b2:	data_out=16'hd;
17'h133b3:	data_out=16'h5;
17'h133b4:	data_out=16'hd;
17'h133b5:	data_out=16'h8001;
17'h133b6:	data_out=16'hf;
17'h133b7:	data_out=16'ha;
17'h133b8:	data_out=16'h8005;
17'h133b9:	data_out=16'h3;
17'h133ba:	data_out=16'h14;
17'h133bb:	data_out=16'hb;
17'h133bc:	data_out=16'ha;
17'h133bd:	data_out=16'h7;
17'h133be:	data_out=16'ha;
17'h133bf:	data_out=16'hd;
17'h133c0:	data_out=16'h2;
17'h133c1:	data_out=16'hd;
17'h133c2:	data_out=16'he;
17'h133c3:	data_out=16'h8004;
17'h133c4:	data_out=16'he;
17'h133c5:	data_out=16'h1;
17'h133c6:	data_out=16'h1;
17'h133c7:	data_out=16'h12;
17'h133c8:	data_out=16'h6;
17'h133c9:	data_out=16'hc;
17'h133ca:	data_out=16'h8;
17'h133cb:	data_out=16'h0;
17'h133cc:	data_out=16'hf;
17'h133cd:	data_out=16'h7;
17'h133ce:	data_out=16'he;
17'h133cf:	data_out=16'ha;
17'h133d0:	data_out=16'h9;
17'h133d1:	data_out=16'h7;
17'h133d2:	data_out=16'h6;
17'h133d3:	data_out=16'h9;
17'h133d4:	data_out=16'h8;
17'h133d5:	data_out=16'hf;
17'h133d6:	data_out=16'h15;
17'h133d7:	data_out=16'h16;
17'h133d8:	data_out=16'h18;
17'h133d9:	data_out=16'hf;
17'h133da:	data_out=16'hf;
17'h133db:	data_out=16'h9;
17'h133dc:	data_out=16'h8001;
17'h133dd:	data_out=16'hc;
17'h133de:	data_out=16'h10;
17'h133df:	data_out=16'h0;
17'h133e0:	data_out=16'h8;
17'h133e1:	data_out=16'h5;
17'h133e2:	data_out=16'h5;
17'h133e3:	data_out=16'h5;
17'h133e4:	data_out=16'h11;
17'h133e5:	data_out=16'h8;
17'h133e6:	data_out=16'h8001;
17'h133e7:	data_out=16'h1;
17'h133e8:	data_out=16'h9;
17'h133e9:	data_out=16'hc;
17'h133ea:	data_out=16'h8006;
17'h133eb:	data_out=16'h6;
17'h133ec:	data_out=16'h19;
17'h133ed:	data_out=16'h10;
17'h133ee:	data_out=16'h8007;
17'h133ef:	data_out=16'h6;
17'h133f0:	data_out=16'h8001;
17'h133f1:	data_out=16'hf;
17'h133f2:	data_out=16'hf;
17'h133f3:	data_out=16'h10;
17'h133f4:	data_out=16'h3;
17'h133f5:	data_out=16'h3;
17'h133f6:	data_out=16'he;
17'h133f7:	data_out=16'h3;
17'h133f8:	data_out=16'hb;
17'h133f9:	data_out=16'h12;
17'h133fa:	data_out=16'h5;
17'h133fb:	data_out=16'h8005;
17'h133fc:	data_out=16'h1;
17'h133fd:	data_out=16'hb;
17'h133fe:	data_out=16'h6;
17'h133ff:	data_out=16'h13;
17'h13400:	data_out=16'h3;
17'h13401:	data_out=16'h6;
17'h13402:	data_out=16'h8001;
17'h13403:	data_out=16'h3;
17'h13404:	data_out=16'hf;
17'h13405:	data_out=16'h0;
17'h13406:	data_out=16'h8000;
17'h13407:	data_out=16'hf;
17'h13408:	data_out=16'h7;
17'h13409:	data_out=16'h3;
17'h1340a:	data_out=16'h5;
17'h1340b:	data_out=16'h5;
17'h1340c:	data_out=16'h2;
17'h1340d:	data_out=16'h7;
17'h1340e:	data_out=16'h6;
17'h1340f:	data_out=16'h6;
17'h13410:	data_out=16'h8001;
17'h13411:	data_out=16'h5;
17'h13412:	data_out=16'h7;
17'h13413:	data_out=16'h3;
17'h13414:	data_out=16'hf;
17'h13415:	data_out=16'h1;
17'h13416:	data_out=16'h6;
17'h13417:	data_out=16'hf;
17'h13418:	data_out=16'h8003;
17'h13419:	data_out=16'h2;
17'h1341a:	data_out=16'h10;
17'h1341b:	data_out=16'h6;
17'h1341c:	data_out=16'h7;
17'h1341d:	data_out=16'h3;
17'h1341e:	data_out=16'h4;
17'h1341f:	data_out=16'h10;
17'h13420:	data_out=16'he;
17'h13421:	data_out=16'h8001;
17'h13422:	data_out=16'h1;
17'h13423:	data_out=16'h9;
17'h13424:	data_out=16'h3;
17'h13425:	data_out=16'h7;
17'h13426:	data_out=16'hc;
17'h13427:	data_out=16'h8000;
17'h13428:	data_out=16'h8;
17'h13429:	data_out=16'h1;
17'h1342a:	data_out=16'h8;
17'h1342b:	data_out=16'hd;
17'h1342c:	data_out=16'hb;
17'h1342d:	data_out=16'h8001;
17'h1342e:	data_out=16'ha;
17'h1342f:	data_out=16'hc;
17'h13430:	data_out=16'h8;
17'h13431:	data_out=16'hc;
17'h13432:	data_out=16'h8000;
17'h13433:	data_out=16'h7;
17'h13434:	data_out=16'h1;
17'h13435:	data_out=16'hc;
17'h13436:	data_out=16'h4;
17'h13437:	data_out=16'h4;
17'h13438:	data_out=16'h8006;
17'h13439:	data_out=16'h3;
17'h1343a:	data_out=16'he;
17'h1343b:	data_out=16'hb;
17'h1343c:	data_out=16'ha;
17'h1343d:	data_out=16'h1;
17'h1343e:	data_out=16'h6;
17'h1343f:	data_out=16'h7;
17'h13440:	data_out=16'h9;
17'h13441:	data_out=16'h10;
17'h13442:	data_out=16'h8;
17'h13443:	data_out=16'h8003;
17'h13444:	data_out=16'h8;
17'h13445:	data_out=16'h0;
17'h13446:	data_out=16'h8003;
17'h13447:	data_out=16'h5;
17'h13448:	data_out=16'h8;
17'h13449:	data_out=16'h8;
17'h1344a:	data_out=16'h6;
17'h1344b:	data_out=16'h4;
17'h1344c:	data_out=16'hc;
17'h1344d:	data_out=16'hb;
17'h1344e:	data_out=16'h8000;
17'h1344f:	data_out=16'h4;
17'h13450:	data_out=16'hd;
17'h13451:	data_out=16'h8001;
17'h13452:	data_out=16'h5;
17'h13453:	data_out=16'h8000;
17'h13454:	data_out=16'ha;
17'h13455:	data_out=16'h8000;
17'h13456:	data_out=16'h6;
17'h13457:	data_out=16'he;
17'h13458:	data_out=16'h6;
17'h13459:	data_out=16'h3;
17'h1345a:	data_out=16'h9;
17'h1345b:	data_out=16'h8005;
17'h1345c:	data_out=16'h4;
17'h1345d:	data_out=16'h5;
17'h1345e:	data_out=16'h9;
17'h1345f:	data_out=16'hd;
17'h13460:	data_out=16'h5;
17'h13461:	data_out=16'h8001;
17'h13462:	data_out=16'h8003;
17'h13463:	data_out=16'he;
17'h13464:	data_out=16'h3;
17'h13465:	data_out=16'h1;
17'h13466:	data_out=16'h8003;
17'h13467:	data_out=16'he;
17'h13468:	data_out=16'h6;
17'h13469:	data_out=16'h6;
17'h1346a:	data_out=16'h8007;
17'h1346b:	data_out=16'h5;
17'h1346c:	data_out=16'h3;
17'h1346d:	data_out=16'h8001;
17'h1346e:	data_out=16'h4;
17'h1346f:	data_out=16'hd;
17'h13470:	data_out=16'h8004;
17'h13471:	data_out=16'h6;
17'h13472:	data_out=16'h8002;
17'h13473:	data_out=16'hd;
17'h13474:	data_out=16'h5;
17'h13475:	data_out=16'h3;
17'h13476:	data_out=16'hc;
17'h13477:	data_out=16'hf;
17'h13478:	data_out=16'h8;
17'h13479:	data_out=16'hb;
17'h1347a:	data_out=16'he;
17'h1347b:	data_out=16'h8005;
17'h1347c:	data_out=16'hb;
17'h1347d:	data_out=16'h4;
17'h1347e:	data_out=16'h8001;
17'h1347f:	data_out=16'h5;
17'h13480:	data_out=16'h2;
17'h13481:	data_out=16'h8001;
17'h13482:	data_out=16'h4;
17'h13483:	data_out=16'h11;
17'h13484:	data_out=16'h7;
17'h13485:	data_out=16'h5;
17'h13486:	data_out=16'hb;
17'h13487:	data_out=16'h3;
17'h13488:	data_out=16'ha;
17'h13489:	data_out=16'ha;
17'h1348a:	data_out=16'h9;
17'h1348b:	data_out=16'hf;
17'h1348c:	data_out=16'h12;
17'h1348d:	data_out=16'h3;
17'h1348e:	data_out=16'h9;
17'h1348f:	data_out=16'h12;
17'h13490:	data_out=16'h9;
17'h13491:	data_out=16'hf;
17'h13492:	data_out=16'h15;
17'h13493:	data_out=16'h12;
17'h13494:	data_out=16'h8;
17'h13495:	data_out=16'ha;
17'h13496:	data_out=16'hb;
17'h13497:	data_out=16'h15;
17'h13498:	data_out=16'h4;
17'h13499:	data_out=16'h5;
17'h1349a:	data_out=16'h4;
17'h1349b:	data_out=16'h5;
17'h1349c:	data_out=16'hf;
17'h1349d:	data_out=16'h3;
17'h1349e:	data_out=16'ha;
17'h1349f:	data_out=16'ha;
17'h134a0:	data_out=16'h4;
17'h134a1:	data_out=16'h6;
17'h134a2:	data_out=16'h6;
17'h134a3:	data_out=16'h6;
17'h134a4:	data_out=16'h9;
17'h134a5:	data_out=16'h2;
17'h134a6:	data_out=16'hc;
17'h134a7:	data_out=16'h7;
17'h134a8:	data_out=16'ha;
17'h134a9:	data_out=16'h5;
17'h134aa:	data_out=16'h9;
17'h134ab:	data_out=16'h9;
17'h134ac:	data_out=16'h7;
17'h134ad:	data_out=16'h1;
17'h134ae:	data_out=16'h13;
17'h134af:	data_out=16'hf;
17'h134b0:	data_out=16'h15;
17'h134b1:	data_out=16'h7;
17'h134b2:	data_out=16'h11;
17'h134b3:	data_out=16'h5;
17'h134b4:	data_out=16'h5;
17'h134b5:	data_out=16'hc;
17'h134b6:	data_out=16'h1;
17'h134b7:	data_out=16'he;
17'h134b8:	data_out=16'ha;
17'h134b9:	data_out=16'h2;
17'h134ba:	data_out=16'hf;
17'h134bb:	data_out=16'hd;
17'h134bc:	data_out=16'h8;
17'h134bd:	data_out=16'h3;
17'h134be:	data_out=16'h1;
17'h134bf:	data_out=16'hf;
17'h134c0:	data_out=16'h14;
17'h134c1:	data_out=16'he;
17'h134c2:	data_out=16'h9;
17'h134c3:	data_out=16'he;
17'h134c4:	data_out=16'h11;
17'h134c5:	data_out=16'h8001;
17'h134c6:	data_out=16'h2;
17'h134c7:	data_out=16'hd;
17'h134c8:	data_out=16'hc;
17'h134c9:	data_out=16'hc;
17'h134ca:	data_out=16'hc;
17'h134cb:	data_out=16'h13;
17'h134cc:	data_out=16'h12;
17'h134cd:	data_out=16'hf;
17'h134ce:	data_out=16'h10;
17'h134cf:	data_out=16'h10;
17'h134d0:	data_out=16'hb;
17'h134d1:	data_out=16'h5;
17'h134d2:	data_out=16'h6;
17'h134d3:	data_out=16'h10;
17'h134d4:	data_out=16'hd;
17'h134d5:	data_out=16'h11;
17'h134d6:	data_out=16'hc;
17'h134d7:	data_out=16'hb;
17'h134d8:	data_out=16'h14;
17'h134d9:	data_out=16'h7;
17'h134da:	data_out=16'h9;
17'h134db:	data_out=16'h3;
17'h134dc:	data_out=16'hc;
17'h134dd:	data_out=16'h10;
17'h134de:	data_out=16'h2;
17'h134df:	data_out=16'ha;
17'h134e0:	data_out=16'hc;
17'h134e1:	data_out=16'h8;
17'h134e2:	data_out=16'h7;
17'h134e3:	data_out=16'h9;
17'h134e4:	data_out=16'ha;
17'h134e5:	data_out=16'h11;
17'h134e6:	data_out=16'h11;
17'h134e7:	data_out=16'h15;
17'h134e8:	data_out=16'h1;
17'h134e9:	data_out=16'h7;
17'h134ea:	data_out=16'h8;
17'h134eb:	data_out=16'h1;
17'h134ec:	data_out=16'h3;
17'h134ed:	data_out=16'ha;
17'h134ee:	data_out=16'h6;
17'h134ef:	data_out=16'he;
17'h134f0:	data_out=16'h8;
17'h134f1:	data_out=16'hb;
17'h134f2:	data_out=16'h10;
17'h134f3:	data_out=16'h9;
17'h134f4:	data_out=16'h7;
17'h134f5:	data_out=16'h2;
17'h134f6:	data_out=16'h8001;
17'h134f7:	data_out=16'h6;
17'h134f8:	data_out=16'h6;
17'h134f9:	data_out=16'h12;
17'h134fa:	data_out=16'hd;
17'h134fb:	data_out=16'h8003;
17'h134fc:	data_out=16'h2;
17'h134fd:	data_out=16'h9;
17'h134fe:	data_out=16'hc;
17'h134ff:	data_out=16'h13;
17'h13500:	data_out=16'h857c;
17'h13501:	data_out=16'h1cb;
17'h13502:	data_out=16'h9b;
17'h13503:	data_out=16'h15c;
17'h13504:	data_out=16'h2c0;
17'h13505:	data_out=16'h720;
17'h13506:	data_out=16'h56f;
17'h13507:	data_out=16'h2a3;
17'h13508:	data_out=16'h57;
17'h13509:	data_out=16'h800c;
17'h1350a:	data_out=16'h98;
17'h1350b:	data_out=16'h5b2;
17'h1350c:	data_out=16'h597;
17'h1350d:	data_out=16'h3c;
17'h1350e:	data_out=16'h10b;
17'h1350f:	data_out=16'h259;
17'h13510:	data_out=16'h8023;
17'h13511:	data_out=16'h538;
17'h13512:	data_out=16'h18d;
17'h13513:	data_out=16'h221;
17'h13514:	data_out=16'h30f;
17'h13515:	data_out=16'h8084;
17'h13516:	data_out=16'h806e;
17'h13517:	data_out=16'h321;
17'h13518:	data_out=16'h8012;
17'h13519:	data_out=16'h425;
17'h1351a:	data_out=16'h362;
17'h1351b:	data_out=16'h5a4;
17'h1351c:	data_out=16'h4f8;
17'h1351d:	data_out=16'h3bb;
17'h1351e:	data_out=16'h2c2;
17'h1351f:	data_out=16'h347;
17'h13520:	data_out=16'h52d;
17'h13521:	data_out=16'h128;
17'h13522:	data_out=16'hae;
17'h13523:	data_out=16'h81ee;
17'h13524:	data_out=16'h81ef;
17'h13525:	data_out=16'h1d9;
17'h13526:	data_out=16'h8083;
17'h13527:	data_out=16'h47d;
17'h13528:	data_out=16'h157;
17'h13529:	data_out=16'h8204;
17'h1352a:	data_out=16'h8051;
17'h1352b:	data_out=16'h7f1;
17'h1352c:	data_out=16'h8059;
17'h1352d:	data_out=16'h845d;
17'h1352e:	data_out=16'h1fe;
17'h1352f:	data_out=16'h4d7;
17'h13530:	data_out=16'h41b;
17'h13531:	data_out=16'h38e;
17'h13532:	data_out=16'h435;
17'h13533:	data_out=16'h31e;
17'h13534:	data_out=16'h28f;
17'h13535:	data_out=16'h8b8;
17'h13536:	data_out=16'h12e;
17'h13537:	data_out=16'h176;
17'h13538:	data_out=16'h4a2;
17'h13539:	data_out=16'h2f8;
17'h1353a:	data_out=16'h828e;
17'h1353b:	data_out=16'h317;
17'h1353c:	data_out=16'h222;
17'h1353d:	data_out=16'h31c;
17'h1353e:	data_out=16'h159;
17'h1353f:	data_out=16'h71f;
17'h13540:	data_out=16'h223;
17'h13541:	data_out=16'h3e1;
17'h13542:	data_out=16'h8240;
17'h13543:	data_out=16'h438;
17'h13544:	data_out=16'h309;
17'h13545:	data_out=16'h80a2;
17'h13546:	data_out=16'h205;
17'h13547:	data_out=16'h8132;
17'h13548:	data_out=16'h3aa;
17'h13549:	data_out=16'h214;
17'h1354a:	data_out=16'h283;
17'h1354b:	data_out=16'h1bd;
17'h1354c:	data_out=16'h9;
17'h1354d:	data_out=16'ha2;
17'h1354e:	data_out=16'h1af;
17'h1354f:	data_out=16'h28;
17'h13550:	data_out=16'h805e;
17'h13551:	data_out=16'h3a8;
17'h13552:	data_out=16'h82e4;
17'h13553:	data_out=16'h67f;
17'h13554:	data_out=16'h3ec;
17'h13555:	data_out=16'h2d3;
17'h13556:	data_out=16'h43;
17'h13557:	data_out=16'h80df;
17'h13558:	data_out=16'h75;
17'h13559:	data_out=16'hf6;
17'h1355a:	data_out=16'h406;
17'h1355b:	data_out=16'h4c9;
17'h1355c:	data_out=16'h59a;
17'h1355d:	data_out=16'h8003;
17'h1355e:	data_out=16'h4b0;
17'h1355f:	data_out=16'h8019;
17'h13560:	data_out=16'h812d;
17'h13561:	data_out=16'h4fc;
17'h13562:	data_out=16'h2e7;
17'h13563:	data_out=16'h36e;
17'h13564:	data_out=16'h3d4;
17'h13565:	data_out=16'h50c;
17'h13566:	data_out=16'h6ce;
17'h13567:	data_out=16'h192;
17'h13568:	data_out=16'h13e;
17'h13569:	data_out=16'h3d;
17'h1356a:	data_out=16'hf4;
17'h1356b:	data_out=16'h48a;
17'h1356c:	data_out=16'h8902;
17'h1356d:	data_out=16'h355;
17'h1356e:	data_out=16'he7;
17'h1356f:	data_out=16'h37b;
17'h13570:	data_out=16'hfa;
17'h13571:	data_out=16'h244;
17'h13572:	data_out=16'h32b;
17'h13573:	data_out=16'h528;
17'h13574:	data_out=16'h41a;
17'h13575:	data_out=16'h4d0;
17'h13576:	data_out=16'h63c;
17'h13577:	data_out=16'h39;
17'h13578:	data_out=16'h40b;
17'h13579:	data_out=16'h1e6;
17'h1357a:	data_out=16'h385;
17'h1357b:	data_out=16'h159;
17'h1357c:	data_out=16'h1b;
17'h1357d:	data_out=16'h60f;
17'h1357e:	data_out=16'h1b4;
17'h1357f:	data_out=16'h8060;
17'h13580:	data_out=16'h89fc;
17'h13581:	data_out=16'h5f5;
17'h13582:	data_out=16'h967;
17'h13583:	data_out=16'h9ec;
17'h13584:	data_out=16'ha00;
17'h13585:	data_out=16'ha00;
17'h13586:	data_out=16'h9fe;
17'h13587:	data_out=16'h772;
17'h13588:	data_out=16'h83c4;
17'h13589:	data_out=16'h4d6;
17'h1358a:	data_out=16'h81d3;
17'h1358b:	data_out=16'h9fa;
17'h1358c:	data_out=16'h6eb;
17'h1358d:	data_out=16'h862;
17'h1358e:	data_out=16'h336;
17'h1358f:	data_out=16'h9f3;
17'h13590:	data_out=16'h7af;
17'h13591:	data_out=16'ha00;
17'h13592:	data_out=16'h9fc;
17'h13593:	data_out=16'h9ff;
17'h13594:	data_out=16'ha00;
17'h13595:	data_out=16'h459;
17'h13596:	data_out=16'h3db;
17'h13597:	data_out=16'h9fb;
17'h13598:	data_out=16'h10a;
17'h13599:	data_out=16'h9ff;
17'h1359a:	data_out=16'ha00;
17'h1359b:	data_out=16'h9fa;
17'h1359c:	data_out=16'h9fe;
17'h1359d:	data_out=16'h9ff;
17'h1359e:	data_out=16'h9fd;
17'h1359f:	data_out=16'ha00;
17'h135a0:	data_out=16'ha00;
17'h135a1:	data_out=16'h357;
17'h135a2:	data_out=16'h9f7;
17'h135a3:	data_out=16'h884a;
17'h135a4:	data_out=16'h884c;
17'h135a5:	data_out=16'h7af;
17'h135a6:	data_out=16'h86e7;
17'h135a7:	data_out=16'ha00;
17'h135a8:	data_out=16'h3c2;
17'h135a9:	data_out=16'h405;
17'h135aa:	data_out=16'h8073;
17'h135ab:	data_out=16'ha00;
17'h135ac:	data_out=16'h536;
17'h135ad:	data_out=16'h8a00;
17'h135ae:	data_out=16'h9f7;
17'h135af:	data_out=16'ha00;
17'h135b0:	data_out=16'h6cd;
17'h135b1:	data_out=16'ha00;
17'h135b2:	data_out=16'h7eb;
17'h135b3:	data_out=16'ha00;
17'h135b4:	data_out=16'h5fe;
17'h135b5:	data_out=16'ha00;
17'h135b6:	data_out=16'h3e9;
17'h135b7:	data_out=16'h97c;
17'h135b8:	data_out=16'h9ff;
17'h135b9:	data_out=16'ha00;
17'h135ba:	data_out=16'h8085;
17'h135bb:	data_out=16'h8b2;
17'h135bc:	data_out=16'h6be;
17'h135bd:	data_out=16'ha00;
17'h135be:	data_out=16'h3c7;
17'h135bf:	data_out=16'ha00;
17'h135c0:	data_out=16'ha00;
17'h135c1:	data_out=16'h9fa;
17'h135c2:	data_out=16'h89fe;
17'h135c3:	data_out=16'ha00;
17'h135c4:	data_out=16'ha00;
17'h135c5:	data_out=16'h477;
17'h135c6:	data_out=16'h8138;
17'h135c7:	data_out=16'h17b;
17'h135c8:	data_out=16'h9ff;
17'h135c9:	data_out=16'h948;
17'h135ca:	data_out=16'h95a;
17'h135cb:	data_out=16'h89e2;
17'h135cc:	data_out=16'h822f;
17'h135cd:	data_out=16'h9f8;
17'h135ce:	data_out=16'h910;
17'h135cf:	data_out=16'h80e9;
17'h135d0:	data_out=16'h9fc;
17'h135d1:	data_out=16'h9fd;
17'h135d2:	data_out=16'h89fb;
17'h135d3:	data_out=16'h9ff;
17'h135d4:	data_out=16'ha00;
17'h135d5:	data_out=16'h9f8;
17'h135d6:	data_out=16'h9de;
17'h135d7:	data_out=16'ha00;
17'h135d8:	data_out=16'h8c8;
17'h135d9:	data_out=16'ha00;
17'h135da:	data_out=16'h9fb;
17'h135db:	data_out=16'ha00;
17'h135dc:	data_out=16'h9ff;
17'h135dd:	data_out=16'h44f;
17'h135de:	data_out=16'ha00;
17'h135df:	data_out=16'h9;
17'h135e0:	data_out=16'h89fb;
17'h135e1:	data_out=16'ha00;
17'h135e2:	data_out=16'h9f7;
17'h135e3:	data_out=16'ha00;
17'h135e4:	data_out=16'h94d;
17'h135e5:	data_out=16'ha00;
17'h135e6:	data_out=16'ha00;
17'h135e7:	data_out=16'h9fb;
17'h135e8:	data_out=16'h37a;
17'h135e9:	data_out=16'h85d6;
17'h135ea:	data_out=16'h322;
17'h135eb:	data_out=16'ha00;
17'h135ec:	data_out=16'h89fc;
17'h135ed:	data_out=16'ha00;
17'h135ee:	data_out=16'h322;
17'h135ef:	data_out=16'ha00;
17'h135f0:	data_out=16'h32c;
17'h135f1:	data_out=16'h9fa;
17'h135f2:	data_out=16'ha00;
17'h135f3:	data_out=16'ha00;
17'h135f4:	data_out=16'h663;
17'h135f5:	data_out=16'h9ff;
17'h135f6:	data_out=16'ha00;
17'h135f7:	data_out=16'h9f0;
17'h135f8:	data_out=16'h9ff;
17'h135f9:	data_out=16'h938;
17'h135fa:	data_out=16'ha00;
17'h135fb:	data_out=16'h3c8;
17'h135fc:	data_out=16'h197;
17'h135fd:	data_out=16'ha00;
17'h135fe:	data_out=16'h9ff;
17'h135ff:	data_out=16'ha00;
17'h13600:	data_out=16'h8468;
17'h13601:	data_out=16'ha00;
17'h13602:	data_out=16'h9b9;
17'h13603:	data_out=16'h611;
17'h13604:	data_out=16'ha00;
17'h13605:	data_out=16'ha00;
17'h13606:	data_out=16'h6cb;
17'h13607:	data_out=16'h8a00;
17'h13608:	data_out=16'h8333;
17'h13609:	data_out=16'h8a00;
17'h1360a:	data_out=16'h1b9;
17'h1360b:	data_out=16'h85fe;
17'h1360c:	data_out=16'h8a00;
17'h1360d:	data_out=16'h581;
17'h1360e:	data_out=16'h57d;
17'h1360f:	data_out=16'h8ac;
17'h13610:	data_out=16'h81d9;
17'h13611:	data_out=16'ha00;
17'h13612:	data_out=16'h810b;
17'h13613:	data_out=16'ha00;
17'h13614:	data_out=16'h9f3;
17'h13615:	data_out=16'ha00;
17'h13616:	data_out=16'h9be;
17'h13617:	data_out=16'h793;
17'h13618:	data_out=16'h275;
17'h13619:	data_out=16'h9fb;
17'h1361a:	data_out=16'ha00;
17'h1361b:	data_out=16'h957;
17'h1361c:	data_out=16'h9fd;
17'h1361d:	data_out=16'h9f3;
17'h1361e:	data_out=16'h9fb;
17'h1361f:	data_out=16'h9f5;
17'h13620:	data_out=16'ha00;
17'h13621:	data_out=16'h5b4;
17'h13622:	data_out=16'h8519;
17'h13623:	data_out=16'h89ff;
17'h13624:	data_out=16'h89ff;
17'h13625:	data_out=16'h89ff;
17'h13626:	data_out=16'h89ff;
17'h13627:	data_out=16'ha00;
17'h13628:	data_out=16'h673;
17'h13629:	data_out=16'h11f;
17'h1362a:	data_out=16'h8a00;
17'h1362b:	data_out=16'ha00;
17'h1362c:	data_out=16'h9ff;
17'h1362d:	data_out=16'h8a00;
17'h1362e:	data_out=16'h195;
17'h1362f:	data_out=16'ha00;
17'h13630:	data_out=16'h79d;
17'h13631:	data_out=16'ha00;
17'h13632:	data_out=16'h90c;
17'h13633:	data_out=16'h9f9;
17'h13634:	data_out=16'h29f;
17'h13635:	data_out=16'h9ff;
17'h13636:	data_out=16'h902;
17'h13637:	data_out=16'h8b6;
17'h13638:	data_out=16'h9fb;
17'h13639:	data_out=16'h9fd;
17'h1363a:	data_out=16'h89f1;
17'h1363b:	data_out=16'h90b;
17'h1363c:	data_out=16'h9fd;
17'h1363d:	data_out=16'ha00;
17'h1363e:	data_out=16'h67b;
17'h1363f:	data_out=16'ha00;
17'h13640:	data_out=16'h82c;
17'h13641:	data_out=16'h9f1;
17'h13642:	data_out=16'h8a00;
17'h13643:	data_out=16'h9f8;
17'h13644:	data_out=16'ha00;
17'h13645:	data_out=16'ha00;
17'h13646:	data_out=16'h853a;
17'h13647:	data_out=16'h89ff;
17'h13648:	data_out=16'h76c;
17'h13649:	data_out=16'h89f8;
17'h1364a:	data_out=16'h81b2;
17'h1364b:	data_out=16'h8a00;
17'h1364c:	data_out=16'h8a00;
17'h1364d:	data_out=16'h811a;
17'h1364e:	data_out=16'h80db;
17'h1364f:	data_out=16'h8a00;
17'h13650:	data_out=16'h9f5;
17'h13651:	data_out=16'h99c;
17'h13652:	data_out=16'h89f8;
17'h13653:	data_out=16'ha00;
17'h13654:	data_out=16'ha00;
17'h13655:	data_out=16'h67f;
17'h13656:	data_out=16'h8;
17'h13657:	data_out=16'h816f;
17'h13658:	data_out=16'h9f9;
17'h13659:	data_out=16'h5a9;
17'h1365a:	data_out=16'h863;
17'h1365b:	data_out=16'ha00;
17'h1365c:	data_out=16'h9d0;
17'h1365d:	data_out=16'h558;
17'h1365e:	data_out=16'ha00;
17'h1365f:	data_out=16'h24b;
17'h13660:	data_out=16'h8a00;
17'h13661:	data_out=16'h9fe;
17'h13662:	data_out=16'h548;
17'h13663:	data_out=16'h9f5;
17'h13664:	data_out=16'h307;
17'h13665:	data_out=16'h64b;
17'h13666:	data_out=16'h9fe;
17'h13667:	data_out=16'h9f3;
17'h13668:	data_out=16'h5ec;
17'h13669:	data_out=16'h896d;
17'h1366a:	data_out=16'h559;
17'h1366b:	data_out=16'ha00;
17'h1366c:	data_out=16'h8848;
17'h1366d:	data_out=16'h9f7;
17'h1366e:	data_out=16'h559;
17'h1366f:	data_out=16'h99f;
17'h13670:	data_out=16'h56c;
17'h13671:	data_out=16'h9e4;
17'h13672:	data_out=16'ha00;
17'h13673:	data_out=16'ha00;
17'h13674:	data_out=16'h682;
17'h13675:	data_out=16'h807;
17'h13676:	data_out=16'h9fe;
17'h13677:	data_out=16'h63b;
17'h13678:	data_out=16'h9a2;
17'h13679:	data_out=16'h1b3;
17'h1367a:	data_out=16'h9f5;
17'h1367b:	data_out=16'h67c;
17'h1367c:	data_out=16'h730;
17'h1367d:	data_out=16'ha00;
17'h1367e:	data_out=16'h86a2;
17'h1367f:	data_out=16'ha00;
17'h13680:	data_out=16'ha00;
17'h13681:	data_out=16'ha00;
17'h13682:	data_out=16'h870a;
17'h13683:	data_out=16'h63a;
17'h13684:	data_out=16'h9f9;
17'h13685:	data_out=16'h9f3;
17'h13686:	data_out=16'h5e9;
17'h13687:	data_out=16'h8a00;
17'h13688:	data_out=16'h8942;
17'h13689:	data_out=16'h8a00;
17'h1368a:	data_out=16'h9f6;
17'h1368b:	data_out=16'h89e9;
17'h1368c:	data_out=16'h8a00;
17'h1368d:	data_out=16'h89e7;
17'h1368e:	data_out=16'h26c;
17'h1368f:	data_out=16'h89f1;
17'h13690:	data_out=16'h89fe;
17'h13691:	data_out=16'ha00;
17'h13692:	data_out=16'hea;
17'h13693:	data_out=16'ha00;
17'h13694:	data_out=16'h9f4;
17'h13695:	data_out=16'ha00;
17'h13696:	data_out=16'h9c5;
17'h13697:	data_out=16'h9f1;
17'h13698:	data_out=16'h89dd;
17'h13699:	data_out=16'h9fb;
17'h1369a:	data_out=16'h9ef;
17'h1369b:	data_out=16'h41c;
17'h1369c:	data_out=16'ha00;
17'h1369d:	data_out=16'ha00;
17'h1369e:	data_out=16'h9fc;
17'h1369f:	data_out=16'h4f9;
17'h136a0:	data_out=16'ha00;
17'h136a1:	data_out=16'h255;
17'h136a2:	data_out=16'h8a00;
17'h136a3:	data_out=16'h88b5;
17'h136a4:	data_out=16'h88b4;
17'h136a5:	data_out=16'h8a00;
17'h136a6:	data_out=16'h89ea;
17'h136a7:	data_out=16'ha00;
17'h136a8:	data_out=16'h2d9;
17'h136a9:	data_out=16'h99c;
17'h136aa:	data_out=16'h89e4;
17'h136ab:	data_out=16'ha00;
17'h136ac:	data_out=16'ha00;
17'h136ad:	data_out=16'h821f;
17'h136ae:	data_out=16'h8966;
17'h136af:	data_out=16'ha00;
17'h136b0:	data_out=16'h64f;
17'h136b1:	data_out=16'ha00;
17'h136b2:	data_out=16'h9d3;
17'h136b3:	data_out=16'h9f8;
17'h136b4:	data_out=16'ha00;
17'h136b5:	data_out=16'h9b1;
17'h136b6:	data_out=16'h88b6;
17'h136b7:	data_out=16'h83a6;
17'h136b8:	data_out=16'h9fb;
17'h136b9:	data_out=16'h9fc;
17'h136ba:	data_out=16'h8a00;
17'h136bb:	data_out=16'hfe;
17'h136bc:	data_out=16'ha00;
17'h136bd:	data_out=16'ha00;
17'h136be:	data_out=16'h2e4;
17'h136bf:	data_out=16'h9f3;
17'h136c0:	data_out=16'h874c;
17'h136c1:	data_out=16'h84e4;
17'h136c2:	data_out=16'h89ff;
17'h136c3:	data_out=16'h9f2;
17'h136c4:	data_out=16'ha00;
17'h136c5:	data_out=16'ha00;
17'h136c6:	data_out=16'h3fb;
17'h136c7:	data_out=16'h89f5;
17'h136c8:	data_out=16'h874f;
17'h136c9:	data_out=16'h8a00;
17'h136ca:	data_out=16'h88cb;
17'h136cb:	data_out=16'h8a00;
17'h136cc:	data_out=16'h8a00;
17'h136cd:	data_out=16'h8a00;
17'h136ce:	data_out=16'h8872;
17'h136cf:	data_out=16'h8a00;
17'h136d0:	data_out=16'h8377;
17'h136d1:	data_out=16'h5c5;
17'h136d2:	data_out=16'h89fe;
17'h136d3:	data_out=16'ha00;
17'h136d4:	data_out=16'ha00;
17'h136d5:	data_out=16'h370;
17'h136d6:	data_out=16'h89ed;
17'h136d7:	data_out=16'h87d5;
17'h136d8:	data_out=16'h65f;
17'h136d9:	data_out=16'h84bc;
17'h136da:	data_out=16'h838;
17'h136db:	data_out=16'ha00;
17'h136dc:	data_out=16'h9e2;
17'h136dd:	data_out=16'h1c5;
17'h136de:	data_out=16'ha00;
17'h136df:	data_out=16'h87e2;
17'h136e0:	data_out=16'h89ec;
17'h136e1:	data_out=16'h9fd;
17'h136e2:	data_out=16'h89b;
17'h136e3:	data_out=16'h9f6;
17'h136e4:	data_out=16'h6d0;
17'h136e5:	data_out=16'h8566;
17'h136e6:	data_out=16'h9f9;
17'h136e7:	data_out=16'h8140;
17'h136e8:	data_out=16'h266;
17'h136e9:	data_out=16'h89e9;
17'h136ea:	data_out=16'h275;
17'h136eb:	data_out=16'h9fd;
17'h136ec:	data_out=16'ha00;
17'h136ed:	data_out=16'h9f7;
17'h136ee:	data_out=16'h274;
17'h136ef:	data_out=16'h95d;
17'h136f0:	data_out=16'h271;
17'h136f1:	data_out=16'h83b9;
17'h136f2:	data_out=16'h9fc;
17'h136f3:	data_out=16'h9f1;
17'h136f4:	data_out=16'h5c5;
17'h136f5:	data_out=16'h8b6;
17'h136f6:	data_out=16'h9fe;
17'h136f7:	data_out=16'h8a00;
17'h136f8:	data_out=16'h9ec;
17'h136f9:	data_out=16'h89f9;
17'h136fa:	data_out=16'h9f6;
17'h136fb:	data_out=16'h2e6;
17'h136fc:	data_out=16'h87d9;
17'h136fd:	data_out=16'h9f2;
17'h136fe:	data_out=16'h8775;
17'h136ff:	data_out=16'h8381;
17'h13700:	data_out=16'ha00;
17'h13701:	data_out=16'ha00;
17'h13702:	data_out=16'h8a00;
17'h13703:	data_out=16'h89fc;
17'h13704:	data_out=16'h2e0;
17'h13705:	data_out=16'h9d7;
17'h13706:	data_out=16'h7dd;
17'h13707:	data_out=16'h8a00;
17'h13708:	data_out=16'h89cb;
17'h13709:	data_out=16'h8a00;
17'h1370a:	data_out=16'ha00;
17'h1370b:	data_out=16'h89c0;
17'h1370c:	data_out=16'h8a00;
17'h1370d:	data_out=16'h8a00;
17'h1370e:	data_out=16'h4f4;
17'h1370f:	data_out=16'h8a00;
17'h13710:	data_out=16'h8a00;
17'h13711:	data_out=16'ha00;
17'h13712:	data_out=16'h8073;
17'h13713:	data_out=16'h9fe;
17'h13714:	data_out=16'h518;
17'h13715:	data_out=16'h3bb;
17'h13716:	data_out=16'h85c7;
17'h13717:	data_out=16'h459;
17'h13718:	data_out=16'h89fb;
17'h13719:	data_out=16'h9f9;
17'h1371a:	data_out=16'h9d2;
17'h1371b:	data_out=16'h8882;
17'h1371c:	data_out=16'h9e3;
17'h1371d:	data_out=16'ha00;
17'h1371e:	data_out=16'h2f5;
17'h1371f:	data_out=16'h8840;
17'h13720:	data_out=16'ha00;
17'h13721:	data_out=16'h423;
17'h13722:	data_out=16'h8a00;
17'h13723:	data_out=16'h65e;
17'h13724:	data_out=16'h63d;
17'h13725:	data_out=16'h8a00;
17'h13726:	data_out=16'h89f9;
17'h13727:	data_out=16'h9ff;
17'h13728:	data_out=16'h415;
17'h13729:	data_out=16'h9d2;
17'h1372a:	data_out=16'h89ee;
17'h1372b:	data_out=16'ha00;
17'h1372c:	data_out=16'h291;
17'h1372d:	data_out=16'h9f3;
17'h1372e:	data_out=16'h899c;
17'h1372f:	data_out=16'ha00;
17'h13730:	data_out=16'h52f;
17'h13731:	data_out=16'ha00;
17'h13732:	data_out=16'h9c0;
17'h13733:	data_out=16'h8a4;
17'h13734:	data_out=16'ha00;
17'h13735:	data_out=16'h6ac;
17'h13736:	data_out=16'h89cb;
17'h13737:	data_out=16'h86e6;
17'h13738:	data_out=16'ha00;
17'h13739:	data_out=16'h799;
17'h1373a:	data_out=16'h8a00;
17'h1373b:	data_out=16'h828b;
17'h1373c:	data_out=16'ha00;
17'h1373d:	data_out=16'ha00;
17'h1373e:	data_out=16'h421;
17'h1373f:	data_out=16'h9d7;
17'h13740:	data_out=16'h89eb;
17'h13741:	data_out=16'h89fa;
17'h13742:	data_out=16'h8a00;
17'h13743:	data_out=16'h82bc;
17'h13744:	data_out=16'ha00;
17'h13745:	data_out=16'h385;
17'h13746:	data_out=16'h971;
17'h13747:	data_out=16'h8a00;
17'h13748:	data_out=16'h89ff;
17'h13749:	data_out=16'h8a00;
17'h1374a:	data_out=16'h8998;
17'h1374b:	data_out=16'h8a00;
17'h1374c:	data_out=16'h8a00;
17'h1374d:	data_out=16'h8a00;
17'h1374e:	data_out=16'h88cb;
17'h1374f:	data_out=16'h8a00;
17'h13750:	data_out=16'h89b1;
17'h13751:	data_out=16'h89fe;
17'h13752:	data_out=16'h8a00;
17'h13753:	data_out=16'ha00;
17'h13754:	data_out=16'ha00;
17'h13755:	data_out=16'h89ff;
17'h13756:	data_out=16'h89f7;
17'h13757:	data_out=16'h88b5;
17'h13758:	data_out=16'h89fd;
17'h13759:	data_out=16'h82e9;
17'h1375a:	data_out=16'h6bb;
17'h1375b:	data_out=16'ha00;
17'h1375c:	data_out=16'h9d9;
17'h1375d:	data_out=16'h882b;
17'h1375e:	data_out=16'ha00;
17'h1375f:	data_out=16'h895d;
17'h13760:	data_out=16'h89f7;
17'h13761:	data_out=16'h9f2;
17'h13762:	data_out=16'h3ba;
17'h13763:	data_out=16'h97d;
17'h13764:	data_out=16'ha00;
17'h13765:	data_out=16'h9f8;
17'h13766:	data_out=16'h7b4;
17'h13767:	data_out=16'h8780;
17'h13768:	data_out=16'h3da;
17'h13769:	data_out=16'h89f8;
17'h1376a:	data_out=16'h573;
17'h1376b:	data_out=16'h9d9;
17'h1376c:	data_out=16'ha00;
17'h1376d:	data_out=16'h98f;
17'h1376e:	data_out=16'h570;
17'h1376f:	data_out=16'h6f2;
17'h13770:	data_out=16'h530;
17'h13771:	data_out=16'h89f6;
17'h13772:	data_out=16'h9f0;
17'h13773:	data_out=16'h9f5;
17'h13774:	data_out=16'h4cf;
17'h13775:	data_out=16'h93d;
17'h13776:	data_out=16'h9fa;
17'h13777:	data_out=16'h8a00;
17'h13778:	data_out=16'h3a2;
17'h13779:	data_out=16'h8a00;
17'h1377a:	data_out=16'h782;
17'h1377b:	data_out=16'h423;
17'h1377c:	data_out=16'h89f7;
17'h1377d:	data_out=16'h8402;
17'h1377e:	data_out=16'ha0;
17'h1377f:	data_out=16'h899a;
17'h13780:	data_out=16'ha00;
17'h13781:	data_out=16'ha00;
17'h13782:	data_out=16'h86b6;
17'h13783:	data_out=16'h89dd;
17'h13784:	data_out=16'h8415;
17'h13785:	data_out=16'h89f;
17'h13786:	data_out=16'h769;
17'h13787:	data_out=16'h8a00;
17'h13788:	data_out=16'h8992;
17'h13789:	data_out=16'h8a00;
17'h1378a:	data_out=16'ha00;
17'h1378b:	data_out=16'h8801;
17'h1378c:	data_out=16'h8a00;
17'h1378d:	data_out=16'h8a00;
17'h1378e:	data_out=16'h9f5;
17'h1378f:	data_out=16'h8a00;
17'h13790:	data_out=16'h89fb;
17'h13791:	data_out=16'ha00;
17'h13792:	data_out=16'h8836;
17'h13793:	data_out=16'ha00;
17'h13794:	data_out=16'h829d;
17'h13795:	data_out=16'h8171;
17'h13796:	data_out=16'h89b8;
17'h13797:	data_out=16'h8383;
17'h13798:	data_out=16'h89fd;
17'h13799:	data_out=16'h9fa;
17'h1379a:	data_out=16'h9ab;
17'h1379b:	data_out=16'h8843;
17'h1379c:	data_out=16'h9cd;
17'h1379d:	data_out=16'ha00;
17'h1379e:	data_out=16'h8165;
17'h1379f:	data_out=16'h8891;
17'h137a0:	data_out=16'ha00;
17'h137a1:	data_out=16'h9f3;
17'h137a2:	data_out=16'h89fc;
17'h137a3:	data_out=16'h6bd;
17'h137a4:	data_out=16'h667;
17'h137a5:	data_out=16'h89fd;
17'h137a6:	data_out=16'h89e1;
17'h137a7:	data_out=16'h9fc;
17'h137a8:	data_out=16'h9f0;
17'h137a9:	data_out=16'h9ec;
17'h137aa:	data_out=16'h88c5;
17'h137ab:	data_out=16'h9f5;
17'h137ac:	data_out=16'h89a2;
17'h137ad:	data_out=16'h9fa;
17'h137ae:	data_out=16'h8067;
17'h137af:	data_out=16'h9f6;
17'h137b0:	data_out=16'h33a;
17'h137b1:	data_out=16'ha00;
17'h137b2:	data_out=16'h9e1;
17'h137b3:	data_out=16'he0;
17'h137b4:	data_out=16'ha00;
17'h137b5:	data_out=16'h3b4;
17'h137b6:	data_out=16'h883d;
17'h137b7:	data_out=16'h385;
17'h137b8:	data_out=16'ha00;
17'h137b9:	data_out=16'h19;
17'h137ba:	data_out=16'h89ff;
17'h137bb:	data_out=16'h86e9;
17'h137bc:	data_out=16'ha00;
17'h137bd:	data_out=16'h9c2;
17'h137be:	data_out=16'h9f0;
17'h137bf:	data_out=16'h894;
17'h137c0:	data_out=16'h83bf;
17'h137c1:	data_out=16'h89fe;
17'h137c2:	data_out=16'h8a00;
17'h137c3:	data_out=16'h1ff;
17'h137c4:	data_out=16'h920;
17'h137c5:	data_out=16'h81ea;
17'h137c6:	data_out=16'h9f8;
17'h137c7:	data_out=16'h89ff;
17'h137c8:	data_out=16'h8a00;
17'h137c9:	data_out=16'h89fc;
17'h137ca:	data_out=16'h8993;
17'h137cb:	data_out=16'h8a00;
17'h137cc:	data_out=16'h8a00;
17'h137cd:	data_out=16'h89f9;
17'h137ce:	data_out=16'h3c2;
17'h137cf:	data_out=16'h8a00;
17'h137d0:	data_out=16'h89e9;
17'h137d1:	data_out=16'h8a00;
17'h137d2:	data_out=16'h8a00;
17'h137d3:	data_out=16'ha00;
17'h137d4:	data_out=16'ha00;
17'h137d5:	data_out=16'h8a00;
17'h137d6:	data_out=16'h87f2;
17'h137d7:	data_out=16'h836b;
17'h137d8:	data_out=16'h8a00;
17'h137d9:	data_out=16'h24c;
17'h137da:	data_out=16'h400;
17'h137db:	data_out=16'ha00;
17'h137dc:	data_out=16'h9d3;
17'h137dd:	data_out=16'h972;
17'h137de:	data_out=16'ha00;
17'h137df:	data_out=16'h88e7;
17'h137e0:	data_out=16'h89e1;
17'h137e1:	data_out=16'h9f6;
17'h137e2:	data_out=16'h82cf;
17'h137e3:	data_out=16'h3ed;
17'h137e4:	data_out=16'ha00;
17'h137e5:	data_out=16'h9e4;
17'h137e6:	data_out=16'h89dc;
17'h137e7:	data_out=16'h8639;
17'h137e8:	data_out=16'h9f1;
17'h137e9:	data_out=16'h89f4;
17'h137ea:	data_out=16'h9f7;
17'h137eb:	data_out=16'h8b8;
17'h137ec:	data_out=16'h9fe;
17'h137ed:	data_out=16'h402;
17'h137ee:	data_out=16'h9f7;
17'h137ef:	data_out=16'h36f;
17'h137f0:	data_out=16'h9f6;
17'h137f1:	data_out=16'h89e8;
17'h137f2:	data_out=16'h9e8;
17'h137f3:	data_out=16'ha00;
17'h137f4:	data_out=16'h315;
17'h137f5:	data_out=16'h712;
17'h137f6:	data_out=16'h9f4;
17'h137f7:	data_out=16'h8a00;
17'h137f8:	data_out=16'h82cb;
17'h137f9:	data_out=16'h8a00;
17'h137fa:	data_out=16'h252;
17'h137fb:	data_out=16'h9f0;
17'h137fc:	data_out=16'h89f8;
17'h137fd:	data_out=16'h894f;
17'h137fe:	data_out=16'h9e8;
17'h137ff:	data_out=16'h89f6;
17'h13800:	data_out=16'h9ea;
17'h13801:	data_out=16'ha00;
17'h13802:	data_out=16'h89ee;
17'h13803:	data_out=16'h8906;
17'h13804:	data_out=16'h854a;
17'h13805:	data_out=16'h37b;
17'h13806:	data_out=16'h2b6;
17'h13807:	data_out=16'h8a00;
17'h13808:	data_out=16'h8934;
17'h13809:	data_out=16'h8a00;
17'h1380a:	data_out=16'ha00;
17'h1380b:	data_out=16'h8310;
17'h1380c:	data_out=16'h8a00;
17'h1380d:	data_out=16'h8a00;
17'h1380e:	data_out=16'h9fe;
17'h1380f:	data_out=16'h89fe;
17'h13810:	data_out=16'h89d2;
17'h13811:	data_out=16'ha00;
17'h13812:	data_out=16'h8a00;
17'h13813:	data_out=16'ha00;
17'h13814:	data_out=16'h88fd;
17'h13815:	data_out=16'h8387;
17'h13816:	data_out=16'h89d4;
17'h13817:	data_out=16'h8908;
17'h13818:	data_out=16'h8a00;
17'h13819:	data_out=16'h9f3;
17'h1381a:	data_out=16'h646;
17'h1381b:	data_out=16'h840e;
17'h1381c:	data_out=16'h92f;
17'h1381d:	data_out=16'ha00;
17'h1381e:	data_out=16'h88e4;
17'h1381f:	data_out=16'h898c;
17'h13820:	data_out=16'h9d8;
17'h13821:	data_out=16'h9fd;
17'h13822:	data_out=16'h8922;
17'h13823:	data_out=16'h9c6;
17'h13824:	data_out=16'h966;
17'h13825:	data_out=16'h89c7;
17'h13826:	data_out=16'h882d;
17'h13827:	data_out=16'h9f1;
17'h13828:	data_out=16'h9f9;
17'h13829:	data_out=16'h9ee;
17'h1382a:	data_out=16'h8831;
17'h1382b:	data_out=16'h9e0;
17'h1382c:	data_out=16'h89c9;
17'h1382d:	data_out=16'ha00;
17'h1382e:	data_out=16'h82bb;
17'h1382f:	data_out=16'h9e9;
17'h13830:	data_out=16'h1cb;
17'h13831:	data_out=16'ha00;
17'h13832:	data_out=16'h9e2;
17'h13833:	data_out=16'h89bb;
17'h13834:	data_out=16'ha00;
17'h13835:	data_out=16'h89ab;
17'h13836:	data_out=16'h871b;
17'h13837:	data_out=16'h897b;
17'h13838:	data_out=16'ha00;
17'h13839:	data_out=16'h89bc;
17'h1383a:	data_out=16'h89fa;
17'h1383b:	data_out=16'h89ee;
17'h1383c:	data_out=16'ha00;
17'h1383d:	data_out=16'h9a2;
17'h1383e:	data_out=16'h9f9;
17'h1383f:	data_out=16'h372;
17'h13840:	data_out=16'h99b;
17'h13841:	data_out=16'h89f3;
17'h13842:	data_out=16'h89d5;
17'h13843:	data_out=16'h7a8;
17'h13844:	data_out=16'h1c9;
17'h13845:	data_out=16'h83e7;
17'h13846:	data_out=16'h9fb;
17'h13847:	data_out=16'h89ff;
17'h13848:	data_out=16'h8a00;
17'h13849:	data_out=16'h8969;
17'h1384a:	data_out=16'h89c2;
17'h1384b:	data_out=16'h8a00;
17'h1384c:	data_out=16'h89f9;
17'h1384d:	data_out=16'h896b;
17'h1384e:	data_out=16'h30d;
17'h1384f:	data_out=16'h89fa;
17'h13850:	data_out=16'h89fb;
17'h13851:	data_out=16'h8a00;
17'h13852:	data_out=16'h8a00;
17'h13853:	data_out=16'h9f9;
17'h13854:	data_out=16'h9ea;
17'h13855:	data_out=16'h89d8;
17'h13856:	data_out=16'h557;
17'h13857:	data_out=16'h832c;
17'h13858:	data_out=16'h89f6;
17'h13859:	data_out=16'h567;
17'h1385a:	data_out=16'h80cd;
17'h1385b:	data_out=16'ha00;
17'h1385c:	data_out=16'h92e;
17'h1385d:	data_out=16'h9c2;
17'h1385e:	data_out=16'ha00;
17'h1385f:	data_out=16'h8978;
17'h13860:	data_out=16'h8762;
17'h13861:	data_out=16'h9e5;
17'h13862:	data_out=16'h8114;
17'h13863:	data_out=16'h89a4;
17'h13864:	data_out=16'ha00;
17'h13865:	data_out=16'h9e1;
17'h13866:	data_out=16'h899c;
17'h13867:	data_out=16'h89a4;
17'h13868:	data_out=16'h9fb;
17'h13869:	data_out=16'h89ce;
17'h1386a:	data_out=16'h9ff;
17'h1386b:	data_out=16'h30e;
17'h1386c:	data_out=16'h9c0;
17'h1386d:	data_out=16'h8997;
17'h1386e:	data_out=16'h9ff;
17'h1386f:	data_out=16'h19a;
17'h13870:	data_out=16'h9fe;
17'h13871:	data_out=16'h89fb;
17'h13872:	data_out=16'h9db;
17'h13873:	data_out=16'ha00;
17'h13874:	data_out=16'h1f6;
17'h13875:	data_out=16'h5e4;
17'h13876:	data_out=16'h47f;
17'h13877:	data_out=16'h8a00;
17'h13878:	data_out=16'h45c;
17'h13879:	data_out=16'h8a00;
17'h1387a:	data_out=16'h893e;
17'h1387b:	data_out=16'h9f9;
17'h1387c:	data_out=16'h89fe;
17'h1387d:	data_out=16'h89fc;
17'h1387e:	data_out=16'h9e4;
17'h1387f:	data_out=16'h89fa;
17'h13880:	data_out=16'h9f9;
17'h13881:	data_out=16'ha00;
17'h13882:	data_out=16'h899c;
17'h13883:	data_out=16'h89f8;
17'h13884:	data_out=16'h38c;
17'h13885:	data_out=16'h648;
17'h13886:	data_out=16'h89ff;
17'h13887:	data_out=16'h8a00;
17'h13888:	data_out=16'h879c;
17'h13889:	data_out=16'h89f6;
17'h1388a:	data_out=16'ha00;
17'h1388b:	data_out=16'h87e8;
17'h1388c:	data_out=16'h89fc;
17'h1388d:	data_out=16'h8a00;
17'h1388e:	data_out=16'h888;
17'h1388f:	data_out=16'h89e8;
17'h13890:	data_out=16'h89eb;
17'h13891:	data_out=16'ha00;
17'h13892:	data_out=16'h8a00;
17'h13893:	data_out=16'ha00;
17'h13894:	data_out=16'h89fa;
17'h13895:	data_out=16'h893e;
17'h13896:	data_out=16'h89f3;
17'h13897:	data_out=16'h89fe;
17'h13898:	data_out=16'h8a00;
17'h13899:	data_out=16'h9f1;
17'h1389a:	data_out=16'h97f;
17'h1389b:	data_out=16'h85aa;
17'h1389c:	data_out=16'h594;
17'h1389d:	data_out=16'ha00;
17'h1389e:	data_out=16'h89f0;
17'h1389f:	data_out=16'h89ef;
17'h138a0:	data_out=16'h9f7;
17'h138a1:	data_out=16'h663;
17'h138a2:	data_out=16'h88fc;
17'h138a3:	data_out=16'h9ff;
17'h138a4:	data_out=16'h9ff;
17'h138a5:	data_out=16'h893c;
17'h138a6:	data_out=16'h869f;
17'h138a7:	data_out=16'h9fb;
17'h138a8:	data_out=16'h4f6;
17'h138a9:	data_out=16'h9eb;
17'h138aa:	data_out=16'h8799;
17'h138ab:	data_out=16'h9dc;
17'h138ac:	data_out=16'h89f4;
17'h138ad:	data_out=16'h74c;
17'h138ae:	data_out=16'h8518;
17'h138af:	data_out=16'h9f6;
17'h138b0:	data_out=16'h29d;
17'h138b1:	data_out=16'ha00;
17'h138b2:	data_out=16'ha00;
17'h138b3:	data_out=16'h89ff;
17'h138b4:	data_out=16'ha00;
17'h138b5:	data_out=16'h818f;
17'h138b6:	data_out=16'h833e;
17'h138b7:	data_out=16'h87e6;
17'h138b8:	data_out=16'ha00;
17'h138b9:	data_out=16'h89ff;
17'h138ba:	data_out=16'h89f5;
17'h138bb:	data_out=16'h871e;
17'h138bc:	data_out=16'ha00;
17'h138bd:	data_out=16'h9fa;
17'h138be:	data_out=16'h4ff;
17'h138bf:	data_out=16'h640;
17'h138c0:	data_out=16'ha00;
17'h138c1:	data_out=16'h89c7;
17'h138c2:	data_out=16'h89a3;
17'h138c3:	data_out=16'h9ea;
17'h138c4:	data_out=16'h807;
17'h138c5:	data_out=16'h896c;
17'h138c6:	data_out=16'h9fc;
17'h138c7:	data_out=16'h8a00;
17'h138c8:	data_out=16'h89ff;
17'h138c9:	data_out=16'h87e9;
17'h138ca:	data_out=16'h86fe;
17'h138cb:	data_out=16'h8a00;
17'h138cc:	data_out=16'h89e0;
17'h138cd:	data_out=16'h894d;
17'h138ce:	data_out=16'h475;
17'h138cf:	data_out=16'h89e5;
17'h138d0:	data_out=16'h89f6;
17'h138d1:	data_out=16'h8a00;
17'h138d2:	data_out=16'h89ce;
17'h138d3:	data_out=16'h9f9;
17'h138d4:	data_out=16'h9f6;
17'h138d5:	data_out=16'h89e1;
17'h138d6:	data_out=16'h211;
17'h138d7:	data_out=16'h8530;
17'h138d8:	data_out=16'h89d4;
17'h138d9:	data_out=16'h9ff;
17'h138da:	data_out=16'h8a00;
17'h138db:	data_out=16'ha00;
17'h138dc:	data_out=16'h9e7;
17'h138dd:	data_out=16'h9fa;
17'h138de:	data_out=16'ha00;
17'h138df:	data_out=16'h89ab;
17'h138e0:	data_out=16'h87b5;
17'h138e1:	data_out=16'ha00;
17'h138e2:	data_out=16'h86de;
17'h138e3:	data_out=16'h8a00;
17'h138e4:	data_out=16'ha00;
17'h138e5:	data_out=16'ha00;
17'h138e6:	data_out=16'h89ad;
17'h138e7:	data_out=16'h89fd;
17'h138e8:	data_out=16'h560;
17'h138e9:	data_out=16'h898d;
17'h138ea:	data_out=16'h9bc;
17'h138eb:	data_out=16'h3ea;
17'h138ec:	data_out=16'h9ee;
17'h138ed:	data_out=16'h8a00;
17'h138ee:	data_out=16'h9b8;
17'h138ef:	data_out=16'h5fb;
17'h138f0:	data_out=16'h923;
17'h138f1:	data_out=16'h89fd;
17'h138f2:	data_out=16'ha00;
17'h138f3:	data_out=16'ha00;
17'h138f4:	data_out=16'h2d2;
17'h138f5:	data_out=16'h78d;
17'h138f6:	data_out=16'h862e;
17'h138f7:	data_out=16'h89fb;
17'h138f8:	data_out=16'h990;
17'h138f9:	data_out=16'h8a00;
17'h138fa:	data_out=16'h89fe;
17'h138fb:	data_out=16'h500;
17'h138fc:	data_out=16'h8a00;
17'h138fd:	data_out=16'h89f2;
17'h138fe:	data_out=16'h9eb;
17'h138ff:	data_out=16'h89fb;
17'h13900:	data_out=16'h9eb;
17'h13901:	data_out=16'ha00;
17'h13902:	data_out=16'h8883;
17'h13903:	data_out=16'h89cf;
17'h13904:	data_out=16'h854f;
17'h13905:	data_out=16'h9f7;
17'h13906:	data_out=16'h89fd;
17'h13907:	data_out=16'h8a00;
17'h13908:	data_out=16'h8631;
17'h13909:	data_out=16'h89f0;
17'h1390a:	data_out=16'ha00;
17'h1390b:	data_out=16'h87ce;
17'h1390c:	data_out=16'h8996;
17'h1390d:	data_out=16'h8a00;
17'h1390e:	data_out=16'h608;
17'h1390f:	data_out=16'h8978;
17'h13910:	data_out=16'h89a2;
17'h13911:	data_out=16'ha00;
17'h13912:	data_out=16'h8a00;
17'h13913:	data_out=16'h839a;
17'h13914:	data_out=16'h89c4;
17'h13915:	data_out=16'h89e2;
17'h13916:	data_out=16'h89d7;
17'h13917:	data_out=16'h89b3;
17'h13918:	data_out=16'h8a00;
17'h13919:	data_out=16'h85d2;
17'h1391a:	data_out=16'ha00;
17'h1391b:	data_out=16'h8909;
17'h1391c:	data_out=16'h850e;
17'h1391d:	data_out=16'ha00;
17'h1391e:	data_out=16'h89b7;
17'h1391f:	data_out=16'h89e4;
17'h13920:	data_out=16'h17;
17'h13921:	data_out=16'h42c;
17'h13922:	data_out=16'h8983;
17'h13923:	data_out=16'h3e3;
17'h13924:	data_out=16'h3bc;
17'h13925:	data_out=16'h88b1;
17'h13926:	data_out=16'h84d6;
17'h13927:	data_out=16'ha00;
17'h13928:	data_out=16'h341;
17'h13929:	data_out=16'h9ed;
17'h1392a:	data_out=16'h8575;
17'h1392b:	data_out=16'h82ec;
17'h1392c:	data_out=16'h89e9;
17'h1392d:	data_out=16'h8873;
17'h1392e:	data_out=16'h85cb;
17'h1392f:	data_out=16'h8540;
17'h13930:	data_out=16'h45d;
17'h13931:	data_out=16'ha00;
17'h13932:	data_out=16'ha00;
17'h13933:	data_out=16'h89f8;
17'h13934:	data_out=16'ha00;
17'h13935:	data_out=16'h846b;
17'h13936:	data_out=16'h82f6;
17'h13937:	data_out=16'h86fb;
17'h13938:	data_out=16'ha00;
17'h13939:	data_out=16'h89ff;
17'h1393a:	data_out=16'h89f1;
17'h1393b:	data_out=16'h8061;
17'h1393c:	data_out=16'ha00;
17'h1393d:	data_out=16'h86e9;
17'h1393e:	data_out=16'h350;
17'h1393f:	data_out=16'h9f7;
17'h13940:	data_out=16'ha00;
17'h13941:	data_out=16'h8976;
17'h13942:	data_out=16'h8894;
17'h13943:	data_out=16'ha00;
17'h13944:	data_out=16'ha00;
17'h13945:	data_out=16'h89e4;
17'h13946:	data_out=16'ha00;
17'h13947:	data_out=16'h8a00;
17'h13948:	data_out=16'h89fc;
17'h13949:	data_out=16'h8718;
17'h1394a:	data_out=16'h300;
17'h1394b:	data_out=16'h89df;
17'h1394c:	data_out=16'h89e0;
17'h1394d:	data_out=16'h89b8;
17'h1394e:	data_out=16'h271;
17'h1394f:	data_out=16'h89d2;
17'h13950:	data_out=16'h89f5;
17'h13951:	data_out=16'h8a00;
17'h13952:	data_out=16'h88d4;
17'h13953:	data_out=16'h9fe;
17'h13954:	data_out=16'h802b;
17'h13955:	data_out=16'h895d;
17'h13956:	data_out=16'h83fd;
17'h13957:	data_out=16'h88bd;
17'h13958:	data_out=16'h89a8;
17'h13959:	data_out=16'h7a1;
17'h1395a:	data_out=16'h89dc;
17'h1395b:	data_out=16'ha00;
17'h1395c:	data_out=16'h9ed;
17'h1395d:	data_out=16'ha00;
17'h1395e:	data_out=16'h8283;
17'h1395f:	data_out=16'h89ee;
17'h13960:	data_out=16'h767;
17'h13961:	data_out=16'ha00;
17'h13962:	data_out=16'h87f0;
17'h13963:	data_out=16'h89df;
17'h13964:	data_out=16'h9f9;
17'h13965:	data_out=16'ha00;
17'h13966:	data_out=16'h87fa;
17'h13967:	data_out=16'h89fb;
17'h13968:	data_out=16'h346;
17'h13969:	data_out=16'h8986;
17'h1396a:	data_out=16'h708;
17'h1396b:	data_out=16'h8686;
17'h1396c:	data_out=16'h9ee;
17'h1396d:	data_out=16'h89e5;
17'h1396e:	data_out=16'h708;
17'h1396f:	data_out=16'ha00;
17'h13970:	data_out=16'h694;
17'h13971:	data_out=16'h899b;
17'h13972:	data_out=16'ha00;
17'h13973:	data_out=16'ha00;
17'h13974:	data_out=16'h4a7;
17'h13975:	data_out=16'h3cf;
17'h13976:	data_out=16'h887a;
17'h13977:	data_out=16'h89b3;
17'h13978:	data_out=16'ha00;
17'h13979:	data_out=16'h89f4;
17'h1397a:	data_out=16'h89b9;
17'h1397b:	data_out=16'h355;
17'h1397c:	data_out=16'h8a00;
17'h1397d:	data_out=16'h89ec;
17'h1397e:	data_out=16'h80cf;
17'h1397f:	data_out=16'h89fe;
17'h13980:	data_out=16'h658;
17'h13981:	data_out=16'ha00;
17'h13982:	data_out=16'h880d;
17'h13983:	data_out=16'h89fe;
17'h13984:	data_out=16'h8265;
17'h13985:	data_out=16'h8253;
17'h13986:	data_out=16'h89ff;
17'h13987:	data_out=16'h886f;
17'h13988:	data_out=16'h8480;
17'h13989:	data_out=16'h89e2;
17'h1398a:	data_out=16'ha00;
17'h1398b:	data_out=16'h8955;
17'h1398c:	data_out=16'h84b2;
17'h1398d:	data_out=16'h8a00;
17'h1398e:	data_out=16'h9ff;
17'h1398f:	data_out=16'h88db;
17'h13990:	data_out=16'h8998;
17'h13991:	data_out=16'ha00;
17'h13992:	data_out=16'h8a00;
17'h13993:	data_out=16'h8953;
17'h13994:	data_out=16'h89e7;
17'h13995:	data_out=16'h89e0;
17'h13996:	data_out=16'h89e3;
17'h13997:	data_out=16'h89d9;
17'h13998:	data_out=16'h8a00;
17'h13999:	data_out=16'h9ee;
17'h1399a:	data_out=16'h6b4;
17'h1399b:	data_out=16'h8935;
17'h1399c:	data_out=16'h89f9;
17'h1399d:	data_out=16'ha00;
17'h1399e:	data_out=16'h89bf;
17'h1399f:	data_out=16'h89c1;
17'h139a0:	data_out=16'h8919;
17'h139a1:	data_out=16'h9ff;
17'h139a2:	data_out=16'h89ac;
17'h139a3:	data_out=16'h9ff;
17'h139a4:	data_out=16'h9ff;
17'h139a5:	data_out=16'h889d;
17'h139a6:	data_out=16'h55d;
17'h139a7:	data_out=16'ha00;
17'h139a8:	data_out=16'h9ff;
17'h139a9:	data_out=16'h9f0;
17'h139aa:	data_out=16'h8595;
17'h139ab:	data_out=16'h84b7;
17'h139ac:	data_out=16'h89eb;
17'h139ad:	data_out=16'h8859;
17'h139ae:	data_out=16'h87fc;
17'h139af:	data_out=16'h886c;
17'h139b0:	data_out=16'h625;
17'h139b1:	data_out=16'ha00;
17'h139b2:	data_out=16'h9ff;
17'h139b3:	data_out=16'h89fe;
17'h139b4:	data_out=16'ha00;
17'h139b5:	data_out=16'hb7;
17'h139b6:	data_out=16'h8360;
17'h139b7:	data_out=16'h8736;
17'h139b8:	data_out=16'h9fd;
17'h139b9:	data_out=16'h8a00;
17'h139ba:	data_out=16'h89da;
17'h139bb:	data_out=16'h9fa;
17'h139bc:	data_out=16'h8297;
17'h139bd:	data_out=16'h8917;
17'h139be:	data_out=16'h9ff;
17'h139bf:	data_out=16'h822a;
17'h139c0:	data_out=16'ha00;
17'h139c1:	data_out=16'h895f;
17'h139c2:	data_out=16'h877a;
17'h139c3:	data_out=16'h9fd;
17'h139c4:	data_out=16'h9ff;
17'h139c5:	data_out=16'h89e2;
17'h139c6:	data_out=16'h9ff;
17'h139c7:	data_out=16'h89ee;
17'h139c8:	data_out=16'h89eb;
17'h139c9:	data_out=16'h869e;
17'h139ca:	data_out=16'h9ff;
17'h139cb:	data_out=16'h89b9;
17'h139cc:	data_out=16'h89d1;
17'h139cd:	data_out=16'h89bd;
17'h139ce:	data_out=16'h88e2;
17'h139cf:	data_out=16'h8971;
17'h139d0:	data_out=16'h89fc;
17'h139d1:	data_out=16'h8a00;
17'h139d2:	data_out=16'h889;
17'h139d3:	data_out=16'h80f2;
17'h139d4:	data_out=16'h88c4;
17'h139d5:	data_out=16'h8980;
17'h139d6:	data_out=16'h8443;
17'h139d7:	data_out=16'h890a;
17'h139d8:	data_out=16'h89cb;
17'h139d9:	data_out=16'ha00;
17'h139da:	data_out=16'h89f3;
17'h139db:	data_out=16'ha00;
17'h139dc:	data_out=16'h1f5;
17'h139dd:	data_out=16'h853f;
17'h139de:	data_out=16'h853a;
17'h139df:	data_out=16'h89d9;
17'h139e0:	data_out=16'h9f6;
17'h139e1:	data_out=16'h9fe;
17'h139e2:	data_out=16'h894b;
17'h139e3:	data_out=16'h89e5;
17'h139e4:	data_out=16'h9fe;
17'h139e5:	data_out=16'ha00;
17'h139e6:	data_out=16'hba;
17'h139e7:	data_out=16'h89f7;
17'h139e8:	data_out=16'h9ff;
17'h139e9:	data_out=16'h8990;
17'h139ea:	data_out=16'ha00;
17'h139eb:	data_out=16'h878a;
17'h139ec:	data_out=16'h9f2;
17'h139ed:	data_out=16'h89e8;
17'h139ee:	data_out=16'ha00;
17'h139ef:	data_out=16'ha00;
17'h139f0:	data_out=16'ha00;
17'h139f1:	data_out=16'h892d;
17'h139f2:	data_out=16'ha00;
17'h139f3:	data_out=16'ha00;
17'h139f4:	data_out=16'h622;
17'h139f5:	data_out=16'he3;
17'h139f6:	data_out=16'h88a8;
17'h139f7:	data_out=16'h8995;
17'h139f8:	data_out=16'h9f5;
17'h139f9:	data_out=16'h89b0;
17'h139fa:	data_out=16'h89d2;
17'h139fb:	data_out=16'h9ff;
17'h139fc:	data_out=16'h89ff;
17'h139fd:	data_out=16'h89e1;
17'h139fe:	data_out=16'h898e;
17'h139ff:	data_out=16'h8a00;
17'h13a00:	data_out=16'h819f;
17'h13a01:	data_out=16'ha00;
17'h13a02:	data_out=16'h6e4;
17'h13a03:	data_out=16'h89ff;
17'h13a04:	data_out=16'h886;
17'h13a05:	data_out=16'h877d;
17'h13a06:	data_out=16'h89ff;
17'h13a07:	data_out=16'h9f4;
17'h13a08:	data_out=16'h664;
17'h13a09:	data_out=16'h89d5;
17'h13a0a:	data_out=16'ha00;
17'h13a0b:	data_out=16'h898c;
17'h13a0c:	data_out=16'ha00;
17'h13a0d:	data_out=16'h8a00;
17'h13a0e:	data_out=16'h9ff;
17'h13a0f:	data_out=16'h8732;
17'h13a10:	data_out=16'h898f;
17'h13a11:	data_out=16'ha00;
17'h13a12:	data_out=16'h89f9;
17'h13a13:	data_out=16'h89b9;
17'h13a14:	data_out=16'h89ee;
17'h13a15:	data_out=16'h89f7;
17'h13a16:	data_out=16'h89f4;
17'h13a17:	data_out=16'h89f9;
17'h13a18:	data_out=16'h89fd;
17'h13a19:	data_out=16'h9fb;
17'h13a1a:	data_out=16'h7a2;
17'h13a1b:	data_out=16'h895c;
17'h13a1c:	data_out=16'h8a00;
17'h13a1d:	data_out=16'ha00;
17'h13a1e:	data_out=16'h89d4;
17'h13a1f:	data_out=16'h89d3;
17'h13a20:	data_out=16'h89ae;
17'h13a21:	data_out=16'h9ff;
17'h13a22:	data_out=16'h8902;
17'h13a23:	data_out=16'h9ff;
17'h13a24:	data_out=16'h9ff;
17'h13a25:	data_out=16'h85f9;
17'h13a26:	data_out=16'h9fc;
17'h13a27:	data_out=16'h683;
17'h13a28:	data_out=16'h9ff;
17'h13a29:	data_out=16'ha00;
17'h13a2a:	data_out=16'h822f;
17'h13a2b:	data_out=16'h88b2;
17'h13a2c:	data_out=16'h89fd;
17'h13a2d:	data_out=16'h882d;
17'h13a2e:	data_out=16'h8861;
17'h13a2f:	data_out=16'h89ab;
17'h13a30:	data_out=16'h9e5;
17'h13a31:	data_out=16'ha00;
17'h13a32:	data_out=16'h9fb;
17'h13a33:	data_out=16'h89f7;
17'h13a34:	data_out=16'ha00;
17'h13a35:	data_out=16'h222;
17'h13a36:	data_out=16'h8103;
17'h13a37:	data_out=16'h8203;
17'h13a38:	data_out=16'h28;
17'h13a39:	data_out=16'h89fe;
17'h13a3a:	data_out=16'h89cf;
17'h13a3b:	data_out=16'h9f1;
17'h13a3c:	data_out=16'h8771;
17'h13a3d:	data_out=16'h895d;
17'h13a3e:	data_out=16'h9ff;
17'h13a3f:	data_out=16'h8782;
17'h13a40:	data_out=16'ha00;
17'h13a41:	data_out=16'h8825;
17'h13a42:	data_out=16'h9fb;
17'h13a43:	data_out=16'h9f7;
17'h13a44:	data_out=16'h8645;
17'h13a45:	data_out=16'h89f9;
17'h13a46:	data_out=16'h9ff;
17'h13a47:	data_out=16'h89d8;
17'h13a48:	data_out=16'h89f7;
17'h13a49:	data_out=16'h82de;
17'h13a4a:	data_out=16'h9fd;
17'h13a4b:	data_out=16'h8303;
17'h13a4c:	data_out=16'h87d7;
17'h13a4d:	data_out=16'h895f;
17'h13a4e:	data_out=16'h8991;
17'h13a4f:	data_out=16'h830d;
17'h13a50:	data_out=16'h8a00;
17'h13a51:	data_out=16'h8a00;
17'h13a52:	data_out=16'h9ff;
17'h13a53:	data_out=16'h84ec;
17'h13a54:	data_out=16'h8953;
17'h13a55:	data_out=16'h896a;
17'h13a56:	data_out=16'h9f5;
17'h13a57:	data_out=16'h8856;
17'h13a58:	data_out=16'h89d6;
17'h13a59:	data_out=16'ha00;
17'h13a5a:	data_out=16'h89f4;
17'h13a5b:	data_out=16'h9fc;
17'h13a5c:	data_out=16'h899e;
17'h13a5d:	data_out=16'h84cd;
17'h13a5e:	data_out=16'h8635;
17'h13a5f:	data_out=16'h89d2;
17'h13a60:	data_out=16'h9f9;
17'h13a61:	data_out=16'h9e1;
17'h13a62:	data_out=16'h8971;
17'h13a63:	data_out=16'h89e7;
17'h13a64:	data_out=16'h9f9;
17'h13a65:	data_out=16'ha00;
17'h13a66:	data_out=16'h9e3;
17'h13a67:	data_out=16'h89df;
17'h13a68:	data_out=16'h9ff;
17'h13a69:	data_out=16'h899b;
17'h13a6a:	data_out=16'h9ff;
17'h13a6b:	data_out=16'h8935;
17'h13a6c:	data_out=16'h9dd;
17'h13a6d:	data_out=16'h89e8;
17'h13a6e:	data_out=16'h9ff;
17'h13a6f:	data_out=16'h9ed;
17'h13a70:	data_out=16'h9ff;
17'h13a71:	data_out=16'h88c0;
17'h13a72:	data_out=16'h952;
17'h13a73:	data_out=16'h9e5;
17'h13a74:	data_out=16'h9da;
17'h13a75:	data_out=16'h320;
17'h13a76:	data_out=16'h883d;
17'h13a77:	data_out=16'h88d5;
17'h13a78:	data_out=16'h9d9;
17'h13a79:	data_out=16'h897e;
17'h13a7a:	data_out=16'h89e0;
17'h13a7b:	data_out=16'h9ff;
17'h13a7c:	data_out=16'h89fa;
17'h13a7d:	data_out=16'h89f3;
17'h13a7e:	data_out=16'h8970;
17'h13a7f:	data_out=16'h8a00;
17'h13a80:	data_out=16'h840e;
17'h13a81:	data_out=16'ha00;
17'h13a82:	data_out=16'h9f6;
17'h13a83:	data_out=16'h8a00;
17'h13a84:	data_out=16'h839;
17'h13a85:	data_out=16'h806c;
17'h13a86:	data_out=16'h89fe;
17'h13a87:	data_out=16'ha00;
17'h13a88:	data_out=16'h5ec;
17'h13a89:	data_out=16'h89c9;
17'h13a8a:	data_out=16'h9c7;
17'h13a8b:	data_out=16'h899c;
17'h13a8c:	data_out=16'ha00;
17'h13a8d:	data_out=16'h8a00;
17'h13a8e:	data_out=16'h9fe;
17'h13a8f:	data_out=16'h85fd;
17'h13a90:	data_out=16'h89e6;
17'h13a91:	data_out=16'ha00;
17'h13a92:	data_out=16'h89ea;
17'h13a93:	data_out=16'h89ed;
17'h13a94:	data_out=16'h89ed;
17'h13a95:	data_out=16'h8a00;
17'h13a96:	data_out=16'h89fe;
17'h13a97:	data_out=16'h89fa;
17'h13a98:	data_out=16'h89f6;
17'h13a99:	data_out=16'h9ef;
17'h13a9a:	data_out=16'h98c;
17'h13a9b:	data_out=16'h89a7;
17'h13a9c:	data_out=16'h8a00;
17'h13a9d:	data_out=16'ha00;
17'h13a9e:	data_out=16'h89e3;
17'h13a9f:	data_out=16'h8995;
17'h13aa0:	data_out=16'h89f2;
17'h13aa1:	data_out=16'h9fe;
17'h13aa2:	data_out=16'h89eb;
17'h13aa3:	data_out=16'h9f7;
17'h13aa4:	data_out=16'h9f7;
17'h13aa5:	data_out=16'h87b5;
17'h13aa6:	data_out=16'h9df;
17'h13aa7:	data_out=16'h89a0;
17'h13aa8:	data_out=16'h9ff;
17'h13aa9:	data_out=16'ha00;
17'h13aaa:	data_out=16'h81e0;
17'h13aab:	data_out=16'h89be;
17'h13aac:	data_out=16'h8a00;
17'h13aad:	data_out=16'h88e3;
17'h13aae:	data_out=16'h88e9;
17'h13aaf:	data_out=16'h89f1;
17'h13ab0:	data_out=16'ha00;
17'h13ab1:	data_out=16'h9d5;
17'h13ab2:	data_out=16'h9b7;
17'h13ab3:	data_out=16'h89f5;
17'h13ab4:	data_out=16'ha00;
17'h13ab5:	data_out=16'h9f5;
17'h13ab6:	data_out=16'h824a;
17'h13ab7:	data_out=16'h9fa;
17'h13ab8:	data_out=16'h89fc;
17'h13ab9:	data_out=16'h8a00;
17'h13aba:	data_out=16'h89d4;
17'h13abb:	data_out=16'h982;
17'h13abc:	data_out=16'h88b5;
17'h13abd:	data_out=16'h89f4;
17'h13abe:	data_out=16'h9ff;
17'h13abf:	data_out=16'h802f;
17'h13ac0:	data_out=16'h9c4;
17'h13ac1:	data_out=16'h84c1;
17'h13ac2:	data_out=16'h9c7;
17'h13ac3:	data_out=16'ha00;
17'h13ac4:	data_out=16'h8080;
17'h13ac5:	data_out=16'h8a00;
17'h13ac6:	data_out=16'h9ff;
17'h13ac7:	data_out=16'h89de;
17'h13ac8:	data_out=16'h89f6;
17'h13ac9:	data_out=16'h8586;
17'h13aca:	data_out=16'h9ec;
17'h13acb:	data_out=16'h8d4;
17'h13acc:	data_out=16'h8836;
17'h13acd:	data_out=16'h89ee;
17'h13ace:	data_out=16'h89a8;
17'h13acf:	data_out=16'h10a;
17'h13ad0:	data_out=16'h8a00;
17'h13ad1:	data_out=16'h89d5;
17'h13ad2:	data_out=16'h9eb;
17'h13ad3:	data_out=16'h882f;
17'h13ad4:	data_out=16'h89dc;
17'h13ad5:	data_out=16'h88ee;
17'h13ad6:	data_out=16'h9e3;
17'h13ad7:	data_out=16'h8912;
17'h13ad8:	data_out=16'h89d7;
17'h13ad9:	data_out=16'h988;
17'h13ada:	data_out=16'h89d6;
17'h13adb:	data_out=16'h98a;
17'h13adc:	data_out=16'h89c3;
17'h13add:	data_out=16'h8818;
17'h13ade:	data_out=16'h881a;
17'h13adf:	data_out=16'h89f5;
17'h13ae0:	data_out=16'h9d6;
17'h13ae1:	data_out=16'h9b3;
17'h13ae2:	data_out=16'h8955;
17'h13ae3:	data_out=16'h89e9;
17'h13ae4:	data_out=16'h820;
17'h13ae5:	data_out=16'h9df;
17'h13ae6:	data_out=16'h9f1;
17'h13ae7:	data_out=16'h8974;
17'h13ae8:	data_out=16'h9ff;
17'h13ae9:	data_out=16'h8998;
17'h13aea:	data_out=16'h9fe;
17'h13aeb:	data_out=16'h89d5;
17'h13aec:	data_out=16'h96f;
17'h13aed:	data_out=16'h89eb;
17'h13aee:	data_out=16'h9fe;
17'h13aef:	data_out=16'h9c1;
17'h13af0:	data_out=16'h9fe;
17'h13af1:	data_out=16'h8817;
17'h13af2:	data_out=16'h8083;
17'h13af3:	data_out=16'h9a9;
17'h13af4:	data_out=16'h9ee;
17'h13af5:	data_out=16'h999;
17'h13af6:	data_out=16'h88ba;
17'h13af7:	data_out=16'h8980;
17'h13af8:	data_out=16'h9d9;
17'h13af9:	data_out=16'h89ad;
17'h13afa:	data_out=16'h89e4;
17'h13afb:	data_out=16'h9ff;
17'h13afc:	data_out=16'h89f5;
17'h13afd:	data_out=16'h89e2;
17'h13afe:	data_out=16'h8987;
17'h13aff:	data_out=16'h8a00;
17'h13b00:	data_out=16'h2e;
17'h13b01:	data_out=16'h9db;
17'h13b02:	data_out=16'h56e;
17'h13b03:	data_out=16'h89bd;
17'h13b04:	data_out=16'h8a00;
17'h13b05:	data_out=16'h86fa;
17'h13b06:	data_out=16'h8a00;
17'h13b07:	data_out=16'h9fb;
17'h13b08:	data_out=16'h86ba;
17'h13b09:	data_out=16'h8999;
17'h13b0a:	data_out=16'h96c;
17'h13b0b:	data_out=16'h89a8;
17'h13b0c:	data_out=16'ha00;
17'h13b0d:	data_out=16'h89d1;
17'h13b0e:	data_out=16'h9fc;
17'h13b0f:	data_out=16'h8442;
17'h13b10:	data_out=16'h89f3;
17'h13b11:	data_out=16'h8a00;
17'h13b12:	data_out=16'h89a9;
17'h13b13:	data_out=16'h89fb;
17'h13b14:	data_out=16'h896c;
17'h13b15:	data_out=16'h89ed;
17'h13b16:	data_out=16'h88ff;
17'h13b17:	data_out=16'h8945;
17'h13b18:	data_out=16'h89e6;
17'h13b19:	data_out=16'h9a8;
17'h13b1a:	data_out=16'h46a;
17'h13b1b:	data_out=16'h8919;
17'h13b1c:	data_out=16'h8a00;
17'h13b1d:	data_out=16'h989;
17'h13b1e:	data_out=16'h899d;
17'h13b1f:	data_out=16'h892b;
17'h13b20:	data_out=16'h89f4;
17'h13b21:	data_out=16'h9fc;
17'h13b22:	data_out=16'h89f9;
17'h13b23:	data_out=16'h742;
17'h13b24:	data_out=16'h72e;
17'h13b25:	data_out=16'h89b1;
17'h13b26:	data_out=16'h3d4;
17'h13b27:	data_out=16'h89f8;
17'h13b28:	data_out=16'h9fd;
17'h13b29:	data_out=16'ha00;
17'h13b2a:	data_out=16'h80ec;
17'h13b2b:	data_out=16'h89ef;
17'h13b2c:	data_out=16'h89bc;
17'h13b2d:	data_out=16'h88de;
17'h13b2e:	data_out=16'h882d;
17'h13b2f:	data_out=16'h89fa;
17'h13b30:	data_out=16'ha00;
17'h13b31:	data_out=16'h990;
17'h13b32:	data_out=16'h572;
17'h13b33:	data_out=16'h89d5;
17'h13b34:	data_out=16'h9ed;
17'h13b35:	data_out=16'h89fb;
17'h13b36:	data_out=16'h85a6;
17'h13b37:	data_out=16'h3e;
17'h13b38:	data_out=16'h8a00;
17'h13b39:	data_out=16'h89f0;
17'h13b3a:	data_out=16'h89cb;
17'h13b3b:	data_out=16'h81ca;
17'h13b3c:	data_out=16'h897a;
17'h13b3d:	data_out=16'h89fb;
17'h13b3e:	data_out=16'h9fd;
17'h13b3f:	data_out=16'h86e0;
17'h13b40:	data_out=16'h816;
17'h13b41:	data_out=16'h820b;
17'h13b42:	data_out=16'h9a7;
17'h13b43:	data_out=16'ha00;
17'h13b44:	data_out=16'h877b;
17'h13b45:	data_out=16'h89ea;
17'h13b46:	data_out=16'h9bc;
17'h13b47:	data_out=16'h89bc;
17'h13b48:	data_out=16'h89de;
17'h13b49:	data_out=16'h89a3;
17'h13b4a:	data_out=16'h99e;
17'h13b4b:	data_out=16'h9bb;
17'h13b4c:	data_out=16'h89d3;
17'h13b4d:	data_out=16'h89fb;
17'h13b4e:	data_out=16'h89c0;
17'h13b4f:	data_out=16'h888c;
17'h13b50:	data_out=16'h8a00;
17'h13b51:	data_out=16'h88ba;
17'h13b52:	data_out=16'h8cc;
17'h13b53:	data_out=16'h89be;
17'h13b54:	data_out=16'h89e4;
17'h13b55:	data_out=16'h83e1;
17'h13b56:	data_out=16'h883a;
17'h13b57:	data_out=16'h89b6;
17'h13b58:	data_out=16'h89a5;
17'h13b59:	data_out=16'h8a00;
17'h13b5a:	data_out=16'h8834;
17'h13b5b:	data_out=16'h8a00;
17'h13b5c:	data_out=16'h8907;
17'h13b5d:	data_out=16'h89a6;
17'h13b5e:	data_out=16'h88a8;
17'h13b5f:	data_out=16'h89f4;
17'h13b60:	data_out=16'h98d;
17'h13b61:	data_out=16'h5e3;
17'h13b62:	data_out=16'h8697;
17'h13b63:	data_out=16'h89c0;
17'h13b64:	data_out=16'h89fc;
17'h13b65:	data_out=16'h89d7;
17'h13b66:	data_out=16'h9fe;
17'h13b67:	data_out=16'h9fa;
17'h13b68:	data_out=16'h9fc;
17'h13b69:	data_out=16'h89d3;
17'h13b6a:	data_out=16'h9fb;
17'h13b6b:	data_out=16'h89c6;
17'h13b6c:	data_out=16'h980;
17'h13b6d:	data_out=16'h89c9;
17'h13b6e:	data_out=16'h9fb;
17'h13b6f:	data_out=16'h9ec;
17'h13b70:	data_out=16'h9fc;
17'h13b71:	data_out=16'h855d;
17'h13b72:	data_out=16'h8a00;
17'h13b73:	data_out=16'h83d6;
17'h13b74:	data_out=16'h9f7;
17'h13b75:	data_out=16'h7b4;
17'h13b76:	data_out=16'h89e5;
17'h13b77:	data_out=16'h89ac;
17'h13b78:	data_out=16'h9a2;
17'h13b79:	data_out=16'h89b1;
17'h13b7a:	data_out=16'h8993;
17'h13b7b:	data_out=16'h9fd;
17'h13b7c:	data_out=16'h89eb;
17'h13b7d:	data_out=16'h89b4;
17'h13b7e:	data_out=16'h898d;
17'h13b7f:	data_out=16'h8a00;
17'h13b80:	data_out=16'h9c9;
17'h13b81:	data_out=16'h9e8;
17'h13b82:	data_out=16'h85a6;
17'h13b83:	data_out=16'h89ae;
17'h13b84:	data_out=16'h861f;
17'h13b85:	data_out=16'h776;
17'h13b86:	data_out=16'h8a00;
17'h13b87:	data_out=16'ha00;
17'h13b88:	data_out=16'h8779;
17'h13b89:	data_out=16'h899c;
17'h13b8a:	data_out=16'h967;
17'h13b8b:	data_out=16'h89d7;
17'h13b8c:	data_out=16'ha00;
17'h13b8d:	data_out=16'h898c;
17'h13b8e:	data_out=16'h9eb;
17'h13b8f:	data_out=16'h8513;
17'h13b90:	data_out=16'h89ff;
17'h13b91:	data_out=16'h8a00;
17'h13b92:	data_out=16'h897b;
17'h13b93:	data_out=16'h8a00;
17'h13b94:	data_out=16'h899e;
17'h13b95:	data_out=16'h863c;
17'h13b96:	data_out=16'h830e;
17'h13b97:	data_out=16'h8951;
17'h13b98:	data_out=16'h89d9;
17'h13b99:	data_out=16'h923;
17'h13b9a:	data_out=16'h946;
17'h13b9b:	data_out=16'h8973;
17'h13b9c:	data_out=16'h89e9;
17'h13b9d:	data_out=16'h221;
17'h13b9e:	data_out=16'h8991;
17'h13b9f:	data_out=16'h8943;
17'h13ba0:	data_out=16'h899a;
17'h13ba1:	data_out=16'h9ce;
17'h13ba2:	data_out=16'h8a00;
17'h13ba3:	data_out=16'h8a00;
17'h13ba4:	data_out=16'h8a00;
17'h13ba5:	data_out=16'h89ff;
17'h13ba6:	data_out=16'h89d6;
17'h13ba7:	data_out=16'h89c9;
17'h13ba8:	data_out=16'h9cf;
17'h13ba9:	data_out=16'ha00;
17'h13baa:	data_out=16'h1de;
17'h13bab:	data_out=16'h89e1;
17'h13bac:	data_out=16'h849a;
17'h13bad:	data_out=16'h89f8;
17'h13bae:	data_out=16'h890f;
17'h13baf:	data_out=16'h899b;
17'h13bb0:	data_out=16'h9fc;
17'h13bb1:	data_out=16'h9e0;
17'h13bb2:	data_out=16'h320;
17'h13bb3:	data_out=16'h89ad;
17'h13bb4:	data_out=16'h9f5;
17'h13bb5:	data_out=16'h89c8;
17'h13bb6:	data_out=16'h8598;
17'h13bb7:	data_out=16'h8651;
17'h13bb8:	data_out=16'h8a00;
17'h13bb9:	data_out=16'h89ca;
17'h13bba:	data_out=16'h89d2;
17'h13bbb:	data_out=16'h249;
17'h13bbc:	data_out=16'h89f9;
17'h13bbd:	data_out=16'h89b6;
17'h13bbe:	data_out=16'h9d3;
17'h13bbf:	data_out=16'h7a7;
17'h13bc0:	data_out=16'h6c5;
17'h13bc1:	data_out=16'h37e;
17'h13bc2:	data_out=16'h657;
17'h13bc3:	data_out=16'h9f3;
17'h13bc4:	data_out=16'h8b6;
17'h13bc5:	data_out=16'h85bb;
17'h13bc6:	data_out=16'h800;
17'h13bc7:	data_out=16'h89c7;
17'h13bc8:	data_out=16'h8999;
17'h13bc9:	data_out=16'h8a00;
17'h13bca:	data_out=16'h9ff;
17'h13bcb:	data_out=16'h9d7;
17'h13bcc:	data_out=16'h89ff;
17'h13bcd:	data_out=16'h8a00;
17'h13bce:	data_out=16'h8770;
17'h13bcf:	data_out=16'h89f9;
17'h13bd0:	data_out=16'h8992;
17'h13bd1:	data_out=16'h883f;
17'h13bd2:	data_out=16'h8937;
17'h13bd3:	data_out=16'h896a;
17'h13bd4:	data_out=16'h8986;
17'h13bd5:	data_out=16'h8674;
17'h13bd6:	data_out=16'h8a00;
17'h13bd7:	data_out=16'h8a00;
17'h13bd8:	data_out=16'h89dd;
17'h13bd9:	data_out=16'h8a00;
17'h13bda:	data_out=16'h8736;
17'h13bdb:	data_out=16'h89f1;
17'h13bdc:	data_out=16'h88eb;
17'h13bdd:	data_out=16'h8748;
17'h13bde:	data_out=16'h886f;
17'h13bdf:	data_out=16'h89dd;
17'h13be0:	data_out=16'h1;
17'h13be1:	data_out=16'h59d;
17'h13be2:	data_out=16'h887d;
17'h13be3:	data_out=16'h8990;
17'h13be4:	data_out=16'h89fc;
17'h13be5:	data_out=16'h8743;
17'h13be6:	data_out=16'ha00;
17'h13be7:	data_out=16'ha00;
17'h13be8:	data_out=16'h9ba;
17'h13be9:	data_out=16'h89e3;
17'h13bea:	data_out=16'h9eb;
17'h13beb:	data_out=16'h88db;
17'h13bec:	data_out=16'h9dd;
17'h13bed:	data_out=16'h8998;
17'h13bee:	data_out=16'h9eb;
17'h13bef:	data_out=16'ha00;
17'h13bf0:	data_out=16'h9eb;
17'h13bf1:	data_out=16'hc8;
17'h13bf2:	data_out=16'h89d3;
17'h13bf3:	data_out=16'h84b6;
17'h13bf4:	data_out=16'h9ef;
17'h13bf5:	data_out=16'h59c;
17'h13bf6:	data_out=16'h8825;
17'h13bf7:	data_out=16'h89b3;
17'h13bf8:	data_out=16'h4b3;
17'h13bf9:	data_out=16'h8932;
17'h13bfa:	data_out=16'h8986;
17'h13bfb:	data_out=16'h9d6;
17'h13bfc:	data_out=16'h89da;
17'h13bfd:	data_out=16'h8967;
17'h13bfe:	data_out=16'h89c8;
17'h13bff:	data_out=16'h89fc;
17'h13c00:	data_out=16'h9bb;
17'h13c01:	data_out=16'h9e5;
17'h13c02:	data_out=16'h89c8;
17'h13c03:	data_out=16'h89ad;
17'h13c04:	data_out=16'h919;
17'h13c05:	data_out=16'h9ef;
17'h13c06:	data_out=16'h89f6;
17'h13c07:	data_out=16'h9f4;
17'h13c08:	data_out=16'h89bd;
17'h13c09:	data_out=16'h89dc;
17'h13c0a:	data_out=16'h9a4;
17'h13c0b:	data_out=16'h89e7;
17'h13c0c:	data_out=16'h9e2;
17'h13c0d:	data_out=16'h895d;
17'h13c0e:	data_out=16'h5c3;
17'h13c0f:	data_out=16'h8976;
17'h13c10:	data_out=16'h89f6;
17'h13c11:	data_out=16'h8a00;
17'h13c12:	data_out=16'h89c6;
17'h13c13:	data_out=16'h8a00;
17'h13c14:	data_out=16'h89b9;
17'h13c15:	data_out=16'h805e;
17'h13c16:	data_out=16'h9ea;
17'h13c17:	data_out=16'h898c;
17'h13c18:	data_out=16'h8988;
17'h13c19:	data_out=16'h9b8;
17'h13c1a:	data_out=16'h9f1;
17'h13c1b:	data_out=16'h89c4;
17'h13c1c:	data_out=16'h89d5;
17'h13c1d:	data_out=16'h88e3;
17'h13c1e:	data_out=16'h89ad;
17'h13c1f:	data_out=16'h89a6;
17'h13c20:	data_out=16'h896d;
17'h13c21:	data_out=16'h490;
17'h13c22:	data_out=16'h8a00;
17'h13c23:	data_out=16'h8a00;
17'h13c24:	data_out=16'h8a00;
17'h13c25:	data_out=16'h8a00;
17'h13c26:	data_out=16'h8a00;
17'h13c27:	data_out=16'h89cd;
17'h13c28:	data_out=16'h2ac;
17'h13c29:	data_out=16'h9fd;
17'h13c2a:	data_out=16'h8779;
17'h13c2b:	data_out=16'h89f0;
17'h13c2c:	data_out=16'h9ed;
17'h13c2d:	data_out=16'h89ff;
17'h13c2e:	data_out=16'h89bb;
17'h13c2f:	data_out=16'h894a;
17'h13c30:	data_out=16'h9f5;
17'h13c31:	data_out=16'h9e3;
17'h13c32:	data_out=16'h458;
17'h13c33:	data_out=16'h89c6;
17'h13c34:	data_out=16'h9e4;
17'h13c35:	data_out=16'h8142;
17'h13c36:	data_out=16'h88e4;
17'h13c37:	data_out=16'h89d1;
17'h13c38:	data_out=16'h8a00;
17'h13c39:	data_out=16'h89d3;
17'h13c3a:	data_out=16'h89ee;
17'h13c3b:	data_out=16'h582;
17'h13c3c:	data_out=16'h89d7;
17'h13c3d:	data_out=16'h897b;
17'h13c3e:	data_out=16'h2aa;
17'h13c3f:	data_out=16'h9ee;
17'h13c40:	data_out=16'h3ac;
17'h13c41:	data_out=16'h41;
17'h13c42:	data_out=16'h89fe;
17'h13c43:	data_out=16'h819d;
17'h13c44:	data_out=16'h9de;
17'h13c45:	data_out=16'h41;
17'h13c46:	data_out=16'h612;
17'h13c47:	data_out=16'h89ff;
17'h13c48:	data_out=16'h89c8;
17'h13c49:	data_out=16'h8a00;
17'h13c4a:	data_out=16'ha00;
17'h13c4b:	data_out=16'h89be;
17'h13c4c:	data_out=16'h8a00;
17'h13c4d:	data_out=16'h89fe;
17'h13c4e:	data_out=16'h89fe;
17'h13c4f:	data_out=16'h8a00;
17'h13c50:	data_out=16'h895d;
17'h13c51:	data_out=16'h8912;
17'h13c52:	data_out=16'h8a00;
17'h13c53:	data_out=16'h89a6;
17'h13c54:	data_out=16'h898b;
17'h13c55:	data_out=16'h8994;
17'h13c56:	data_out=16'h8a00;
17'h13c57:	data_out=16'h8a00;
17'h13c58:	data_out=16'h89e0;
17'h13c59:	data_out=16'h89f1;
17'h13c5a:	data_out=16'h89b2;
17'h13c5b:	data_out=16'h809f;
17'h13c5c:	data_out=16'h8930;
17'h13c5d:	data_out=16'h8533;
17'h13c5e:	data_out=16'h8852;
17'h13c5f:	data_out=16'h89e7;
17'h13c60:	data_out=16'h8a00;
17'h13c61:	data_out=16'h97c;
17'h13c62:	data_out=16'h89b7;
17'h13c63:	data_out=16'h89b0;
17'h13c64:	data_out=16'h8a00;
17'h13c65:	data_out=16'h86a0;
17'h13c66:	data_out=16'ha00;
17'h13c67:	data_out=16'ha00;
17'h13c68:	data_out=16'h39d;
17'h13c69:	data_out=16'h89f8;
17'h13c6a:	data_out=16'h672;
17'h13c6b:	data_out=16'h8163;
17'h13c6c:	data_out=16'h9e0;
17'h13c6d:	data_out=16'h89b6;
17'h13c6e:	data_out=16'h674;
17'h13c6f:	data_out=16'ha00;
17'h13c70:	data_out=16'h627;
17'h13c71:	data_out=16'h859a;
17'h13c72:	data_out=16'h8955;
17'h13c73:	data_out=16'h343;
17'h13c74:	data_out=16'h9e7;
17'h13c75:	data_out=16'h9da;
17'h13c76:	data_out=16'h1df;
17'h13c77:	data_out=16'h89d5;
17'h13c78:	data_out=16'h8100;
17'h13c79:	data_out=16'h89da;
17'h13c7a:	data_out=16'h89a7;
17'h13c7b:	data_out=16'h2af;
17'h13c7c:	data_out=16'h890c;
17'h13c7d:	data_out=16'h88c7;
17'h13c7e:	data_out=16'h89d7;
17'h13c7f:	data_out=16'h8735;
17'h13c80:	data_out=16'h801b;
17'h13c81:	data_out=16'h9ff;
17'h13c82:	data_out=16'h89d4;
17'h13c83:	data_out=16'h899e;
17'h13c84:	data_out=16'h9f2;
17'h13c85:	data_out=16'ha00;
17'h13c86:	data_out=16'h89eb;
17'h13c87:	data_out=16'h800e;
17'h13c88:	data_out=16'h89bc;
17'h13c89:	data_out=16'h89fe;
17'h13c8a:	data_out=16'h9e9;
17'h13c8b:	data_out=16'h89ec;
17'h13c8c:	data_out=16'h89c6;
17'h13c8d:	data_out=16'h8948;
17'h13c8e:	data_out=16'h478;
17'h13c8f:	data_out=16'h89d0;
17'h13c90:	data_out=16'h89ee;
17'h13c91:	data_out=16'h8a00;
17'h13c92:	data_out=16'h89ec;
17'h13c93:	data_out=16'h89ee;
17'h13c94:	data_out=16'h89c2;
17'h13c95:	data_out=16'h9f7;
17'h13c96:	data_out=16'h9f3;
17'h13c97:	data_out=16'h8990;
17'h13c98:	data_out=16'h895f;
17'h13c99:	data_out=16'h9fc;
17'h13c9a:	data_out=16'ha00;
17'h13c9b:	data_out=16'h89ce;
17'h13c9c:	data_out=16'h897a;
17'h13c9d:	data_out=16'h89cc;
17'h13c9e:	data_out=16'h89b3;
17'h13c9f:	data_out=16'h89c0;
17'h13ca0:	data_out=16'h8857;
17'h13ca1:	data_out=16'h381;
17'h13ca2:	data_out=16'h89ef;
17'h13ca3:	data_out=16'h89f8;
17'h13ca4:	data_out=16'h89f8;
17'h13ca5:	data_out=16'h8a00;
17'h13ca6:	data_out=16'h8a00;
17'h13ca7:	data_out=16'h89e6;
17'h13ca8:	data_out=16'h1bd;
17'h13ca9:	data_out=16'h43a;
17'h13caa:	data_out=16'h8979;
17'h13cab:	data_out=16'h89ef;
17'h13cac:	data_out=16'h9f6;
17'h13cad:	data_out=16'h8a00;
17'h13cae:	data_out=16'h89f2;
17'h13caf:	data_out=16'h883e;
17'h13cb0:	data_out=16'ha00;
17'h13cb1:	data_out=16'h9f8;
17'h13cb2:	data_out=16'h833;
17'h13cb3:	data_out=16'h89c7;
17'h13cb4:	data_out=16'h3e1;
17'h13cb5:	data_out=16'h50;
17'h13cb6:	data_out=16'h899d;
17'h13cb7:	data_out=16'h89e8;
17'h13cb8:	data_out=16'h89f1;
17'h13cb9:	data_out=16'h89d3;
17'h13cba:	data_out=16'h89fa;
17'h13cbb:	data_out=16'h804;
17'h13cbc:	data_out=16'h892a;
17'h13cbd:	data_out=16'h8959;
17'h13cbe:	data_out=16'h1b5;
17'h13cbf:	data_out=16'ha00;
17'h13cc0:	data_out=16'h3b4;
17'h13cc1:	data_out=16'h8729;
17'h13cc2:	data_out=16'h89ff;
17'h13cc3:	data_out=16'h882c;
17'h13cc4:	data_out=16'h9f3;
17'h13cc5:	data_out=16'h9f7;
17'h13cc6:	data_out=16'h89d2;
17'h13cc7:	data_out=16'h8a00;
17'h13cc8:	data_out=16'h89f3;
17'h13cc9:	data_out=16'h89ff;
17'h13cca:	data_out=16'h849c;
17'h13ccb:	data_out=16'h89e2;
17'h13ccc:	data_out=16'h8a00;
17'h13ccd:	data_out=16'h89e1;
17'h13cce:	data_out=16'h89fc;
17'h13ccf:	data_out=16'h8a00;
17'h13cd0:	data_out=16'h8673;
17'h13cd1:	data_out=16'h2f5;
17'h13cd2:	data_out=16'h8a00;
17'h13cd3:	data_out=16'h89ac;
17'h13cd4:	data_out=16'h8987;
17'h13cd5:	data_out=16'h89a9;
17'h13cd6:	data_out=16'h89fb;
17'h13cd7:	data_out=16'h89fc;
17'h13cd8:	data_out=16'h8290;
17'h13cd9:	data_out=16'h89c1;
17'h13cda:	data_out=16'h89bc;
17'h13cdb:	data_out=16'h6fc;
17'h13cdc:	data_out=16'h8170;
17'h13cdd:	data_out=16'h85cc;
17'h13cde:	data_out=16'h883c;
17'h13cdf:	data_out=16'h89eb;
17'h13ce0:	data_out=16'h8a00;
17'h13ce1:	data_out=16'h9f8;
17'h13ce2:	data_out=16'h89cd;
17'h13ce3:	data_out=16'h89c0;
17'h13ce4:	data_out=16'h8a00;
17'h13ce5:	data_out=16'h8938;
17'h13ce6:	data_out=16'ha00;
17'h13ce7:	data_out=16'ha00;
17'h13ce8:	data_out=16'h2c1;
17'h13ce9:	data_out=16'h89fd;
17'h13cea:	data_out=16'h51f;
17'h13ceb:	data_out=16'h9ff;
17'h13cec:	data_out=16'h9fc;
17'h13ced:	data_out=16'h89c2;
17'h13cee:	data_out=16'h51f;
17'h13cef:	data_out=16'ha00;
17'h13cf0:	data_out=16'h4cd;
17'h13cf1:	data_out=16'h8763;
17'h13cf2:	data_out=16'h28f;
17'h13cf3:	data_out=16'h9ff;
17'h13cf4:	data_out=16'h9fb;
17'h13cf5:	data_out=16'h9f9;
17'h13cf6:	data_out=16'h7fb;
17'h13cf7:	data_out=16'h89f1;
17'h13cf8:	data_out=16'h89f3;
17'h13cf9:	data_out=16'h89cf;
17'h13cfa:	data_out=16'h89c0;
17'h13cfb:	data_out=16'h1b6;
17'h13cfc:	data_out=16'h88f6;
17'h13cfd:	data_out=16'h8295;
17'h13cfe:	data_out=16'h89e9;
17'h13cff:	data_out=16'h4d0;
17'h13d00:	data_out=16'h8796;
17'h13d01:	data_out=16'h8606;
17'h13d02:	data_out=16'h89b1;
17'h13d03:	data_out=16'h8987;
17'h13d04:	data_out=16'ha00;
17'h13d05:	data_out=16'ha00;
17'h13d06:	data_out=16'h89dc;
17'h13d07:	data_out=16'h89e1;
17'h13d08:	data_out=16'h89d9;
17'h13d09:	data_out=16'h89df;
17'h13d0a:	data_out=16'h9dc;
17'h13d0b:	data_out=16'h89eb;
17'h13d0c:	data_out=16'h89ff;
17'h13d0d:	data_out=16'h897d;
17'h13d0e:	data_out=16'h7b8;
17'h13d0f:	data_out=16'h89a1;
17'h13d10:	data_out=16'h89e1;
17'h13d11:	data_out=16'h8a00;
17'h13d12:	data_out=16'h89ac;
17'h13d13:	data_out=16'h89a0;
17'h13d14:	data_out=16'h89a5;
17'h13d15:	data_out=16'ha00;
17'h13d16:	data_out=16'h6d3;
17'h13d17:	data_out=16'h8987;
17'h13d18:	data_out=16'h890b;
17'h13d19:	data_out=16'h9e5;
17'h13d1a:	data_out=16'ha00;
17'h13d1b:	data_out=16'h89c2;
17'h13d1c:	data_out=16'h8980;
17'h13d1d:	data_out=16'h8a00;
17'h13d1e:	data_out=16'h8988;
17'h13d1f:	data_out=16'h8924;
17'h13d20:	data_out=16'h87e9;
17'h13d21:	data_out=16'h6ac;
17'h13d22:	data_out=16'h89de;
17'h13d23:	data_out=16'h8a00;
17'h13d24:	data_out=16'h8a00;
17'h13d25:	data_out=16'h89e0;
17'h13d26:	data_out=16'h89f9;
17'h13d27:	data_out=16'h89eb;
17'h13d28:	data_out=16'h4a7;
17'h13d29:	data_out=16'h9a;
17'h13d2a:	data_out=16'h89a0;
17'h13d2b:	data_out=16'h88b8;
17'h13d2c:	data_out=16'ha00;
17'h13d2d:	data_out=16'h8a00;
17'h13d2e:	data_out=16'h89e4;
17'h13d2f:	data_out=16'h8984;
17'h13d30:	data_out=16'h9ff;
17'h13d31:	data_out=16'h9f8;
17'h13d32:	data_out=16'h48c;
17'h13d33:	data_out=16'h899f;
17'h13d34:	data_out=16'h88d9;
17'h13d35:	data_out=16'h83c8;
17'h13d36:	data_out=16'h89b2;
17'h13d37:	data_out=16'h89c9;
17'h13d38:	data_out=16'h89f7;
17'h13d39:	data_out=16'h89a1;
17'h13d3a:	data_out=16'h89e3;
17'h13d3b:	data_out=16'h44e;
17'h13d3c:	data_out=16'h8827;
17'h13d3d:	data_out=16'h87ee;
17'h13d3e:	data_out=16'h496;
17'h13d3f:	data_out=16'ha00;
17'h13d40:	data_out=16'h8508;
17'h13d41:	data_out=16'h898a;
17'h13d42:	data_out=16'h8a00;
17'h13d43:	data_out=16'h89cd;
17'h13d44:	data_out=16'h9fd;
17'h13d45:	data_out=16'ha00;
17'h13d46:	data_out=16'h89e2;
17'h13d47:	data_out=16'h89fa;
17'h13d48:	data_out=16'h89e4;
17'h13d49:	data_out=16'h89e1;
17'h13d4a:	data_out=16'h8983;
17'h13d4b:	data_out=16'h8a00;
17'h13d4c:	data_out=16'h89f9;
17'h13d4d:	data_out=16'h89ad;
17'h13d4e:	data_out=16'h89f1;
17'h13d4f:	data_out=16'h8a00;
17'h13d50:	data_out=16'h805c;
17'h13d51:	data_out=16'h9eb;
17'h13d52:	data_out=16'h87bf;
17'h13d53:	data_out=16'h89d9;
17'h13d54:	data_out=16'h896b;
17'h13d55:	data_out=16'h8992;
17'h13d56:	data_out=16'hf;
17'h13d57:	data_out=16'h8986;
17'h13d58:	data_out=16'h16;
17'h13d59:	data_out=16'h89d7;
17'h13d5a:	data_out=16'h89c6;
17'h13d5b:	data_out=16'h978;
17'h13d5c:	data_out=16'h8784;
17'h13d5d:	data_out=16'h87e5;
17'h13d5e:	data_out=16'h899f;
17'h13d5f:	data_out=16'h89d5;
17'h13d60:	data_out=16'h8a00;
17'h13d61:	data_out=16'h9fa;
17'h13d62:	data_out=16'h89c8;
17'h13d63:	data_out=16'h89a0;
17'h13d64:	data_out=16'h8a00;
17'h13d65:	data_out=16'h89e9;
17'h13d66:	data_out=16'ha00;
17'h13d67:	data_out=16'ha00;
17'h13d68:	data_out=16'h5f3;
17'h13d69:	data_out=16'h89fd;
17'h13d6a:	data_out=16'h88c;
17'h13d6b:	data_out=16'ha00;
17'h13d6c:	data_out=16'h81c3;
17'h13d6d:	data_out=16'h89a1;
17'h13d6e:	data_out=16'h889;
17'h13d6f:	data_out=16'ha00;
17'h13d70:	data_out=16'h815;
17'h13d71:	data_out=16'h8914;
17'h13d72:	data_out=16'h4ef;
17'h13d73:	data_out=16'h9fe;
17'h13d74:	data_out=16'h9e1;
17'h13d75:	data_out=16'h9ff;
17'h13d76:	data_out=16'h9e0;
17'h13d77:	data_out=16'h89e0;
17'h13d78:	data_out=16'h89f3;
17'h13d79:	data_out=16'h89c2;
17'h13d7a:	data_out=16'h89b1;
17'h13d7b:	data_out=16'h490;
17'h13d7c:	data_out=16'h84de;
17'h13d7d:	data_out=16'h414;
17'h13d7e:	data_out=16'h89f7;
17'h13d7f:	data_out=16'h9ff;
17'h13d80:	data_out=16'h895a;
17'h13d81:	data_out=16'h8906;
17'h13d82:	data_out=16'h89db;
17'h13d83:	data_out=16'h89c7;
17'h13d84:	data_out=16'ha00;
17'h13d85:	data_out=16'ha00;
17'h13d86:	data_out=16'h89e6;
17'h13d87:	data_out=16'h89ec;
17'h13d88:	data_out=16'h89f4;
17'h13d89:	data_out=16'h89e9;
17'h13d8a:	data_out=16'h9f5;
17'h13d8b:	data_out=16'h89ee;
17'h13d8c:	data_out=16'h89fd;
17'h13d8d:	data_out=16'h89bb;
17'h13d8e:	data_out=16'h9ff;
17'h13d8f:	data_out=16'h89d7;
17'h13d90:	data_out=16'h89e8;
17'h13d91:	data_out=16'h89fd;
17'h13d92:	data_out=16'h89f0;
17'h13d93:	data_out=16'h8995;
17'h13d94:	data_out=16'h89d2;
17'h13d95:	data_out=16'ha00;
17'h13d96:	data_out=16'h869d;
17'h13d97:	data_out=16'h89d3;
17'h13d98:	data_out=16'h961;
17'h13d99:	data_out=16'h9f0;
17'h13d9a:	data_out=16'ha00;
17'h13d9b:	data_out=16'h89e4;
17'h13d9c:	data_out=16'h89c7;
17'h13d9d:	data_out=16'h8a00;
17'h13d9e:	data_out=16'h8963;
17'h13d9f:	data_out=16'h57a;
17'h13da0:	data_out=16'h87cd;
17'h13da1:	data_out=16'h9ff;
17'h13da2:	data_out=16'h8648;
17'h13da3:	data_out=16'h192;
17'h13da4:	data_out=16'h197;
17'h13da5:	data_out=16'h89a1;
17'h13da6:	data_out=16'h89fd;
17'h13da7:	data_out=16'h89b9;
17'h13da8:	data_out=16'ha00;
17'h13da9:	data_out=16'h53a;
17'h13daa:	data_out=16'h89f0;
17'h13dab:	data_out=16'h9d8;
17'h13dac:	data_out=16'h38a;
17'h13dad:	data_out=16'h8a00;
17'h13dae:	data_out=16'h89f2;
17'h13daf:	data_out=16'h89cb;
17'h13db0:	data_out=16'ha00;
17'h13db1:	data_out=16'h823b;
17'h13db2:	data_out=16'h8fd;
17'h13db3:	data_out=16'h89b3;
17'h13db4:	data_out=16'h89fe;
17'h13db5:	data_out=16'h9f5;
17'h13db6:	data_out=16'h89ed;
17'h13db7:	data_out=16'h89e7;
17'h13db8:	data_out=16'h89fd;
17'h13db9:	data_out=16'h89ac;
17'h13dba:	data_out=16'h89ab;
17'h13dbb:	data_out=16'h8b6;
17'h13dbc:	data_out=16'h8747;
17'h13dbd:	data_out=16'h8503;
17'h13dbe:	data_out=16'ha00;
17'h13dbf:	data_out=16'ha00;
17'h13dc0:	data_out=16'h8332;
17'h13dc1:	data_out=16'h89bd;
17'h13dc2:	data_out=16'h8a00;
17'h13dc3:	data_out=16'h824a;
17'h13dc4:	data_out=16'ha00;
17'h13dc5:	data_out=16'ha00;
17'h13dc6:	data_out=16'h89e4;
17'h13dc7:	data_out=16'h89f4;
17'h13dc8:	data_out=16'h89f1;
17'h13dc9:	data_out=16'h862c;
17'h13dca:	data_out=16'h89b0;
17'h13dcb:	data_out=16'h8a00;
17'h13dcc:	data_out=16'h89e8;
17'h13dcd:	data_out=16'h469;
17'h13dce:	data_out=16'h89fc;
17'h13dcf:	data_out=16'h89fd;
17'h13dd0:	data_out=16'hd3;
17'h13dd1:	data_out=16'h9ff;
17'h13dd2:	data_out=16'h82b;
17'h13dd3:	data_out=16'h89df;
17'h13dd4:	data_out=16'h897f;
17'h13dd5:	data_out=16'h899d;
17'h13dd6:	data_out=16'h9db;
17'h13dd7:	data_out=16'ha00;
17'h13dd8:	data_out=16'h187;
17'h13dd9:	data_out=16'h8e2;
17'h13dda:	data_out=16'h89e7;
17'h13ddb:	data_out=16'h9fa;
17'h13ddc:	data_out=16'h88d6;
17'h13ddd:	data_out=16'h88e3;
17'h13dde:	data_out=16'h89ee;
17'h13ddf:	data_out=16'h89da;
17'h13de0:	data_out=16'h8a00;
17'h13de1:	data_out=16'ha00;
17'h13de2:	data_out=16'h89f7;
17'h13de3:	data_out=16'h89c9;
17'h13de4:	data_out=16'h8a00;
17'h13de5:	data_out=16'h89ec;
17'h13de6:	data_out=16'ha00;
17'h13de7:	data_out=16'ha00;
17'h13de8:	data_out=16'h9ff;
17'h13de9:	data_out=16'h89f9;
17'h13dea:	data_out=16'h9ff;
17'h13deb:	data_out=16'h9c3;
17'h13dec:	data_out=16'h87e2;
17'h13ded:	data_out=16'h89c6;
17'h13dee:	data_out=16'h9ff;
17'h13def:	data_out=16'h61b;
17'h13df0:	data_out=16'h9ff;
17'h13df1:	data_out=16'h8951;
17'h13df2:	data_out=16'h9ab;
17'h13df3:	data_out=16'h9fd;
17'h13df4:	data_out=16'h9eb;
17'h13df5:	data_out=16'ha00;
17'h13df6:	data_out=16'h9f5;
17'h13df7:	data_out=16'h89f2;
17'h13df8:	data_out=16'h8836;
17'h13df9:	data_out=16'h86ae;
17'h13dfa:	data_out=16'h89cf;
17'h13dfb:	data_out=16'ha00;
17'h13dfc:	data_out=16'h7a2;
17'h13dfd:	data_out=16'ha00;
17'h13dfe:	data_out=16'h89fb;
17'h13dff:	data_out=16'ha00;
17'h13e00:	data_out=16'h8773;
17'h13e01:	data_out=16'h89fe;
17'h13e02:	data_out=16'h89ee;
17'h13e03:	data_out=16'h89a2;
17'h13e04:	data_out=16'ha00;
17'h13e05:	data_out=16'ha00;
17'h13e06:	data_out=16'h89fc;
17'h13e07:	data_out=16'h89fa;
17'h13e08:	data_out=16'h89f3;
17'h13e09:	data_out=16'h89f7;
17'h13e0a:	data_out=16'h9f7;
17'h13e0b:	data_out=16'h89f3;
17'h13e0c:	data_out=16'h89fc;
17'h13e0d:	data_out=16'h89a4;
17'h13e0e:	data_out=16'ha00;
17'h13e0f:	data_out=16'h89f2;
17'h13e10:	data_out=16'h89c5;
17'h13e11:	data_out=16'h8a00;
17'h13e12:	data_out=16'h89f4;
17'h13e13:	data_out=16'h890a;
17'h13e14:	data_out=16'h8956;
17'h13e15:	data_out=16'ha00;
17'h13e16:	data_out=16'h521;
17'h13e17:	data_out=16'h89eb;
17'h13e18:	data_out=16'h9fd;
17'h13e19:	data_out=16'h9ee;
17'h13e1a:	data_out=16'ha00;
17'h13e1b:	data_out=16'h89c3;
17'h13e1c:	data_out=16'h73e;
17'h13e1d:	data_out=16'h8a00;
17'h13e1e:	data_out=16'h899f;
17'h13e1f:	data_out=16'h874;
17'h13e20:	data_out=16'h84d0;
17'h13e21:	data_out=16'ha00;
17'h13e22:	data_out=16'ha00;
17'h13e23:	data_out=16'h9fb;
17'h13e24:	data_out=16'h9fb;
17'h13e25:	data_out=16'h83ea;
17'h13e26:	data_out=16'h89eb;
17'h13e27:	data_out=16'h89ed;
17'h13e28:	data_out=16'ha00;
17'h13e29:	data_out=16'h9ff;
17'h13e2a:	data_out=16'h89f6;
17'h13e2b:	data_out=16'h9da;
17'h13e2c:	data_out=16'ha00;
17'h13e2d:	data_out=16'h8a00;
17'h13e2e:	data_out=16'h89fc;
17'h13e2f:	data_out=16'h89ee;
17'h13e30:	data_out=16'h8445;
17'h13e31:	data_out=16'h8734;
17'h13e32:	data_out=16'h893d;
17'h13e33:	data_out=16'h895a;
17'h13e34:	data_out=16'h8a00;
17'h13e35:	data_out=16'h9ea;
17'h13e36:	data_out=16'h89f0;
17'h13e37:	data_out=16'h89f5;
17'h13e38:	data_out=16'h89ff;
17'h13e39:	data_out=16'h8937;
17'h13e3a:	data_out=16'h89bc;
17'h13e3b:	data_out=16'h784;
17'h13e3c:	data_out=16'h86b6;
17'h13e3d:	data_out=16'ha00;
17'h13e3e:	data_out=16'ha00;
17'h13e3f:	data_out=16'ha00;
17'h13e40:	data_out=16'h858c;
17'h13e41:	data_out=16'h89b8;
17'h13e42:	data_out=16'h89ff;
17'h13e43:	data_out=16'h82bb;
17'h13e44:	data_out=16'ha00;
17'h13e45:	data_out=16'ha00;
17'h13e46:	data_out=16'h89e6;
17'h13e47:	data_out=16'h89f9;
17'h13e48:	data_out=16'h89f9;
17'h13e49:	data_out=16'h4d2;
17'h13e4a:	data_out=16'h89f8;
17'h13e4b:	data_out=16'h89fe;
17'h13e4c:	data_out=16'h89ea;
17'h13e4d:	data_out=16'ha00;
17'h13e4e:	data_out=16'h89fb;
17'h13e4f:	data_out=16'h89fd;
17'h13e50:	data_out=16'h879;
17'h13e51:	data_out=16'ha00;
17'h13e52:	data_out=16'h92d;
17'h13e53:	data_out=16'h89f3;
17'h13e54:	data_out=16'h89e0;
17'h13e55:	data_out=16'h5e6;
17'h13e56:	data_out=16'h9f8;
17'h13e57:	data_out=16'ha00;
17'h13e58:	data_out=16'h8df;
17'h13e59:	data_out=16'h9e1;
17'h13e5a:	data_out=16'h89f8;
17'h13e5b:	data_out=16'ha00;
17'h13e5c:	data_out=16'h8906;
17'h13e5d:	data_out=16'h89ca;
17'h13e5e:	data_out=16'h89f8;
17'h13e5f:	data_out=16'h89f7;
17'h13e60:	data_out=16'h89fd;
17'h13e61:	data_out=16'h9ff;
17'h13e62:	data_out=16'h89f8;
17'h13e63:	data_out=16'h89da;
17'h13e64:	data_out=16'h8a00;
17'h13e65:	data_out=16'h89fe;
17'h13e66:	data_out=16'h9ff;
17'h13e67:	data_out=16'ha00;
17'h13e68:	data_out=16'ha00;
17'h13e69:	data_out=16'h89f4;
17'h13e6a:	data_out=16'ha00;
17'h13e6b:	data_out=16'h9fb;
17'h13e6c:	data_out=16'h8992;
17'h13e6d:	data_out=16'h89d3;
17'h13e6e:	data_out=16'ha00;
17'h13e6f:	data_out=16'h8701;
17'h13e70:	data_out=16'ha00;
17'h13e71:	data_out=16'h89f4;
17'h13e72:	data_out=16'h9e4;
17'h13e73:	data_out=16'h9f7;
17'h13e74:	data_out=16'h8474;
17'h13e75:	data_out=16'ha00;
17'h13e76:	data_out=16'h9f8;
17'h13e77:	data_out=16'h89f4;
17'h13e78:	data_out=16'h8223;
17'h13e79:	data_out=16'h82c2;
17'h13e7a:	data_out=16'h89cf;
17'h13e7b:	data_out=16'ha00;
17'h13e7c:	data_out=16'h74e;
17'h13e7d:	data_out=16'ha00;
17'h13e7e:	data_out=16'h89fc;
17'h13e7f:	data_out=16'ha00;
17'h13e80:	data_out=16'h88f;
17'h13e81:	data_out=16'h8a00;
17'h13e82:	data_out=16'h89c9;
17'h13e83:	data_out=16'h89aa;
17'h13e84:	data_out=16'ha00;
17'h13e85:	data_out=16'h445;
17'h13e86:	data_out=16'h89fe;
17'h13e87:	data_out=16'h89fe;
17'h13e88:	data_out=16'h89f7;
17'h13e89:	data_out=16'h79;
17'h13e8a:	data_out=16'h9fc;
17'h13e8b:	data_out=16'h89f9;
17'h13e8c:	data_out=16'h89fe;
17'h13e8d:	data_out=16'h89b8;
17'h13e8e:	data_out=16'ha00;
17'h13e8f:	data_out=16'h89fa;
17'h13e90:	data_out=16'h8010;
17'h13e91:	data_out=16'h824e;
17'h13e92:	data_out=16'h89fb;
17'h13e93:	data_out=16'h8933;
17'h13e94:	data_out=16'h8996;
17'h13e95:	data_out=16'ha00;
17'h13e96:	data_out=16'h6bb;
17'h13e97:	data_out=16'h89f6;
17'h13e98:	data_out=16'ha00;
17'h13e99:	data_out=16'h3c4;
17'h13e9a:	data_out=16'h56f;
17'h13e9b:	data_out=16'h89ba;
17'h13e9c:	data_out=16'h9ee;
17'h13e9d:	data_out=16'h8a00;
17'h13e9e:	data_out=16'h899c;
17'h13e9f:	data_out=16'h9fd;
17'h13ea0:	data_out=16'h9de;
17'h13ea1:	data_out=16'ha00;
17'h13ea2:	data_out=16'ha00;
17'h13ea3:	data_out=16'ha00;
17'h13ea4:	data_out=16'ha00;
17'h13ea5:	data_out=16'ha00;
17'h13ea6:	data_out=16'h89c5;
17'h13ea7:	data_out=16'h89f6;
17'h13ea8:	data_out=16'ha00;
17'h13ea9:	data_out=16'h887;
17'h13eaa:	data_out=16'h89fb;
17'h13eab:	data_out=16'h9f2;
17'h13eac:	data_out=16'h9ff;
17'h13ead:	data_out=16'h8a00;
17'h13eae:	data_out=16'h89fe;
17'h13eaf:	data_out=16'h89fb;
17'h13eb0:	data_out=16'h87c3;
17'h13eb1:	data_out=16'h89ce;
17'h13eb2:	data_out=16'h8976;
17'h13eb3:	data_out=16'h27e;
17'h13eb4:	data_out=16'h8a00;
17'h13eb5:	data_out=16'h9e4;
17'h13eb6:	data_out=16'h89f7;
17'h13eb7:	data_out=16'h89c8;
17'h13eb8:	data_out=16'h809b;
17'h13eb9:	data_out=16'h6e;
17'h13eba:	data_out=16'h81fd;
17'h13ebb:	data_out=16'h679;
17'h13ebc:	data_out=16'h8880;
17'h13ebd:	data_out=16'ha00;
17'h13ebe:	data_out=16'ha00;
17'h13ebf:	data_out=16'h509;
17'h13ec0:	data_out=16'h9e6;
17'h13ec1:	data_out=16'h89a0;
17'h13ec2:	data_out=16'h89fe;
17'h13ec3:	data_out=16'h86fb;
17'h13ec4:	data_out=16'h9e6;
17'h13ec5:	data_out=16'ha00;
17'h13ec6:	data_out=16'h89e3;
17'h13ec7:	data_out=16'h89fc;
17'h13ec8:	data_out=16'h89fd;
17'h13ec9:	data_out=16'ha00;
17'h13eca:	data_out=16'h89fd;
17'h13ecb:	data_out=16'h89fe;
17'h13ecc:	data_out=16'h889e;
17'h13ecd:	data_out=16'ha00;
17'h13ece:	data_out=16'h89fe;
17'h13ecf:	data_out=16'h160;
17'h13ed0:	data_out=16'h9a8;
17'h13ed1:	data_out=16'ha00;
17'h13ed2:	data_out=16'h9ff;
17'h13ed3:	data_out=16'h89f8;
17'h13ed4:	data_out=16'h89ea;
17'h13ed5:	data_out=16'h70c;
17'h13ed6:	data_out=16'ha00;
17'h13ed7:	data_out=16'ha00;
17'h13ed8:	data_out=16'h9df;
17'h13ed9:	data_out=16'h9fd;
17'h13eda:	data_out=16'h89fc;
17'h13edb:	data_out=16'h9fa;
17'h13edc:	data_out=16'h89d1;
17'h13edd:	data_out=16'h89d9;
17'h13ede:	data_out=16'h89fc;
17'h13edf:	data_out=16'h87f0;
17'h13ee0:	data_out=16'h89fa;
17'h13ee1:	data_out=16'h9f2;
17'h13ee2:	data_out=16'h89f9;
17'h13ee3:	data_out=16'h8743;
17'h13ee4:	data_out=16'h89f5;
17'h13ee5:	data_out=16'h89ff;
17'h13ee6:	data_out=16'h8e;
17'h13ee7:	data_out=16'ha00;
17'h13ee8:	data_out=16'ha00;
17'h13ee9:	data_out=16'h89f6;
17'h13eea:	data_out=16'ha00;
17'h13eeb:	data_out=16'h9eb;
17'h13eec:	data_out=16'h88d4;
17'h13eed:	data_out=16'h84e0;
17'h13eee:	data_out=16'ha00;
17'h13eef:	data_out=16'h89df;
17'h13ef0:	data_out=16'ha00;
17'h13ef1:	data_out=16'h89fc;
17'h13ef2:	data_out=16'h9fc;
17'h13ef3:	data_out=16'h9fb;
17'h13ef4:	data_out=16'h87a6;
17'h13ef5:	data_out=16'h9c8;
17'h13ef6:	data_out=16'ha00;
17'h13ef7:	data_out=16'h2bb;
17'h13ef8:	data_out=16'h867c;
17'h13ef9:	data_out=16'h82bf;
17'h13efa:	data_out=16'h89de;
17'h13efb:	data_out=16'ha00;
17'h13efc:	data_out=16'h91e;
17'h13efd:	data_out=16'h470;
17'h13efe:	data_out=16'h163;
17'h13eff:	data_out=16'ha00;
17'h13f00:	data_out=16'h9fb;
17'h13f01:	data_out=16'h8a00;
17'h13f02:	data_out=16'h89d1;
17'h13f03:	data_out=16'h89cc;
17'h13f04:	data_out=16'ha00;
17'h13f05:	data_out=16'h819a;
17'h13f06:	data_out=16'h89ff;
17'h13f07:	data_out=16'h8a00;
17'h13f08:	data_out=16'h89df;
17'h13f09:	data_out=16'h728;
17'h13f0a:	data_out=16'h9f6;
17'h13f0b:	data_out=16'h89c2;
17'h13f0c:	data_out=16'h89ff;
17'h13f0d:	data_out=16'h89f5;
17'h13f0e:	data_out=16'ha00;
17'h13f0f:	data_out=16'h89fe;
17'h13f10:	data_out=16'ha00;
17'h13f11:	data_out=16'h80a;
17'h13f12:	data_out=16'h89fc;
17'h13f13:	data_out=16'h89cb;
17'h13f14:	data_out=16'h826d;
17'h13f15:	data_out=16'ha00;
17'h13f16:	data_out=16'h815e;
17'h13f17:	data_out=16'h89fc;
17'h13f18:	data_out=16'ha00;
17'h13f19:	data_out=16'h5e2;
17'h13f1a:	data_out=16'h375;
17'h13f1b:	data_out=16'h89b5;
17'h13f1c:	data_out=16'h9e9;
17'h13f1d:	data_out=16'h8a00;
17'h13f1e:	data_out=16'h8923;
17'h13f1f:	data_out=16'h893;
17'h13f20:	data_out=16'h9f5;
17'h13f21:	data_out=16'ha00;
17'h13f22:	data_out=16'ha00;
17'h13f23:	data_out=16'ha00;
17'h13f24:	data_out=16'ha00;
17'h13f25:	data_out=16'ha00;
17'h13f26:	data_out=16'h9e9;
17'h13f27:	data_out=16'h897e;
17'h13f28:	data_out=16'ha00;
17'h13f29:	data_out=16'h36e;
17'h13f2a:	data_out=16'h89ff;
17'h13f2b:	data_out=16'ha00;
17'h13f2c:	data_out=16'h92e;
17'h13f2d:	data_out=16'h81aa;
17'h13f2e:	data_out=16'h89ff;
17'h13f2f:	data_out=16'h89fe;
17'h13f30:	data_out=16'h89f0;
17'h13f31:	data_out=16'h89df;
17'h13f32:	data_out=16'h8a00;
17'h13f33:	data_out=16'h9a7;
17'h13f34:	data_out=16'h8a00;
17'h13f35:	data_out=16'ha00;
17'h13f36:	data_out=16'h89cc;
17'h13f37:	data_out=16'h89d8;
17'h13f38:	data_out=16'h88c;
17'h13f39:	data_out=16'h9fe;
17'h13f3a:	data_out=16'ha00;
17'h13f3b:	data_out=16'h4dd;
17'h13f3c:	data_out=16'h88a8;
17'h13f3d:	data_out=16'ha00;
17'h13f3e:	data_out=16'ha00;
17'h13f3f:	data_out=16'h80ef;
17'h13f40:	data_out=16'h9f1;
17'h13f41:	data_out=16'h8998;
17'h13f42:	data_out=16'h89fe;
17'h13f43:	data_out=16'h89da;
17'h13f44:	data_out=16'h9fc;
17'h13f45:	data_out=16'ha00;
17'h13f46:	data_out=16'h9f6;
17'h13f47:	data_out=16'h1ac;
17'h13f48:	data_out=16'h89ff;
17'h13f49:	data_out=16'ha00;
17'h13f4a:	data_out=16'h89ff;
17'h13f4b:	data_out=16'h89ff;
17'h13f4c:	data_out=16'h88b2;
17'h13f4d:	data_out=16'ha00;
17'h13f4e:	data_out=16'h89f5;
17'h13f4f:	data_out=16'h6d1;
17'h13f50:	data_out=16'h852;
17'h13f51:	data_out=16'h4dc;
17'h13f52:	data_out=16'ha00;
17'h13f53:	data_out=16'h89ef;
17'h13f54:	data_out=16'h898;
17'h13f55:	data_out=16'h90a;
17'h13f56:	data_out=16'ha00;
17'h13f57:	data_out=16'ha00;
17'h13f58:	data_out=16'h9e9;
17'h13f59:	data_out=16'h9fb;
17'h13f5a:	data_out=16'h89fa;
17'h13f5b:	data_out=16'ha00;
17'h13f5c:	data_out=16'h89fd;
17'h13f5d:	data_out=16'h89d0;
17'h13f5e:	data_out=16'h89fe;
17'h13f5f:	data_out=16'h41;
17'h13f60:	data_out=16'h89d1;
17'h13f61:	data_out=16'h9f3;
17'h13f62:	data_out=16'h89fb;
17'h13f63:	data_out=16'h66b;
17'h13f64:	data_out=16'h68f;
17'h13f65:	data_out=16'h8a00;
17'h13f66:	data_out=16'h22c;
17'h13f67:	data_out=16'ha00;
17'h13f68:	data_out=16'ha00;
17'h13f69:	data_out=16'h89e0;
17'h13f6a:	data_out=16'ha00;
17'h13f6b:	data_out=16'h9e4;
17'h13f6c:	data_out=16'h886d;
17'h13f6d:	data_out=16'h78d;
17'h13f6e:	data_out=16'ha00;
17'h13f6f:	data_out=16'h8a00;
17'h13f70:	data_out=16'ha00;
17'h13f71:	data_out=16'h89ff;
17'h13f72:	data_out=16'h9f1;
17'h13f73:	data_out=16'h98d;
17'h13f74:	data_out=16'h89f1;
17'h13f75:	data_out=16'h8945;
17'h13f76:	data_out=16'ha00;
17'h13f77:	data_out=16'h7f1;
17'h13f78:	data_out=16'h8960;
17'h13f79:	data_out=16'h8505;
17'h13f7a:	data_out=16'h80a9;
17'h13f7b:	data_out=16'ha00;
17'h13f7c:	data_out=16'h9c2;
17'h13f7d:	data_out=16'h82de;
17'h13f7e:	data_out=16'h75c;
17'h13f7f:	data_out=16'ha00;
17'h13f80:	data_out=16'ha00;
17'h13f81:	data_out=16'h89b0;
17'h13f82:	data_out=16'h8035;
17'h13f83:	data_out=16'h9bc;
17'h13f84:	data_out=16'h9fa;
17'h13f85:	data_out=16'h3a6;
17'h13f86:	data_out=16'h8319;
17'h13f87:	data_out=16'h80d4;
17'h13f88:	data_out=16'h8c8;
17'h13f89:	data_out=16'h94e;
17'h13f8a:	data_out=16'h53a;
17'h13f8b:	data_out=16'h820f;
17'h13f8c:	data_out=16'h8a00;
17'h13f8d:	data_out=16'h89f7;
17'h13f8e:	data_out=16'h699;
17'h13f8f:	data_out=16'h8447;
17'h13f90:	data_out=16'ha00;
17'h13f91:	data_out=16'h4f7;
17'h13f92:	data_out=16'h89fd;
17'h13f93:	data_out=16'h1c6;
17'h13f94:	data_out=16'h99f;
17'h13f95:	data_out=16'ha00;
17'h13f96:	data_out=16'h9a2;
17'h13f97:	data_out=16'h89fa;
17'h13f98:	data_out=16'h9ff;
17'h13f99:	data_out=16'h8127;
17'h13f9a:	data_out=16'h736;
17'h13f9b:	data_out=16'h89d1;
17'h13f9c:	data_out=16'h9fd;
17'h13f9d:	data_out=16'h558;
17'h13f9e:	data_out=16'h2bf;
17'h13f9f:	data_out=16'h7d6;
17'h13fa0:	data_out=16'h9f5;
17'h13fa1:	data_out=16'h663;
17'h13fa2:	data_out=16'ha00;
17'h13fa3:	data_out=16'ha00;
17'h13fa4:	data_out=16'ha00;
17'h13fa5:	data_out=16'ha00;
17'h13fa6:	data_out=16'h9fe;
17'h13fa7:	data_out=16'h5fa;
17'h13fa8:	data_out=16'h683;
17'h13fa9:	data_out=16'ha00;
17'h13faa:	data_out=16'h8a00;
17'h13fab:	data_out=16'h9fe;
17'h13fac:	data_out=16'h9fa;
17'h13fad:	data_out=16'h80fc;
17'h13fae:	data_out=16'h84ae;
17'h13faf:	data_out=16'h4d0;
17'h13fb0:	data_out=16'h89d2;
17'h13fb1:	data_out=16'h89f8;
17'h13fb2:	data_out=16'h89ff;
17'h13fb3:	data_out=16'h9f4;
17'h13fb4:	data_out=16'h80bb;
17'h13fb5:	data_out=16'h30a;
17'h13fb6:	data_out=16'h746;
17'h13fb7:	data_out=16'h821c;
17'h13fb8:	data_out=16'h825;
17'h13fb9:	data_out=16'h9fc;
17'h13fba:	data_out=16'ha00;
17'h13fbb:	data_out=16'h536;
17'h13fbc:	data_out=16'h8941;
17'h13fbd:	data_out=16'ha00;
17'h13fbe:	data_out=16'h685;
17'h13fbf:	data_out=16'h3f1;
17'h13fc0:	data_out=16'h9f2;
17'h13fc1:	data_out=16'h28c;
17'h13fc2:	data_out=16'h89fe;
17'h13fc3:	data_out=16'h813d;
17'h13fc4:	data_out=16'h9f2;
17'h13fc5:	data_out=16'ha00;
17'h13fc6:	data_out=16'ha00;
17'h13fc7:	data_out=16'h9f7;
17'h13fc8:	data_out=16'h8a00;
17'h13fc9:	data_out=16'ha00;
17'h13fca:	data_out=16'h8a00;
17'h13fcb:	data_out=16'h89ff;
17'h13fcc:	data_out=16'h86bd;
17'h13fcd:	data_out=16'ha00;
17'h13fce:	data_out=16'h89f9;
17'h13fcf:	data_out=16'h556;
17'h13fd0:	data_out=16'h9a6;
17'h13fd1:	data_out=16'h9c3;
17'h13fd2:	data_out=16'ha00;
17'h13fd3:	data_out=16'h89ff;
17'h13fd4:	data_out=16'h9f2;
17'h13fd5:	data_out=16'h930;
17'h13fd6:	data_out=16'ha00;
17'h13fd7:	data_out=16'ha00;
17'h13fd8:	data_out=16'h9f9;
17'h13fd9:	data_out=16'h9f5;
17'h13fda:	data_out=16'h89fd;
17'h13fdb:	data_out=16'h9f7;
17'h13fdc:	data_out=16'h8a00;
17'h13fdd:	data_out=16'h8478;
17'h13fde:	data_out=16'h410;
17'h13fdf:	data_out=16'h219;
17'h13fe0:	data_out=16'h995;
17'h13fe1:	data_out=16'h90c;
17'h13fe2:	data_out=16'h89f8;
17'h13fe3:	data_out=16'h8fa;
17'h13fe4:	data_out=16'ha00;
17'h13fe5:	data_out=16'h89ff;
17'h13fe6:	data_out=16'h820e;
17'h13fe7:	data_out=16'h9f2;
17'h13fe8:	data_out=16'h66e;
17'h13fe9:	data_out=16'h5da;
17'h13fea:	data_out=16'h67e;
17'h13feb:	data_out=16'h9ed;
17'h13fec:	data_out=16'h8007;
17'h13fed:	data_out=16'h949;
17'h13fee:	data_out=16'h67c;
17'h13fef:	data_out=16'h8a00;
17'h13ff0:	data_out=16'h6a2;
17'h13ff1:	data_out=16'h8a00;
17'h13ff2:	data_out=16'h9f2;
17'h13ff3:	data_out=16'h768;
17'h13ff4:	data_out=16'h89bf;
17'h13ff5:	data_out=16'h8a00;
17'h13ff6:	data_out=16'ha00;
17'h13ff7:	data_out=16'h9a4;
17'h13ff8:	data_out=16'h89ab;
17'h13ff9:	data_out=16'h86f9;
17'h13ffa:	data_out=16'h8ea;
17'h13ffb:	data_out=16'h68e;
17'h13ffc:	data_out=16'h522;
17'h13ffd:	data_out=16'h801c;
17'h13ffe:	data_out=16'h9be;
17'h13fff:	data_out=16'ha00;
17'h14000:	data_out=16'h9fe;
17'h14001:	data_out=16'h50;
17'h14002:	data_out=16'h168;
17'h14003:	data_out=16'h9fb;
17'h14004:	data_out=16'h9ff;
17'h14005:	data_out=16'h45d;
17'h14006:	data_out=16'h26c;
17'h14007:	data_out=16'h5ef;
17'h14008:	data_out=16'h988;
17'h14009:	data_out=16'ha00;
17'h1400a:	data_out=16'h223;
17'h1400b:	data_out=16'h3ff;
17'h1400c:	data_out=16'h8a00;
17'h1400d:	data_out=16'h24;
17'h1400e:	data_out=16'h362;
17'h1400f:	data_out=16'h52;
17'h14010:	data_out=16'ha00;
17'h14011:	data_out=16'h320;
17'h14012:	data_out=16'h8201;
17'h14013:	data_out=16'h9fe;
17'h14014:	data_out=16'h9fa;
17'h14015:	data_out=16'ha00;
17'h14016:	data_out=16'h9fc;
17'h14017:	data_out=16'h31a;
17'h14018:	data_out=16'h622;
17'h14019:	data_out=16'h8194;
17'h1401a:	data_out=16'h3ea;
17'h1401b:	data_out=16'h888f;
17'h1401c:	data_out=16'h9ff;
17'h1401d:	data_out=16'h69f;
17'h1401e:	data_out=16'h956;
17'h1401f:	data_out=16'h8ff;
17'h14020:	data_out=16'h9fc;
17'h14021:	data_out=16'h351;
17'h14022:	data_out=16'ha00;
17'h14023:	data_out=16'h3c;
17'h14024:	data_out=16'h41;
17'h14025:	data_out=16'ha00;
17'h14026:	data_out=16'h9fb;
17'h14027:	data_out=16'h853;
17'h14028:	data_out=16'h34d;
17'h14029:	data_out=16'ha00;
17'h1402a:	data_out=16'h157;
17'h1402b:	data_out=16'h955;
17'h1402c:	data_out=16'h9fd;
17'h1402d:	data_out=16'h9fe;
17'h1402e:	data_out=16'h3f2;
17'h1402f:	data_out=16'h9de;
17'h14030:	data_out=16'h89f9;
17'h14031:	data_out=16'h8775;
17'h14032:	data_out=16'h8a00;
17'h14033:	data_out=16'h9ff;
17'h14034:	data_out=16'h630;
17'h14035:	data_out=16'h835b;
17'h14036:	data_out=16'h96b;
17'h14037:	data_out=16'h5d;
17'h14038:	data_out=16'h533;
17'h14039:	data_out=16'ha00;
17'h1403a:	data_out=16'ha00;
17'h1403b:	data_out=16'h64c;
17'h1403c:	data_out=16'h804e;
17'h1403d:	data_out=16'ha00;
17'h1403e:	data_out=16'h34c;
17'h1403f:	data_out=16'h49c;
17'h14040:	data_out=16'h9f9;
17'h14041:	data_out=16'h596;
17'h14042:	data_out=16'h89ee;
17'h14043:	data_out=16'h28c;
17'h14044:	data_out=16'h9f7;
17'h14045:	data_out=16'ha00;
17'h14046:	data_out=16'h7e3;
17'h14047:	data_out=16'ha00;
17'h14048:	data_out=16'h80;
17'h14049:	data_out=16'ha00;
17'h1404a:	data_out=16'h8037;
17'h1404b:	data_out=16'h89ff;
17'h1404c:	data_out=16'h46e;
17'h1404d:	data_out=16'ha00;
17'h1404e:	data_out=16'h82c0;
17'h1404f:	data_out=16'h7ea;
17'h14050:	data_out=16'h9fb;
17'h14051:	data_out=16'h83a;
17'h14052:	data_out=16'h4af;
17'h14053:	data_out=16'h8a00;
17'h14054:	data_out=16'h9fa;
17'h14055:	data_out=16'h9be;
17'h14056:	data_out=16'h9fe;
17'h14057:	data_out=16'ha00;
17'h14058:	data_out=16'h9f9;
17'h14059:	data_out=16'h9fb;
17'h1405a:	data_out=16'h89ff;
17'h1405b:	data_out=16'h8a2;
17'h1405c:	data_out=16'h8598;
17'h1405d:	data_out=16'h511;
17'h1405e:	data_out=16'h9c6;
17'h1405f:	data_out=16'h38a;
17'h14060:	data_out=16'h91c;
17'h14061:	data_out=16'h8f1;
17'h14062:	data_out=16'h892c;
17'h14063:	data_out=16'h9e9;
17'h14064:	data_out=16'ha00;
17'h14065:	data_out=16'h3e1;
17'h14066:	data_out=16'h8017;
17'h14067:	data_out=16'h8e6;
17'h14068:	data_out=16'h352;
17'h14069:	data_out=16'h61a;
17'h1406a:	data_out=16'h373;
17'h1406b:	data_out=16'h9fa;
17'h1406c:	data_out=16'h81f6;
17'h1406d:	data_out=16'h9fc;
17'h1406e:	data_out=16'h372;
17'h1406f:	data_out=16'h8256;
17'h14070:	data_out=16'h367;
17'h14071:	data_out=16'h8a00;
17'h14072:	data_out=16'h9fb;
17'h14073:	data_out=16'h971;
17'h14074:	data_out=16'h89ef;
17'h14075:	data_out=16'h8a00;
17'h14076:	data_out=16'h8b2;
17'h14077:	data_out=16'h9fe;
17'h14078:	data_out=16'h8085;
17'h14079:	data_out=16'h206;
17'h1407a:	data_out=16'h9dc;
17'h1407b:	data_out=16'h34b;
17'h1407c:	data_out=16'h22b;
17'h1407d:	data_out=16'he5;
17'h1407e:	data_out=16'ha00;
17'h1407f:	data_out=16'ha00;
17'h14080:	data_out=16'ha00;
17'h14081:	data_out=16'h2ba;
17'h14082:	data_out=16'h808e;
17'h14083:	data_out=16'h49b;
17'h14084:	data_out=16'h34d;
17'h14085:	data_out=16'h32d;
17'h14086:	data_out=16'h8389;
17'h14087:	data_out=16'h150;
17'h14088:	data_out=16'h468;
17'h14089:	data_out=16'h92d;
17'h1408a:	data_out=16'h3c1;
17'h1408b:	data_out=16'h86cf;
17'h1408c:	data_out=16'h879a;
17'h1408d:	data_out=16'h184;
17'h1408e:	data_out=16'ha0;
17'h1408f:	data_out=16'h8066;
17'h14090:	data_out=16'h6d1;
17'h14091:	data_out=16'h15;
17'h14092:	data_out=16'h87bc;
17'h14093:	data_out=16'h2c4;
17'h14094:	data_out=16'hf7;
17'h14095:	data_out=16'h644;
17'h14096:	data_out=16'h630;
17'h14097:	data_out=16'h827c;
17'h14098:	data_out=16'h340;
17'h14099:	data_out=16'h80dc;
17'h1409a:	data_out=16'hed;
17'h1409b:	data_out=16'h8669;
17'h1409c:	data_out=16'h654;
17'h1409d:	data_out=16'h13c;
17'h1409e:	data_out=16'h169;
17'h1409f:	data_out=16'h397;
17'h140a0:	data_out=16'h9ff;
17'h140a1:	data_out=16'h99;
17'h140a2:	data_out=16'h749;
17'h140a3:	data_out=16'h8191;
17'h140a4:	data_out=16'h818c;
17'h140a5:	data_out=16'h3a1;
17'h140a6:	data_out=16'h308;
17'h140a7:	data_out=16'h15f;
17'h140a8:	data_out=16'hbf;
17'h140a9:	data_out=16'h2a5;
17'h140aa:	data_out=16'h835d;
17'h140ab:	data_out=16'h1a9;
17'h140ac:	data_out=16'h6c2;
17'h140ad:	data_out=16'h80b5;
17'h140ae:	data_out=16'h81c3;
17'h140af:	data_out=16'h298;
17'h140b0:	data_out=16'h8534;
17'h140b1:	data_out=16'h50;
17'h140b2:	data_out=16'h858e;
17'h140b3:	data_out=16'h2f2;
17'h140b4:	data_out=16'h93;
17'h140b5:	data_out=16'h8076;
17'h140b6:	data_out=16'h3fb;
17'h140b7:	data_out=16'h819c;
17'h140b8:	data_out=16'h27e;
17'h140b9:	data_out=16'h3ec;
17'h140ba:	data_out=16'h417;
17'h140bb:	data_out=16'h567;
17'h140bc:	data_out=16'h8349;
17'h140bd:	data_out=16'ha00;
17'h140be:	data_out=16'hbf;
17'h140bf:	data_out=16'h3b8;
17'h140c0:	data_out=16'h56c;
17'h140c1:	data_out=16'h1b8;
17'h140c2:	data_out=16'h880c;
17'h140c3:	data_out=16'h80c0;
17'h140c4:	data_out=16'h777;
17'h140c5:	data_out=16'h652;
17'h140c6:	data_out=16'h8064;
17'h140c7:	data_out=16'h35e;
17'h140c8:	data_out=16'h8384;
17'h140c9:	data_out=16'h40d;
17'h140ca:	data_out=16'h80c6;
17'h140cb:	data_out=16'h8a00;
17'h140cc:	data_out=16'h8231;
17'h140cd:	data_out=16'h77e;
17'h140ce:	data_out=16'h8401;
17'h140cf:	data_out=16'h80d1;
17'h140d0:	data_out=16'h731;
17'h140d1:	data_out=16'h492;
17'h140d2:	data_out=16'he6;
17'h140d3:	data_out=16'h86cc;
17'h140d4:	data_out=16'h73f;
17'h140d5:	data_out=16'h2ce;
17'h140d6:	data_out=16'h55f;
17'h140d7:	data_out=16'h600;
17'h140d8:	data_out=16'h2c2;
17'h140d9:	data_out=16'h5b6;
17'h140da:	data_out=16'h89c2;
17'h140db:	data_out=16'h65b;
17'h140dc:	data_out=16'ha5;
17'h140dd:	data_out=16'h227;
17'h140de:	data_out=16'h2b5;
17'h140df:	data_out=16'h230;
17'h140e0:	data_out=16'h816b;
17'h140e1:	data_out=16'h842;
17'h140e2:	data_out=16'h85ff;
17'h140e3:	data_out=16'h237;
17'h140e4:	data_out=16'h28a;
17'h140e5:	data_out=16'h8356;
17'h140e6:	data_out=16'h8087;
17'h140e7:	data_out=16'h80ff;
17'h140e8:	data_out=16'h9d;
17'h140e9:	data_out=16'h29b;
17'h140ea:	data_out=16'h7c;
17'h140eb:	data_out=16'h629;
17'h140ec:	data_out=16'h3a1;
17'h140ed:	data_out=16'h2c3;
17'h140ee:	data_out=16'h87;
17'h140ef:	data_out=16'h80f7;
17'h140f0:	data_out=16'h98;
17'h140f1:	data_out=16'h8186;
17'h140f2:	data_out=16'h5e7;
17'h140f3:	data_out=16'h663;
17'h140f4:	data_out=16'h8568;
17'h140f5:	data_out=16'h86ce;
17'h140f6:	data_out=16'h184;
17'h140f7:	data_out=16'h6e6;
17'h140f8:	data_out=16'h81c1;
17'h140f9:	data_out=16'h80b2;
17'h140fa:	data_out=16'h160;
17'h140fb:	data_out=16'hcb;
17'h140fc:	data_out=16'h258;
17'h140fd:	data_out=16'h82fb;
17'h140fe:	data_out=16'h998;
17'h140ff:	data_out=16'h726;
17'h14100:	data_out=16'h11d;
17'h14101:	data_out=16'h15a;
17'h14102:	data_out=16'h118;
17'h14103:	data_out=16'h57;
17'h14104:	data_out=16'h100;
17'h14105:	data_out=16'h85;
17'h14106:	data_out=16'h801e;
17'h14107:	data_out=16'hfb;
17'h14108:	data_out=16'h188;
17'h14109:	data_out=16'h74;
17'h1410a:	data_out=16'h14c;
17'h1410b:	data_out=16'h80c0;
17'h1410c:	data_out=16'h153;
17'h1410d:	data_out=16'h65;
17'h1410e:	data_out=16'h2f;
17'h1410f:	data_out=16'h101;
17'h14110:	data_out=16'h6f;
17'h14111:	data_out=16'h99;
17'h14112:	data_out=16'h8012;
17'h14113:	data_out=16'h8014;
17'h14114:	data_out=16'h5b;
17'h14115:	data_out=16'hc5;
17'h14116:	data_out=16'h143;
17'h14117:	data_out=16'h8000;
17'h14118:	data_out=16'hb4;
17'h14119:	data_out=16'h806e;
17'h1411a:	data_out=16'hc5;
17'h1411b:	data_out=16'h8083;
17'h1411c:	data_out=16'h4c;
17'h1411d:	data_out=16'he8;
17'h1411e:	data_out=16'h800a;
17'h1411f:	data_out=16'hd8;
17'h14120:	data_out=16'he3;
17'h14121:	data_out=16'h3a;
17'h14122:	data_out=16'h3;
17'h14123:	data_out=16'h1a0;
17'h14124:	data_out=16'h1a1;
17'h14125:	data_out=16'h60;
17'h14126:	data_out=16'h68;
17'h14127:	data_out=16'hd6;
17'h14128:	data_out=16'h3a;
17'h14129:	data_out=16'h8001;
17'h1412a:	data_out=16'h68;
17'h1412b:	data_out=16'h8005;
17'h1412c:	data_out=16'h14e;
17'h1412d:	data_out=16'h8054;
17'h1412e:	data_out=16'h68;
17'h1412f:	data_out=16'ha0;
17'h14130:	data_out=16'h54;
17'h14131:	data_out=16'h8000;
17'h14132:	data_out=16'h2b;
17'h14133:	data_out=16'h7c;
17'h14134:	data_out=16'h802c;
17'h14135:	data_out=16'h1af;
17'h14136:	data_out=16'h22f;
17'h14137:	data_out=16'h110;
17'h14138:	data_out=16'h16;
17'h14139:	data_out=16'h44;
17'h1413a:	data_out=16'h12c;
17'h1413b:	data_out=16'h186;
17'h1413c:	data_out=16'h82;
17'h1413d:	data_out=16'hd1;
17'h1413e:	data_out=16'h33;
17'h1413f:	data_out=16'h80;
17'h14140:	data_out=16'hee;
17'h14141:	data_out=16'h127;
17'h14142:	data_out=16'h804e;
17'h14143:	data_out=16'h8012;
17'h14144:	data_out=16'h11c;
17'h14145:	data_out=16'h11f;
17'h14146:	data_out=16'h802d;
17'h14147:	data_out=16'hf2;
17'h14148:	data_out=16'h805b;
17'h14149:	data_out=16'h70;
17'h1414a:	data_out=16'hcd;
17'h1414b:	data_out=16'h20;
17'h1414c:	data_out=16'h38;
17'h1414d:	data_out=16'h28;
17'h1414e:	data_out=16'hb2;
17'h1414f:	data_out=16'h56;
17'h14150:	data_out=16'hfe;
17'h14151:	data_out=16'h162;
17'h14152:	data_out=16'h19d;
17'h14153:	data_out=16'h2;
17'h14154:	data_out=16'h137;
17'h14155:	data_out=16'h18c;
17'h14156:	data_out=16'h12e;
17'h14157:	data_out=16'h10e;
17'h14158:	data_out=16'h16f;
17'h14159:	data_out=16'he4;
17'h1415a:	data_out=16'h80d7;
17'h1415b:	data_out=16'h246;
17'h1415c:	data_out=16'hcf;
17'h1415d:	data_out=16'h6a;
17'h1415e:	data_out=16'h5e;
17'h1415f:	data_out=16'h99;
17'h14160:	data_out=16'h4c;
17'h14161:	data_out=16'h197;
17'h14162:	data_out=16'h8046;
17'h14163:	data_out=16'h73;
17'h14164:	data_out=16'h8040;
17'h14165:	data_out=16'h808f;
17'h14166:	data_out=16'h801d;
17'h14167:	data_out=16'h8037;
17'h14168:	data_out=16'h35;
17'h14169:	data_out=16'h1f8;
17'h1416a:	data_out=16'h33;
17'h1416b:	data_out=16'h85;
17'h1416c:	data_out=16'h188;
17'h1416d:	data_out=16'h81;
17'h1416e:	data_out=16'h3d;
17'h1416f:	data_out=16'h8064;
17'h14170:	data_out=16'h3c;
17'h14171:	data_out=16'h131;
17'h14172:	data_out=16'h16;
17'h14173:	data_out=16'h65;
17'h14174:	data_out=16'h55;
17'h14175:	data_out=16'h8006;
17'h14176:	data_out=16'h7;
17'h14177:	data_out=16'hd8;
17'h14178:	data_out=16'h8057;
17'h14179:	data_out=16'h117;
17'h1417a:	data_out=16'h72;
17'h1417b:	data_out=16'h3c;
17'h1417c:	data_out=16'hee;
17'h1417d:	data_out=16'h40;
17'h1417e:	data_out=16'h46;
17'h1417f:	data_out=16'hfd;
17'h14180:	data_out=16'h17;
17'h14181:	data_out=16'h2;
17'h14182:	data_out=16'h13;
17'h14183:	data_out=16'he;
17'h14184:	data_out=16'h9;
17'h14185:	data_out=16'h5;
17'h14186:	data_out=16'he;
17'h14187:	data_out=16'h19;
17'h14188:	data_out=16'he;
17'h14189:	data_out=16'h8;
17'h1418a:	data_out=16'h1f;
17'h1418b:	data_out=16'h6;
17'h1418c:	data_out=16'h8;
17'h1418d:	data_out=16'h12;
17'h1418e:	data_out=16'hc;
17'h1418f:	data_out=16'h11;
17'h14190:	data_out=16'h12;
17'h14191:	data_out=16'h8000;
17'h14192:	data_out=16'h18;
17'h14193:	data_out=16'h11;
17'h14194:	data_out=16'h1d;
17'h14195:	data_out=16'h8001;
17'h14196:	data_out=16'hc;
17'h14197:	data_out=16'h1b;
17'h14198:	data_out=16'hc;
17'h14199:	data_out=16'he;
17'h1419a:	data_out=16'h4;
17'h1419b:	data_out=16'h15;
17'h1419c:	data_out=16'h10;
17'h1419d:	data_out=16'hf;
17'h1419e:	data_out=16'he;
17'h1419f:	data_out=16'h15;
17'h141a0:	data_out=16'h7;
17'h141a1:	data_out=16'h7;
17'h141a2:	data_out=16'hc;
17'h141a3:	data_out=16'ha;
17'h141a4:	data_out=16'hc;
17'h141a5:	data_out=16'hf;
17'h141a6:	data_out=16'h13;
17'h141a7:	data_out=16'hc;
17'h141a8:	data_out=16'h1;
17'h141a9:	data_out=16'hd;
17'h141aa:	data_out=16'hf;
17'h141ab:	data_out=16'h5;
17'h141ac:	data_out=16'h7;
17'h141ad:	data_out=16'h3;
17'h141ae:	data_out=16'h12;
17'h141af:	data_out=16'h13;
17'h141b0:	data_out=16'h7;
17'h141b1:	data_out=16'h7;
17'h141b2:	data_out=16'hb;
17'h141b3:	data_out=16'h1a;
17'h141b4:	data_out=16'h12;
17'h141b5:	data_out=16'h11;
17'h141b6:	data_out=16'hd;
17'h141b7:	data_out=16'h16;
17'h141b8:	data_out=16'h8004;
17'h141b9:	data_out=16'h10;
17'h141ba:	data_out=16'h17;
17'h141bb:	data_out=16'h8;
17'h141bc:	data_out=16'h29;
17'h141bd:	data_out=16'he;
17'h141be:	data_out=16'h1;
17'h141bf:	data_out=16'h3;
17'h141c0:	data_out=16'hd;
17'h141c1:	data_out=16'h12;
17'h141c2:	data_out=16'h1c;
17'h141c3:	data_out=16'h0;
17'h141c4:	data_out=16'h12;
17'h141c5:	data_out=16'h1;
17'h141c6:	data_out=16'ha;
17'h141c7:	data_out=16'h1a;
17'h141c8:	data_out=16'h17;
17'h141c9:	data_out=16'h12;
17'h141ca:	data_out=16'h15;
17'h141cb:	data_out=16'h15;
17'h141cc:	data_out=16'h10;
17'h141cd:	data_out=16'hb;
17'h141ce:	data_out=16'h13;
17'h141cf:	data_out=16'h12;
17'h141d0:	data_out=16'h14;
17'h141d1:	data_out=16'h13;
17'h141d2:	data_out=16'h1;
17'h141d3:	data_out=16'h14;
17'h141d4:	data_out=16'he;
17'h141d5:	data_out=16'h1d;
17'h141d6:	data_out=16'h27;
17'h141d7:	data_out=16'h13;
17'h141d8:	data_out=16'h20;
17'h141d9:	data_out=16'h15;
17'h141da:	data_out=16'h13;
17'h141db:	data_out=16'h8001;
17'h141dc:	data_out=16'h13;
17'h141dd:	data_out=16'h16;
17'h141de:	data_out=16'h10;
17'h141df:	data_out=16'h4;
17'h141e0:	data_out=16'h12;
17'h141e1:	data_out=16'h7;
17'h141e2:	data_out=16'hd;
17'h141e3:	data_out=16'hd;
17'h141e4:	data_out=16'h14;
17'h141e5:	data_out=16'h13;
17'h141e6:	data_out=16'h2;
17'h141e7:	data_out=16'ha;
17'h141e8:	data_out=16'h9;
17'h141e9:	data_out=16'h17;
17'h141ea:	data_out=16'h9;
17'h141eb:	data_out=16'h8001;
17'h141ec:	data_out=16'h25;
17'h141ed:	data_out=16'h12;
17'h141ee:	data_out=16'h1;
17'h141ef:	data_out=16'hd;
17'h141f0:	data_out=16'h1;
17'h141f1:	data_out=16'h18;
17'h141f2:	data_out=16'h1a;
17'h141f3:	data_out=16'h16;
17'h141f4:	data_out=16'ha;
17'h141f5:	data_out=16'hd;
17'h141f6:	data_out=16'h7;
17'h141f7:	data_out=16'h16;
17'h141f8:	data_out=16'h8004;
17'h141f9:	data_out=16'h1f;
17'h141fa:	data_out=16'h10;
17'h141fb:	data_out=16'hc;
17'h141fc:	data_out=16'h9;
17'h141fd:	data_out=16'h7;
17'h141fe:	data_out=16'ha;
17'h141ff:	data_out=16'h14;
17'h14200:	data_out=16'h8;
17'h14201:	data_out=16'h8001;
17'h14202:	data_out=16'h8002;
17'h14203:	data_out=16'h8002;
17'h14204:	data_out=16'h9;
17'h14205:	data_out=16'h8001;
17'h14206:	data_out=16'h8001;
17'h14207:	data_out=16'h5;
17'h14208:	data_out=16'h4;
17'h14209:	data_out=16'h8005;
17'h1420a:	data_out=16'h5;
17'h1420b:	data_out=16'h8004;
17'h1420c:	data_out=16'h4;
17'h1420d:	data_out=16'h8007;
17'h1420e:	data_out=16'h4;
17'h1420f:	data_out=16'h8009;
17'h14210:	data_out=16'h2;
17'h14211:	data_out=16'h2;
17'h14212:	data_out=16'h9;
17'h14213:	data_out=16'h6;
17'h14214:	data_out=16'h8001;
17'h14215:	data_out=16'h8007;
17'h14216:	data_out=16'h2;
17'h14217:	data_out=16'h0;
17'h14218:	data_out=16'h7;
17'h14219:	data_out=16'h5;
17'h1421a:	data_out=16'h8002;
17'h1421b:	data_out=16'h3;
17'h1421c:	data_out=16'h8001;
17'h1421d:	data_out=16'h0;
17'h1421e:	data_out=16'h7;
17'h1421f:	data_out=16'h8003;
17'h14220:	data_out=16'h9;
17'h14221:	data_out=16'h8004;
17'h14222:	data_out=16'h4;
17'h14223:	data_out=16'h9;
17'h14224:	data_out=16'h4;
17'h14225:	data_out=16'h8006;
17'h14226:	data_out=16'h4;
17'h14227:	data_out=16'h8002;
17'h14228:	data_out=16'h8002;
17'h14229:	data_out=16'h0;
17'h1422a:	data_out=16'h4;
17'h1422b:	data_out=16'h8007;
17'h1422c:	data_out=16'h2;
17'h1422d:	data_out=16'h8002;
17'h1422e:	data_out=16'h8007;
17'h1422f:	data_out=16'h8005;
17'h14230:	data_out=16'h9;
17'h14231:	data_out=16'h8007;
17'h14232:	data_out=16'h8008;
17'h14233:	data_out=16'h8001;
17'h14234:	data_out=16'h8005;
17'h14235:	data_out=16'h4;
17'h14236:	data_out=16'h8;
17'h14237:	data_out=16'h8007;
17'h14238:	data_out=16'h8000;
17'h14239:	data_out=16'h8003;
17'h1423a:	data_out=16'h5;
17'h1423b:	data_out=16'h8;
17'h1423c:	data_out=16'h7;
17'h1423d:	data_out=16'h4;
17'h1423e:	data_out=16'h8004;
17'h1423f:	data_out=16'h7;
17'h14240:	data_out=16'h8;
17'h14241:	data_out=16'h9;
17'h14242:	data_out=16'h6;
17'h14243:	data_out=16'h3;
17'h14244:	data_out=16'h8006;
17'h14245:	data_out=16'h2;
17'h14246:	data_out=16'h8008;
17'h14247:	data_out=16'h1;
17'h14248:	data_out=16'h8007;
17'h14249:	data_out=16'h5;
17'h1424a:	data_out=16'h3;
17'h1424b:	data_out=16'h4;
17'h1424c:	data_out=16'h8006;
17'h1424d:	data_out=16'h5;
17'h1424e:	data_out=16'h8;
17'h1424f:	data_out=16'h8007;
17'h14250:	data_out=16'h7;
17'h14251:	data_out=16'h8009;
17'h14252:	data_out=16'h1;
17'h14253:	data_out=16'h8007;
17'h14254:	data_out=16'h4;
17'h14255:	data_out=16'h0;
17'h14256:	data_out=16'h8004;
17'h14257:	data_out=16'h8005;
17'h14258:	data_out=16'h7;
17'h14259:	data_out=16'h8008;
17'h1425a:	data_out=16'h8007;
17'h1425b:	data_out=16'h5;
17'h1425c:	data_out=16'h5;
17'h1425d:	data_out=16'h8002;
17'h1425e:	data_out=16'h3;
17'h1425f:	data_out=16'h4;
17'h14260:	data_out=16'h8002;
17'h14261:	data_out=16'h0;
17'h14262:	data_out=16'h8002;
17'h14263:	data_out=16'h1;
17'h14264:	data_out=16'h8007;
17'h14265:	data_out=16'h8001;
17'h14266:	data_out=16'h8007;
17'h14267:	data_out=16'h8006;
17'h14268:	data_out=16'h8006;
17'h14269:	data_out=16'h5;
17'h1426a:	data_out=16'h7;
17'h1426b:	data_out=16'h8003;
17'h1426c:	data_out=16'h1;
17'h1426d:	data_out=16'h7;
17'h1426e:	data_out=16'h8001;
17'h1426f:	data_out=16'h8001;
17'h14270:	data_out=16'h7;
17'h14271:	data_out=16'h8008;
17'h14272:	data_out=16'h2;
17'h14273:	data_out=16'h2;
17'h14274:	data_out=16'h1;
17'h14275:	data_out=16'h6;
17'h14276:	data_out=16'h6;
17'h14277:	data_out=16'h8001;
17'h14278:	data_out=16'h7;
17'h14279:	data_out=16'h8;
17'h1427a:	data_out=16'h8005;
17'h1427b:	data_out=16'h3;
17'h1427c:	data_out=16'h8003;
17'h1427d:	data_out=16'h7;
17'h1427e:	data_out=16'h8002;
17'h1427f:	data_out=16'h3;
17'h14280:	data_out=16'h8002;
17'h14281:	data_out=16'h4;
17'h14282:	data_out=16'h8005;
17'h14283:	data_out=16'h8000;
17'h14284:	data_out=16'h8006;
17'h14285:	data_out=16'h8003;
17'h14286:	data_out=16'h3;
17'h14287:	data_out=16'h8003;
17'h14288:	data_out=16'h8007;
17'h14289:	data_out=16'h1;
17'h1428a:	data_out=16'h3;
17'h1428b:	data_out=16'h3;
17'h1428c:	data_out=16'h8001;
17'h1428d:	data_out=16'h8007;
17'h1428e:	data_out=16'h8007;
17'h1428f:	data_out=16'h8003;
17'h14290:	data_out=16'h8006;
17'h14291:	data_out=16'h4;
17'h14292:	data_out=16'h8;
17'h14293:	data_out=16'h4;
17'h14294:	data_out=16'h1;
17'h14295:	data_out=16'h5;
17'h14296:	data_out=16'h8006;
17'h14297:	data_out=16'h8000;
17'h14298:	data_out=16'h4;
17'h14299:	data_out=16'h8002;
17'h1429a:	data_out=16'h8007;
17'h1429b:	data_out=16'h8009;
17'h1429c:	data_out=16'h8004;
17'h1429d:	data_out=16'h0;
17'h1429e:	data_out=16'h4;
17'h1429f:	data_out=16'h3;
17'h142a0:	data_out=16'h8005;
17'h142a1:	data_out=16'h8;
17'h142a2:	data_out=16'h8006;
17'h142a3:	data_out=16'h8002;
17'h142a4:	data_out=16'h8004;
17'h142a5:	data_out=16'h6;
17'h142a6:	data_out=16'h4;
17'h142a7:	data_out=16'h8002;
17'h142a8:	data_out=16'h8002;
17'h142a9:	data_out=16'h8002;
17'h142aa:	data_out=16'h8008;
17'h142ab:	data_out=16'h6;
17'h142ac:	data_out=16'h8000;
17'h142ad:	data_out=16'h8006;
17'h142ae:	data_out=16'h8006;
17'h142af:	data_out=16'h3;
17'h142b0:	data_out=16'h7;
17'h142b1:	data_out=16'h8007;
17'h142b2:	data_out=16'h8002;
17'h142b3:	data_out=16'h8001;
17'h142b4:	data_out=16'h7;
17'h142b5:	data_out=16'h1;
17'h142b6:	data_out=16'h8;
17'h142b7:	data_out=16'h1;
17'h142b8:	data_out=16'h9;
17'h142b9:	data_out=16'h8008;
17'h142ba:	data_out=16'h1;
17'h142bb:	data_out=16'h8004;
17'h142bc:	data_out=16'h2;
17'h142bd:	data_out=16'h8005;
17'h142be:	data_out=16'h8;
17'h142bf:	data_out=16'h6;
17'h142c0:	data_out=16'h8006;
17'h142c1:	data_out=16'h8007;
17'h142c2:	data_out=16'h8005;
17'h142c3:	data_out=16'h8001;
17'h142c4:	data_out=16'h8;
17'h142c5:	data_out=16'h8;
17'h142c6:	data_out=16'h6;
17'h142c7:	data_out=16'h8003;
17'h142c8:	data_out=16'h8003;
17'h142c9:	data_out=16'h6;
17'h142ca:	data_out=16'h8006;
17'h142cb:	data_out=16'h6;
17'h142cc:	data_out=16'h8009;
17'h142cd:	data_out=16'h8003;
17'h142ce:	data_out=16'h8001;
17'h142cf:	data_out=16'h7;
17'h142d0:	data_out=16'h8002;
17'h142d1:	data_out=16'h6;
17'h142d2:	data_out=16'h8002;
17'h142d3:	data_out=16'h8004;
17'h142d4:	data_out=16'h8002;
17'h142d5:	data_out=16'h8003;
17'h142d6:	data_out=16'h6;
17'h142d7:	data_out=16'h8002;
17'h142d8:	data_out=16'h8002;
17'h142d9:	data_out=16'h8002;
17'h142da:	data_out=16'h2;
17'h142db:	data_out=16'h9;
17'h142dc:	data_out=16'h2;
17'h142dd:	data_out=16'h1;
17'h142de:	data_out=16'h6;
17'h142df:	data_out=16'h6;
17'h142e0:	data_out=16'h3;
17'h142e1:	data_out=16'h8009;
17'h142e2:	data_out=16'h8005;
17'h142e3:	data_out=16'h2;
17'h142e4:	data_out=16'h8;
17'h142e5:	data_out=16'h8008;
17'h142e6:	data_out=16'h8;
17'h142e7:	data_out=16'h8004;
17'h142e8:	data_out=16'h7;
17'h142e9:	data_out=16'h8007;
17'h142ea:	data_out=16'h8008;
17'h142eb:	data_out=16'h8;
17'h142ec:	data_out=16'h8002;
17'h142ed:	data_out=16'h0;
17'h142ee:	data_out=16'h6;
17'h142ef:	data_out=16'h6;
17'h142f0:	data_out=16'h8003;
17'h142f1:	data_out=16'h8006;
17'h142f2:	data_out=16'h8007;
17'h142f3:	data_out=16'h4;
17'h142f4:	data_out=16'h0;
17'h142f5:	data_out=16'h8;
17'h142f6:	data_out=16'h8007;
17'h142f7:	data_out=16'h8;
17'h142f8:	data_out=16'h8004;
17'h142f9:	data_out=16'h4;
17'h142fa:	data_out=16'h8;
17'h142fb:	data_out=16'h8;
17'h142fc:	data_out=16'h8003;
17'h142fd:	data_out=16'h4;
17'h142fe:	data_out=16'h4;
17'h142ff:	data_out=16'h9;
17'h14300:	data_out=16'h810b;
17'h14301:	data_out=16'h141;
17'h14302:	data_out=16'h152;
17'h14303:	data_out=16'h13d;
17'h14304:	data_out=16'h222;
17'h14305:	data_out=16'h3ee;
17'h14306:	data_out=16'h2c5;
17'h14307:	data_out=16'h26d;
17'h14308:	data_out=16'h21d;
17'h14309:	data_out=16'h84;
17'h1430a:	data_out=16'hf1;
17'h1430b:	data_out=16'h1fd;
17'h1430c:	data_out=16'h349;
17'h1430d:	data_out=16'h51;
17'h1430e:	data_out=16'ha7;
17'h1430f:	data_out=16'h236;
17'h14310:	data_out=16'h8032;
17'h14311:	data_out=16'h2e8;
17'h14312:	data_out=16'h11e;
17'h14313:	data_out=16'he9;
17'h14314:	data_out=16'hf2;
17'h14315:	data_out=16'h7;
17'h14316:	data_out=16'hb9;
17'h14317:	data_out=16'hcf;
17'h14318:	data_out=16'h9f;
17'h14319:	data_out=16'h127;
17'h1431a:	data_out=16'h23f;
17'h1431b:	data_out=16'h15b;
17'h1431c:	data_out=16'h34b;
17'h1431d:	data_out=16'h1ad;
17'h1431e:	data_out=16'h1c5;
17'h1431f:	data_out=16'h2c3;
17'h14320:	data_out=16'h1ac;
17'h14321:	data_out=16'ha3;
17'h14322:	data_out=16'h8022;
17'h14323:	data_out=16'h804b;
17'h14324:	data_out=16'h805c;
17'h14325:	data_out=16'hfd;
17'h14326:	data_out=16'h1d2;
17'h14327:	data_out=16'h216;
17'h14328:	data_out=16'hb9;
17'h14329:	data_out=16'h8070;
17'h1432a:	data_out=16'hf7;
17'h1432b:	data_out=16'hf6;
17'h1432c:	data_out=16'h199;
17'h1432d:	data_out=16'h8198;
17'h1432e:	data_out=16'hee;
17'h1432f:	data_out=16'h16b;
17'h14330:	data_out=16'h32f;
17'h14331:	data_out=16'h247;
17'h14332:	data_out=16'h31e;
17'h14333:	data_out=16'h143;
17'h14334:	data_out=16'h15b;
17'h14335:	data_out=16'h4e9;
17'h14336:	data_out=16'h1a8;
17'h14337:	data_out=16'h18c;
17'h14338:	data_out=16'h26c;
17'h14339:	data_out=16'h18a;
17'h1433a:	data_out=16'h811a;
17'h1433b:	data_out=16'h32b;
17'h1433c:	data_out=16'h1a6;
17'h1433d:	data_out=16'h173;
17'h1433e:	data_out=16'hc8;
17'h1433f:	data_out=16'h3ed;
17'h14340:	data_out=16'hda;
17'h14341:	data_out=16'h28f;
17'h14342:	data_out=16'ha;
17'h14343:	data_out=16'h26c;
17'h14344:	data_out=16'h23f;
17'h14345:	data_out=16'h802c;
17'h14346:	data_out=16'hde;
17'h14347:	data_out=16'h5c;
17'h14348:	data_out=16'h85;
17'h14349:	data_out=16'hfd;
17'h1434a:	data_out=16'h24c;
17'h1434b:	data_out=16'h14e;
17'h1434c:	data_out=16'h9f;
17'h1434d:	data_out=16'h803e;
17'h1434e:	data_out=16'h178;
17'h1434f:	data_out=16'hde;
17'h14350:	data_out=16'h56;
17'h14351:	data_out=16'h2c6;
17'h14352:	data_out=16'h8005;
17'h14353:	data_out=16'h225;
17'h14354:	data_out=16'h13c;
17'h14355:	data_out=16'h346;
17'h14356:	data_out=16'h17e;
17'h14357:	data_out=16'ha3;
17'h14358:	data_out=16'h1de;
17'h14359:	data_out=16'h143;
17'h1435a:	data_out=16'h5c;
17'h1435b:	data_out=16'h416;
17'h1435c:	data_out=16'h25b;
17'h1435d:	data_out=16'h8a;
17'h1435e:	data_out=16'h166;
17'h1435f:	data_out=16'h43;
17'h14360:	data_out=16'h140;
17'h14361:	data_out=16'h3cd;
17'h14362:	data_out=16'h1f4;
17'h14363:	data_out=16'h109;
17'h14364:	data_out=16'h198;
17'h14365:	data_out=16'h1bc;
17'h14366:	data_out=16'h13d;
17'h14367:	data_out=16'h6e;
17'h14368:	data_out=16'hac;
17'h14369:	data_out=16'h21b;
17'h1436a:	data_out=16'h9f;
17'h1436b:	data_out=16'h309;
17'h1436c:	data_out=16'h81b7;
17'h1436d:	data_out=16'h158;
17'h1436e:	data_out=16'h96;
17'h1436f:	data_out=16'h22a;
17'h14370:	data_out=16'h9d;
17'h14371:	data_out=16'h1df;
17'h14372:	data_out=16'h1df;
17'h14373:	data_out=16'h2b3;
17'h14374:	data_out=16'h332;
17'h14375:	data_out=16'h3c6;
17'h14376:	data_out=16'h155;
17'h14377:	data_out=16'h114;
17'h14378:	data_out=16'h267;
17'h14379:	data_out=16'h21e;
17'h1437a:	data_out=16'h110;
17'h1437b:	data_out=16'hc2;
17'h1437c:	data_out=16'hed;
17'h1437d:	data_out=16'h367;
17'h1437e:	data_out=16'h125;
17'h1437f:	data_out=16'h13d;
17'h14380:	data_out=16'h89fe;
17'h14381:	data_out=16'h26b;
17'h14382:	data_out=16'h4a5;
17'h14383:	data_out=16'h810d;
17'h14384:	data_out=16'h3f8;
17'h14385:	data_out=16'ha00;
17'h14386:	data_out=16'h80d;
17'h14387:	data_out=16'h80ef;
17'h14388:	data_out=16'h244;
17'h14389:	data_out=16'h8772;
17'h1438a:	data_out=16'h8541;
17'h1438b:	data_out=16'h8f2;
17'h1438c:	data_out=16'h9ab;
17'h1438d:	data_out=16'hd6;
17'h1438e:	data_out=16'h19f;
17'h1438f:	data_out=16'h473;
17'h14390:	data_out=16'h81e1;
17'h14391:	data_out=16'ha00;
17'h14392:	data_out=16'h165;
17'h14393:	data_out=16'h818a;
17'h14394:	data_out=16'h642;
17'h14395:	data_out=16'h81ca;
17'h14396:	data_out=16'h8249;
17'h14397:	data_out=16'h512;
17'h14398:	data_out=16'h89;
17'h14399:	data_out=16'ha00;
17'h1439a:	data_out=16'h4b7;
17'h1439b:	data_out=16'h9ff;
17'h1439c:	data_out=16'h9fd;
17'h1439d:	data_out=16'h674;
17'h1439e:	data_out=16'h5fc;
17'h1439f:	data_out=16'h603;
17'h143a0:	data_out=16'ha00;
17'h143a1:	data_out=16'h1b9;
17'h143a2:	data_out=16'h8779;
17'h143a3:	data_out=16'h83f8;
17'h143a4:	data_out=16'h83f6;
17'h143a5:	data_out=16'h82f9;
17'h143a6:	data_out=16'h8685;
17'h143a7:	data_out=16'ha00;
17'h143a8:	data_out=16'h1fd;
17'h143a9:	data_out=16'h857b;
17'h143aa:	data_out=16'h85a0;
17'h143ab:	data_out=16'ha00;
17'h143ac:	data_out=16'h825e;
17'h143ad:	data_out=16'h8a00;
17'h143ae:	data_out=16'h25b;
17'h143af:	data_out=16'h8e0;
17'h143b0:	data_out=16'h26a;
17'h143b1:	data_out=16'h64f;
17'h143b2:	data_out=16'h1bd;
17'h143b3:	data_out=16'h769;
17'h143b4:	data_out=16'h86;
17'h143b5:	data_out=16'h9fe;
17'h143b6:	data_out=16'h464;
17'h143b7:	data_out=16'h48e;
17'h143b8:	data_out=16'h6a0;
17'h143b9:	data_out=16'h7ec;
17'h143ba:	data_out=16'h8a00;
17'h143bb:	data_out=16'h794;
17'h143bc:	data_out=16'h5d5;
17'h143bd:	data_out=16'h804d;
17'h143be:	data_out=16'h200;
17'h143bf:	data_out=16'ha00;
17'h143c0:	data_out=16'h8201;
17'h143c1:	data_out=16'ha00;
17'h143c2:	data_out=16'h8a00;
17'h143c3:	data_out=16'h869;
17'h143c4:	data_out=16'h80c;
17'h143c5:	data_out=16'h81d5;
17'h143c6:	data_out=16'h8030;
17'h143c7:	data_out=16'h88ea;
17'h143c8:	data_out=16'h347;
17'h143c9:	data_out=16'h828a;
17'h143ca:	data_out=16'h375;
17'h143cb:	data_out=16'h9a;
17'h143cc:	data_out=16'h87a6;
17'h143cd:	data_out=16'h8737;
17'h143ce:	data_out=16'h295;
17'h143cf:	data_out=16'h8707;
17'h143d0:	data_out=16'h81a8;
17'h143d1:	data_out=16'h9fe;
17'h143d2:	data_out=16'h8748;
17'h143d3:	data_out=16'ha00;
17'h143d4:	data_out=16'h882;
17'h143d5:	data_out=16'h9f7;
17'h143d6:	data_out=16'h8496;
17'h143d7:	data_out=16'h856a;
17'h143d8:	data_out=16'h90a;
17'h143d9:	data_out=16'h82e5;
17'h143da:	data_out=16'h9fe;
17'h143db:	data_out=16'ha00;
17'h143dc:	data_out=16'ha00;
17'h143dd:	data_out=16'h8397;
17'h143de:	data_out=16'h784;
17'h143df:	data_out=16'h812c;
17'h143e0:	data_out=16'h8a00;
17'h143e1:	data_out=16'ha00;
17'h143e2:	data_out=16'h74b;
17'h143e3:	data_out=16'h856;
17'h143e4:	data_out=16'h498;
17'h143e5:	data_out=16'h5be;
17'h143e6:	data_out=16'ha00;
17'h143e7:	data_out=16'h8174;
17'h143e8:	data_out=16'h1cf;
17'h143e9:	data_out=16'hf6;
17'h143ea:	data_out=16'h170;
17'h143eb:	data_out=16'h7e3;
17'h143ec:	data_out=16'h89fe;
17'h143ed:	data_out=16'h802;
17'h143ee:	data_out=16'h180;
17'h143ef:	data_out=16'h23c;
17'h143f0:	data_out=16'h198;
17'h143f1:	data_out=16'h52c;
17'h143f2:	data_out=16'h8242;
17'h143f3:	data_out=16'h3dd;
17'h143f4:	data_out=16'h249;
17'h143f5:	data_out=16'ha00;
17'h143f6:	data_out=16'h9ff;
17'h143f7:	data_out=16'h82f8;
17'h143f8:	data_out=16'h7e1;
17'h143f9:	data_out=16'h36a;
17'h143fa:	data_out=16'h76b;
17'h143fb:	data_out=16'h201;
17'h143fc:	data_out=16'h176;
17'h143fd:	data_out=16'ha00;
17'h143fe:	data_out=16'h8300;
17'h143ff:	data_out=16'h83b4;
17'h14400:	data_out=16'h8857;
17'h14401:	data_out=16'ha00;
17'h14402:	data_out=16'h78a;
17'h14403:	data_out=16'h181;
17'h14404:	data_out=16'h81a3;
17'h14405:	data_out=16'h9fa;
17'h14406:	data_out=16'h3f4;
17'h14407:	data_out=16'h8a00;
17'h14408:	data_out=16'h7d8;
17'h14409:	data_out=16'h8a00;
17'h1440a:	data_out=16'h8a00;
17'h1440b:	data_out=16'h747;
17'h1440c:	data_out=16'h333;
17'h1440d:	data_out=16'h78a;
17'h1440e:	data_out=16'h8229;
17'h1440f:	data_out=16'h283;
17'h14410:	data_out=16'h8260;
17'h14411:	data_out=16'h9fc;
17'h14412:	data_out=16'h8562;
17'h14413:	data_out=16'h83ff;
17'h14414:	data_out=16'h9b9;
17'h14415:	data_out=16'h81a0;
17'h14416:	data_out=16'h8807;
17'h14417:	data_out=16'h8fc;
17'h14418:	data_out=16'hd1;
17'h14419:	data_out=16'h9fb;
17'h1441a:	data_out=16'h92;
17'h1441b:	data_out=16'h9f2;
17'h1441c:	data_out=16'h9f5;
17'h1441d:	data_out=16'h9fa;
17'h1441e:	data_out=16'h9bc;
17'h1441f:	data_out=16'hd2;
17'h14420:	data_out=16'ha00;
17'h14421:	data_out=16'h81e0;
17'h14422:	data_out=16'h8a00;
17'h14423:	data_out=16'h89fe;
17'h14424:	data_out=16'h89ff;
17'h14425:	data_out=16'h8a00;
17'h14426:	data_out=16'h8a00;
17'h14427:	data_out=16'ha00;
17'h14428:	data_out=16'h8146;
17'h14429:	data_out=16'hb;
17'h1442a:	data_out=16'h89f9;
17'h1442b:	data_out=16'ha00;
17'h1442c:	data_out=16'h875d;
17'h1442d:	data_out=16'h8a00;
17'h1442e:	data_out=16'h481;
17'h1442f:	data_out=16'ha00;
17'h14430:	data_out=16'h8a00;
17'h14431:	data_out=16'h9ff;
17'h14432:	data_out=16'h8a00;
17'h14433:	data_out=16'h9f6;
17'h14434:	data_out=16'h8952;
17'h14435:	data_out=16'h9b2;
17'h14436:	data_out=16'ha00;
17'h14437:	data_out=16'h64b;
17'h14438:	data_out=16'h9f7;
17'h14439:	data_out=16'h9fb;
17'h1443a:	data_out=16'h8a00;
17'h1443b:	data_out=16'hdd;
17'h1443c:	data_out=16'h937;
17'h1443d:	data_out=16'h256;
17'h1443e:	data_out=16'h8122;
17'h1443f:	data_out=16'h9fa;
17'h14440:	data_out=16'h8a00;
17'h14441:	data_out=16'ha00;
17'h14442:	data_out=16'h8a00;
17'h14443:	data_out=16'h833;
17'h14444:	data_out=16'h9ff;
17'h14445:	data_out=16'h827f;
17'h14446:	data_out=16'h83b2;
17'h14447:	data_out=16'h8a00;
17'h14448:	data_out=16'h772;
17'h14449:	data_out=16'h8a00;
17'h1444a:	data_out=16'h4ea;
17'h1444b:	data_out=16'h8a00;
17'h1444c:	data_out=16'h8a00;
17'h1444d:	data_out=16'h89ff;
17'h1444e:	data_out=16'h8016;
17'h1444f:	data_out=16'h8a00;
17'h14450:	data_out=16'h878d;
17'h14451:	data_out=16'h7b7;
17'h14452:	data_out=16'h8a00;
17'h14453:	data_out=16'ha00;
17'h14454:	data_out=16'ha00;
17'h14455:	data_out=16'h44f;
17'h14456:	data_out=16'h89f0;
17'h14457:	data_out=16'h89f8;
17'h14458:	data_out=16'h9ff;
17'h14459:	data_out=16'h8a00;
17'h1445a:	data_out=16'h9fa;
17'h1445b:	data_out=16'h9ff;
17'h1445c:	data_out=16'h9fb;
17'h1445d:	data_out=16'h810a;
17'h1445e:	data_out=16'h9fe;
17'h1445f:	data_out=16'h321;
17'h14460:	data_out=16'h8a00;
17'h14461:	data_out=16'h972;
17'h14462:	data_out=16'h6cc;
17'h14463:	data_out=16'h9f5;
17'h14464:	data_out=16'h1bd;
17'h14465:	data_out=16'h82b7;
17'h14466:	data_out=16'h9f5;
17'h14467:	data_out=16'h878b;
17'h14468:	data_out=16'h81ae;
17'h14469:	data_out=16'hfa;
17'h1446a:	data_out=16'h825e;
17'h1446b:	data_out=16'h9e9;
17'h1446c:	data_out=16'h89e8;
17'h1446d:	data_out=16'h9f6;
17'h1446e:	data_out=16'h825e;
17'h1446f:	data_out=16'h8766;
17'h14470:	data_out=16'h8240;
17'h14471:	data_out=16'h33c;
17'h14472:	data_out=16'h8a00;
17'h14473:	data_out=16'h820b;
17'h14474:	data_out=16'h8a00;
17'h14475:	data_out=16'h9fd;
17'h14476:	data_out=16'h9f3;
17'h14477:	data_out=16'h8a00;
17'h14478:	data_out=16'h56e;
17'h14479:	data_out=16'h4ed;
17'h1447a:	data_out=16'h9f2;
17'h1447b:	data_out=16'h80ea;
17'h1447c:	data_out=16'h699;
17'h1447d:	data_out=16'h9f9;
17'h1447e:	data_out=16'h8a00;
17'h1447f:	data_out=16'h86ef;
17'h14480:	data_out=16'h977;
17'h14481:	data_out=16'ha00;
17'h14482:	data_out=16'h89ed;
17'h14483:	data_out=16'h52b;
17'h14484:	data_out=16'h899a;
17'h14485:	data_out=16'h9eb;
17'h14486:	data_out=16'h8a00;
17'h14487:	data_out=16'h8a00;
17'h14488:	data_out=16'hff;
17'h14489:	data_out=16'h8a00;
17'h1448a:	data_out=16'h89fe;
17'h1448b:	data_out=16'h6b2;
17'h1448c:	data_out=16'h89fe;
17'h1448d:	data_out=16'h600;
17'h1448e:	data_out=16'h89ff;
17'h1448f:	data_out=16'h89ee;
17'h14490:	data_out=16'h89fd;
17'h14491:	data_out=16'h8715;
17'h14492:	data_out=16'h841e;
17'h14493:	data_out=16'h587;
17'h14494:	data_out=16'h9d7;
17'h14495:	data_out=16'h840d;
17'h14496:	data_out=16'h843b;
17'h14497:	data_out=16'h9a0;
17'h14498:	data_out=16'h887c;
17'h14499:	data_out=16'h6c9;
17'h1449a:	data_out=16'h849e;
17'h1449b:	data_out=16'h8cd;
17'h1449c:	data_out=16'ha00;
17'h1449d:	data_out=16'h659;
17'h1449e:	data_out=16'h944;
17'h1449f:	data_out=16'h855a;
17'h144a0:	data_out=16'ha00;
17'h144a1:	data_out=16'h89fb;
17'h144a2:	data_out=16'h8a00;
17'h144a3:	data_out=16'h89f4;
17'h144a4:	data_out=16'h89f4;
17'h144a5:	data_out=16'h8a00;
17'h144a6:	data_out=16'h8a00;
17'h144a7:	data_out=16'h9fe;
17'h144a8:	data_out=16'h8960;
17'h144a9:	data_out=16'h6c9;
17'h144aa:	data_out=16'h89e7;
17'h144ab:	data_out=16'ha00;
17'h144ac:	data_out=16'h830f;
17'h144ad:	data_out=16'h8a00;
17'h144ae:	data_out=16'h889c;
17'h144af:	data_out=16'ha00;
17'h144b0:	data_out=16'h8a00;
17'h144b1:	data_out=16'h9ff;
17'h144b2:	data_out=16'h8a00;
17'h144b3:	data_out=16'h9f9;
17'h144b4:	data_out=16'h8374;
17'h144b5:	data_out=16'h6f2;
17'h144b6:	data_out=16'h9ff;
17'h144b7:	data_out=16'h89fa;
17'h144b8:	data_out=16'h9f6;
17'h144b9:	data_out=16'ha00;
17'h144ba:	data_out=16'h8a00;
17'h144bb:	data_out=16'h884a;
17'h144bc:	data_out=16'h9cd;
17'h144bd:	data_out=16'h82d3;
17'h144be:	data_out=16'h895b;
17'h144bf:	data_out=16'h9ec;
17'h144c0:	data_out=16'h8a00;
17'h144c1:	data_out=16'h9fe;
17'h144c2:	data_out=16'h8a00;
17'h144c3:	data_out=16'h848a;
17'h144c4:	data_out=16'ha00;
17'h144c5:	data_out=16'h849a;
17'h144c6:	data_out=16'h89f7;
17'h144c7:	data_out=16'h89fa;
17'h144c8:	data_out=16'h862c;
17'h144c9:	data_out=16'h8a00;
17'h144ca:	data_out=16'h4e8;
17'h144cb:	data_out=16'h8a00;
17'h144cc:	data_out=16'h8a00;
17'h144cd:	data_out=16'h8a00;
17'h144ce:	data_out=16'h8860;
17'h144cf:	data_out=16'h8a00;
17'h144d0:	data_out=16'h8595;
17'h144d1:	data_out=16'h4e3;
17'h144d2:	data_out=16'h8a00;
17'h144d3:	data_out=16'h9ff;
17'h144d4:	data_out=16'ha00;
17'h144d5:	data_out=16'h812b;
17'h144d6:	data_out=16'h89e3;
17'h144d7:	data_out=16'h89f8;
17'h144d8:	data_out=16'ha00;
17'h144d9:	data_out=16'h8a00;
17'h144da:	data_out=16'h9bb;
17'h144db:	data_out=16'h9fe;
17'h144dc:	data_out=16'h9f0;
17'h144dd:	data_out=16'h8839;
17'h144de:	data_out=16'ha00;
17'h144df:	data_out=16'h8183;
17'h144e0:	data_out=16'h8a00;
17'h144e1:	data_out=16'h676;
17'h144e2:	data_out=16'h5e6;
17'h144e3:	data_out=16'h9f7;
17'h144e4:	data_out=16'h8903;
17'h144e5:	data_out=16'h8a00;
17'h144e6:	data_out=16'h62;
17'h144e7:	data_out=16'h8a00;
17'h144e8:	data_out=16'h89c9;
17'h144e9:	data_out=16'h882f;
17'h144ea:	data_out=16'h89ff;
17'h144eb:	data_out=16'h75a;
17'h144ec:	data_out=16'h8528;
17'h144ed:	data_out=16'h9f8;
17'h144ee:	data_out=16'h89ff;
17'h144ef:	data_out=16'h8a00;
17'h144f0:	data_out=16'h89ff;
17'h144f1:	data_out=16'h809f;
17'h144f2:	data_out=16'h8a00;
17'h144f3:	data_out=16'h8a00;
17'h144f4:	data_out=16'h8a00;
17'h144f5:	data_out=16'h981;
17'h144f6:	data_out=16'h723;
17'h144f7:	data_out=16'h8a00;
17'h144f8:	data_out=16'h85be;
17'h144f9:	data_out=16'h897d;
17'h144fa:	data_out=16'h9f3;
17'h144fb:	data_out=16'h895a;
17'h144fc:	data_out=16'ha2;
17'h144fd:	data_out=16'h82b7;
17'h144fe:	data_out=16'h8a00;
17'h144ff:	data_out=16'h8630;
17'h14500:	data_out=16'ha00;
17'h14501:	data_out=16'ha00;
17'h14502:	data_out=16'h89f6;
17'h14503:	data_out=16'h808a;
17'h14504:	data_out=16'h89dd;
17'h14505:	data_out=16'h7a3;
17'h14506:	data_out=16'h8a00;
17'h14507:	data_out=16'h8a00;
17'h14508:	data_out=16'h80bb;
17'h14509:	data_out=16'h8a00;
17'h1450a:	data_out=16'h8a00;
17'h1450b:	data_out=16'h861;
17'h1450c:	data_out=16'h89f6;
17'h1450d:	data_out=16'h88a9;
17'h1450e:	data_out=16'h8a00;
17'h1450f:	data_out=16'h89e7;
17'h14510:	data_out=16'h89fe;
17'h14511:	data_out=16'h8057;
17'h14512:	data_out=16'h8245;
17'h14513:	data_out=16'h1e2;
17'h14514:	data_out=16'h7e6;
17'h14515:	data_out=16'h89c8;
17'h14516:	data_out=16'h89dd;
17'h14517:	data_out=16'h8da;
17'h14518:	data_out=16'h89d5;
17'h14519:	data_out=16'h9c5;
17'h1451a:	data_out=16'h89e1;
17'h1451b:	data_out=16'h4ef;
17'h1451c:	data_out=16'h9f8;
17'h1451d:	data_out=16'h9fd;
17'h1451e:	data_out=16'h60a;
17'h1451f:	data_out=16'h89ff;
17'h14520:	data_out=16'ha00;
17'h14521:	data_out=16'h8a00;
17'h14522:	data_out=16'h8a00;
17'h14523:	data_out=16'h89f7;
17'h14524:	data_out=16'h89f9;
17'h14525:	data_out=16'h8a00;
17'h14526:	data_out=16'h89f2;
17'h14527:	data_out=16'h9fc;
17'h14528:	data_out=16'h8a00;
17'h14529:	data_out=16'h9b7;
17'h1452a:	data_out=16'h89d4;
17'h1452b:	data_out=16'ha00;
17'h1452c:	data_out=16'h89cc;
17'h1452d:	data_out=16'h1ad;
17'h1452e:	data_out=16'h8409;
17'h1452f:	data_out=16'ha00;
17'h14530:	data_out=16'h8a00;
17'h14531:	data_out=16'h9fd;
17'h14532:	data_out=16'h8a00;
17'h14533:	data_out=16'h9f3;
17'h14534:	data_out=16'h9f9;
17'h14535:	data_out=16'h8270;
17'h14536:	data_out=16'h9ff;
17'h14537:	data_out=16'h89fe;
17'h14538:	data_out=16'h9fd;
17'h14539:	data_out=16'h9fd;
17'h1453a:	data_out=16'h8a00;
17'h1453b:	data_out=16'h89fd;
17'h1453c:	data_out=16'h9fc;
17'h1453d:	data_out=16'h83d5;
17'h1453e:	data_out=16'h8a00;
17'h1453f:	data_out=16'h78d;
17'h14540:	data_out=16'h8a00;
17'h14541:	data_out=16'h2d4;
17'h14542:	data_out=16'h8a00;
17'h14543:	data_out=16'h8806;
17'h14544:	data_out=16'h9f7;
17'h14545:	data_out=16'h89c8;
17'h14546:	data_out=16'h973;
17'h14547:	data_out=16'h89ea;
17'h14548:	data_out=16'h8614;
17'h14549:	data_out=16'h8a00;
17'h1454a:	data_out=16'h83e;
17'h1454b:	data_out=16'h8a00;
17'h1454c:	data_out=16'h8a00;
17'h1454d:	data_out=16'h8a00;
17'h1454e:	data_out=16'h8422;
17'h1454f:	data_out=16'h8a00;
17'h14550:	data_out=16'h89f1;
17'h14551:	data_out=16'h89fd;
17'h14552:	data_out=16'h8a00;
17'h14553:	data_out=16'h9ff;
17'h14554:	data_out=16'ha00;
17'h14555:	data_out=16'h8a00;
17'h14556:	data_out=16'h89f1;
17'h14557:	data_out=16'h8a00;
17'h14558:	data_out=16'h89bb;
17'h14559:	data_out=16'h8a00;
17'h1455a:	data_out=16'h986;
17'h1455b:	data_out=16'h9f3;
17'h1455c:	data_out=16'h9e1;
17'h1455d:	data_out=16'h88ed;
17'h1455e:	data_out=16'ha00;
17'h1455f:	data_out=16'h85d3;
17'h14560:	data_out=16'h8a00;
17'h14561:	data_out=16'h18;
17'h14562:	data_out=16'h60b;
17'h14563:	data_out=16'h9f2;
17'h14564:	data_out=16'h87a7;
17'h14565:	data_out=16'h8a00;
17'h14566:	data_out=16'h869e;
17'h14567:	data_out=16'h87ef;
17'h14568:	data_out=16'h8a00;
17'h14569:	data_out=16'h892c;
17'h1456a:	data_out=16'h8a00;
17'h1456b:	data_out=16'h82e6;
17'h1456c:	data_out=16'ha00;
17'h1456d:	data_out=16'h9f4;
17'h1456e:	data_out=16'h8a00;
17'h1456f:	data_out=16'h89ff;
17'h14570:	data_out=16'h8a00;
17'h14571:	data_out=16'h805c;
17'h14572:	data_out=16'h89ff;
17'h14573:	data_out=16'h8a00;
17'h14574:	data_out=16'h8a00;
17'h14575:	data_out=16'h43b;
17'h14576:	data_out=16'h9e7;
17'h14577:	data_out=16'h8a00;
17'h14578:	data_out=16'h898a;
17'h14579:	data_out=16'h89c6;
17'h1457a:	data_out=16'h9ea;
17'h1457b:	data_out=16'h8a00;
17'h1457c:	data_out=16'h82fb;
17'h1457d:	data_out=16'h888b;
17'h1457e:	data_out=16'h871d;
17'h1457f:	data_out=16'h8987;
17'h14580:	data_out=16'ha00;
17'h14581:	data_out=16'ha00;
17'h14582:	data_out=16'h89e1;
17'h14583:	data_out=16'h8794;
17'h14584:	data_out=16'h89e9;
17'h14585:	data_out=16'h358;
17'h14586:	data_out=16'h8a00;
17'h14587:	data_out=16'h8a00;
17'h14588:	data_out=16'h371;
17'h14589:	data_out=16'h8a00;
17'h1458a:	data_out=16'h89f6;
17'h1458b:	data_out=16'h9ef;
17'h1458c:	data_out=16'h8a00;
17'h1458d:	data_out=16'h8a00;
17'h1458e:	data_out=16'h89f9;
17'h1458f:	data_out=16'h8a00;
17'h14590:	data_out=16'h8a00;
17'h14591:	data_out=16'ha00;
17'h14592:	data_out=16'h5e6;
17'h14593:	data_out=16'h84ea;
17'h14594:	data_out=16'h3c6;
17'h14595:	data_out=16'h89e0;
17'h14596:	data_out=16'h89ff;
17'h14597:	data_out=16'h36a;
17'h14598:	data_out=16'h89f4;
17'h14599:	data_out=16'h9ce;
17'h1459a:	data_out=16'h89fa;
17'h1459b:	data_out=16'h5c6;
17'h1459c:	data_out=16'h9e5;
17'h1459d:	data_out=16'h9f5;
17'h1459e:	data_out=16'h363;
17'h1459f:	data_out=16'h89ff;
17'h145a0:	data_out=16'h9e9;
17'h145a1:	data_out=16'h89fa;
17'h145a2:	data_out=16'h8a00;
17'h145a3:	data_out=16'h8006;
17'h145a4:	data_out=16'h8038;
17'h145a5:	data_out=16'h8a00;
17'h145a6:	data_out=16'h89bd;
17'h145a7:	data_out=16'h9e2;
17'h145a8:	data_out=16'h89fb;
17'h145a9:	data_out=16'h9fa;
17'h145aa:	data_out=16'h89c8;
17'h145ab:	data_out=16'h9f3;
17'h145ac:	data_out=16'h89ff;
17'h145ad:	data_out=16'h9e3;
17'h145ae:	data_out=16'h9b1;
17'h145af:	data_out=16'h9dd;
17'h145b0:	data_out=16'h8a00;
17'h145b1:	data_out=16'h9de;
17'h145b2:	data_out=16'h89ff;
17'h145b3:	data_out=16'h9c0;
17'h145b4:	data_out=16'ha00;
17'h145b5:	data_out=16'h87cb;
17'h145b6:	data_out=16'h9f8;
17'h145b7:	data_out=16'h89e2;
17'h145b8:	data_out=16'h9f4;
17'h145b9:	data_out=16'h9d0;
17'h145ba:	data_out=16'h8a00;
17'h145bb:	data_out=16'h89f0;
17'h145bc:	data_out=16'ha00;
17'h145bd:	data_out=16'h851b;
17'h145be:	data_out=16'h89fb;
17'h145bf:	data_out=16'h33d;
17'h145c0:	data_out=16'h89ff;
17'h145c1:	data_out=16'h8023;
17'h145c2:	data_out=16'h89fd;
17'h145c3:	data_out=16'h861a;
17'h145c4:	data_out=16'h441;
17'h145c5:	data_out=16'h89e2;
17'h145c6:	data_out=16'h9ff;
17'h145c7:	data_out=16'h8a00;
17'h145c8:	data_out=16'h8a00;
17'h145c9:	data_out=16'h8a00;
17'h145ca:	data_out=16'h80e1;
17'h145cb:	data_out=16'h8934;
17'h145cc:	data_out=16'h8a00;
17'h145cd:	data_out=16'h8a00;
17'h145ce:	data_out=16'h871;
17'h145cf:	data_out=16'h8a00;
17'h145d0:	data_out=16'h89ff;
17'h145d1:	data_out=16'h8a00;
17'h145d2:	data_out=16'h8a00;
17'h145d3:	data_out=16'ha00;
17'h145d4:	data_out=16'h9ed;
17'h145d5:	data_out=16'h8a00;
17'h145d6:	data_out=16'h89be;
17'h145d7:	data_out=16'h89e3;
17'h145d8:	data_out=16'h897c;
17'h145d9:	data_out=16'h89fe;
17'h145da:	data_out=16'h963;
17'h145db:	data_out=16'h9de;
17'h145dc:	data_out=16'h9e1;
17'h145dd:	data_out=16'h8941;
17'h145de:	data_out=16'h9da;
17'h145df:	data_out=16'h865e;
17'h145e0:	data_out=16'h89e9;
17'h145e1:	data_out=16'h81cf;
17'h145e2:	data_out=16'h86f;
17'h145e3:	data_out=16'h9c0;
17'h145e4:	data_out=16'h809;
17'h145e5:	data_out=16'h89ff;
17'h145e6:	data_out=16'h8a00;
17'h145e7:	data_out=16'h811d;
17'h145e8:	data_out=16'h89fb;
17'h145e9:	data_out=16'h874b;
17'h145ea:	data_out=16'h89f8;
17'h145eb:	data_out=16'h89c5;
17'h145ec:	data_out=16'h9da;
17'h145ed:	data_out=16'h9c2;
17'h145ee:	data_out=16'h89f8;
17'h145ef:	data_out=16'h8a00;
17'h145f0:	data_out=16'h89f8;
17'h145f1:	data_out=16'h87d8;
17'h145f2:	data_out=16'h89fd;
17'h145f3:	data_out=16'h89fe;
17'h145f4:	data_out=16'h8a00;
17'h145f5:	data_out=16'h808c;
17'h145f6:	data_out=16'h9d0;
17'h145f7:	data_out=16'h8a00;
17'h145f8:	data_out=16'h89fe;
17'h145f9:	data_out=16'h88cf;
17'h145fa:	data_out=16'h81a;
17'h145fb:	data_out=16'h89fb;
17'h145fc:	data_out=16'h879b;
17'h145fd:	data_out=16'h89cd;
17'h145fe:	data_out=16'h1a;
17'h145ff:	data_out=16'h89fc;
17'h14600:	data_out=16'h9da;
17'h14601:	data_out=16'ha00;
17'h14602:	data_out=16'h987;
17'h14603:	data_out=16'h86b0;
17'h14604:	data_out=16'h89d4;
17'h14605:	data_out=16'hcc;
17'h14606:	data_out=16'h8a00;
17'h14607:	data_out=16'h8a00;
17'h14608:	data_out=16'h834e;
17'h14609:	data_out=16'h8a00;
17'h1460a:	data_out=16'h81a4;
17'h1460b:	data_out=16'h9e0;
17'h1460c:	data_out=16'h8a00;
17'h1460d:	data_out=16'h8a00;
17'h1460e:	data_out=16'h6dc;
17'h1460f:	data_out=16'h89fc;
17'h14610:	data_out=16'h8928;
17'h14611:	data_out=16'ha00;
17'h14612:	data_out=16'h8455;
17'h14613:	data_out=16'h88c;
17'h14614:	data_out=16'h3c;
17'h14615:	data_out=16'h89e6;
17'h14616:	data_out=16'h89fd;
17'h14617:	data_out=16'h8404;
17'h14618:	data_out=16'h89f8;
17'h14619:	data_out=16'h8458;
17'h1461a:	data_out=16'h89f8;
17'h1461b:	data_out=16'h97a;
17'h1461c:	data_out=16'h9eb;
17'h1461d:	data_out=16'h9fc;
17'h1461e:	data_out=16'h81f5;
17'h1461f:	data_out=16'h89e3;
17'h14620:	data_out=16'h9a7;
17'h14621:	data_out=16'h598;
17'h14622:	data_out=16'h88c7;
17'h14623:	data_out=16'ha00;
17'h14624:	data_out=16'ha00;
17'h14625:	data_out=16'h898b;
17'h14626:	data_out=16'ha00;
17'h14627:	data_out=16'h785;
17'h14628:	data_out=16'h4ef;
17'h14629:	data_out=16'ha00;
17'h1462a:	data_out=16'h85e5;
17'h1462b:	data_out=16'h9d2;
17'h1462c:	data_out=16'h89fd;
17'h1462d:	data_out=16'h9de;
17'h1462e:	data_out=16'h98c;
17'h1462f:	data_out=16'hb3;
17'h14630:	data_out=16'h8a00;
17'h14631:	data_out=16'h9f3;
17'h14632:	data_out=16'h89d0;
17'h14633:	data_out=16'h24d;
17'h14634:	data_out=16'h9fe;
17'h14635:	data_out=16'h898d;
17'h14636:	data_out=16'h121;
17'h14637:	data_out=16'h9f8;
17'h14638:	data_out=16'h9f7;
17'h14639:	data_out=16'h288;
17'h1463a:	data_out=16'h89ff;
17'h1463b:	data_out=16'h89db;
17'h1463c:	data_out=16'ha00;
17'h1463d:	data_out=16'h587;
17'h1463e:	data_out=16'h4f9;
17'h1463f:	data_out=16'hb6;
17'h14640:	data_out=16'h89f7;
17'h14641:	data_out=16'h81de;
17'h14642:	data_out=16'h89c1;
17'h14643:	data_out=16'h8f6;
17'h14644:	data_out=16'h827d;
17'h14645:	data_out=16'h89ea;
17'h14646:	data_out=16'ha00;
17'h14647:	data_out=16'h8a00;
17'h14648:	data_out=16'h8a00;
17'h14649:	data_out=16'h8903;
17'h1464a:	data_out=16'h89e7;
17'h1464b:	data_out=16'h8a00;
17'h1464c:	data_out=16'h89fe;
17'h1464d:	data_out=16'h89ca;
17'h1464e:	data_out=16'h675;
17'h1464f:	data_out=16'h89fe;
17'h14650:	data_out=16'h8a00;
17'h14651:	data_out=16'h8a00;
17'h14652:	data_out=16'h89ed;
17'h14653:	data_out=16'h9fc;
17'h14654:	data_out=16'h99b;
17'h14655:	data_out=16'h8384;
17'h14656:	data_out=16'h80d0;
17'h14657:	data_out=16'h37b;
17'h14658:	data_out=16'h8814;
17'h14659:	data_out=16'h89a9;
17'h1465a:	data_out=16'h68c;
17'h1465b:	data_out=16'ha00;
17'h1465c:	data_out=16'h99a;
17'h1465d:	data_out=16'h88df;
17'h1465e:	data_out=16'h8224;
17'h1465f:	data_out=16'h8940;
17'h14660:	data_out=16'h745;
17'h14661:	data_out=16'h442;
17'h14662:	data_out=16'h9d4;
17'h14663:	data_out=16'h2fd;
17'h14664:	data_out=16'h9ff;
17'h14665:	data_out=16'h89fa;
17'h14666:	data_out=16'h8a00;
17'h14667:	data_out=16'h859a;
17'h14668:	data_out=16'h505;
17'h14669:	data_out=16'h855f;
17'h1466a:	data_out=16'h7af;
17'h1466b:	data_out=16'h89e4;
17'h1466c:	data_out=16'h98d;
17'h1466d:	data_out=16'h33c;
17'h1466e:	data_out=16'h7ac;
17'h1466f:	data_out=16'h8a00;
17'h14670:	data_out=16'h744;
17'h14671:	data_out=16'h8a00;
17'h14672:	data_out=16'h8962;
17'h14673:	data_out=16'h61a;
17'h14674:	data_out=16'h89ff;
17'h14675:	data_out=16'h301;
17'h14676:	data_out=16'h9b6;
17'h14677:	data_out=16'h8a00;
17'h14678:	data_out=16'h89fe;
17'h14679:	data_out=16'h89e0;
17'h1467a:	data_out=16'h319;
17'h1467b:	data_out=16'h4fc;
17'h1467c:	data_out=16'h89f7;
17'h1467d:	data_out=16'h89ff;
17'h1467e:	data_out=16'h9ee;
17'h1467f:	data_out=16'h8a00;
17'h14680:	data_out=16'h9b5;
17'h14681:	data_out=16'ha00;
17'h14682:	data_out=16'h9e5;
17'h14683:	data_out=16'h899b;
17'h14684:	data_out=16'h88c1;
17'h14685:	data_out=16'h6dc;
17'h14686:	data_out=16'h8a00;
17'h14687:	data_out=16'h8a00;
17'h14688:	data_out=16'h9bc;
17'h14689:	data_out=16'h8a00;
17'h1468a:	data_out=16'h8a2;
17'h1468b:	data_out=16'h9e4;
17'h1468c:	data_out=16'h8a00;
17'h1468d:	data_out=16'h8a00;
17'h1468e:	data_out=16'ha00;
17'h1468f:	data_out=16'h950;
17'h14690:	data_out=16'h89fc;
17'h14691:	data_out=16'ha00;
17'h14692:	data_out=16'h82d0;
17'h14693:	data_out=16'h80bf;
17'h14694:	data_out=16'h828d;
17'h14695:	data_out=16'h89f2;
17'h14696:	data_out=16'h89fd;
17'h14697:	data_out=16'h822d;
17'h14698:	data_out=16'h8a00;
17'h14699:	data_out=16'h8984;
17'h1469a:	data_out=16'h892a;
17'h1469b:	data_out=16'h9f5;
17'h1469c:	data_out=16'h873;
17'h1469d:	data_out=16'ha00;
17'h1469e:	data_out=16'h628;
17'h1469f:	data_out=16'h897c;
17'h146a0:	data_out=16'h9b9;
17'h146a1:	data_out=16'ha00;
17'h146a2:	data_out=16'h8740;
17'h146a3:	data_out=16'h7be;
17'h146a4:	data_out=16'h79b;
17'h146a5:	data_out=16'h86f1;
17'h146a6:	data_out=16'h9fb;
17'h146a7:	data_out=16'h9fb;
17'h146a8:	data_out=16'ha00;
17'h146a9:	data_out=16'ha00;
17'h146aa:	data_out=16'h97f;
17'h146ab:	data_out=16'h9ce;
17'h146ac:	data_out=16'h89fd;
17'h146ad:	data_out=16'h9f5;
17'h146ae:	data_out=16'h9da;
17'h146af:	data_out=16'h9c5;
17'h146b0:	data_out=16'h8157;
17'h146b1:	data_out=16'ha00;
17'h146b2:	data_out=16'h97a;
17'h146b3:	data_out=16'h8609;
17'h146b4:	data_out=16'ha00;
17'h146b5:	data_out=16'h367;
17'h146b6:	data_out=16'h9f2;
17'h146b7:	data_out=16'h9f8;
17'h146b8:	data_out=16'ha00;
17'h146b9:	data_out=16'h8604;
17'h146ba:	data_out=16'h89ff;
17'h146bb:	data_out=16'h3ae;
17'h146bc:	data_out=16'ha00;
17'h146bd:	data_out=16'h986;
17'h146be:	data_out=16'ha00;
17'h146bf:	data_out=16'h6d0;
17'h146c0:	data_out=16'h87d7;
17'h146c1:	data_out=16'h335;
17'h146c2:	data_out=16'h8298;
17'h146c3:	data_out=16'h9db;
17'h146c4:	data_out=16'h532;
17'h146c5:	data_out=16'h89f3;
17'h146c6:	data_out=16'ha00;
17'h146c7:	data_out=16'h8a00;
17'h146c8:	data_out=16'h8a00;
17'h146c9:	data_out=16'h85fa;
17'h146ca:	data_out=16'h8799;
17'h146cb:	data_out=16'h41;
17'h146cc:	data_out=16'h89fa;
17'h146cd:	data_out=16'h88a8;
17'h146ce:	data_out=16'h9dc;
17'h146cf:	data_out=16'h8986;
17'h146d0:	data_out=16'h8a00;
17'h146d1:	data_out=16'h89ff;
17'h146d2:	data_out=16'h883d;
17'h146d3:	data_out=16'h9fe;
17'h146d4:	data_out=16'h9af;
17'h146d5:	data_out=16'h372;
17'h146d6:	data_out=16'h9f7;
17'h146d7:	data_out=16'h9ed;
17'h146d8:	data_out=16'h88f0;
17'h146d9:	data_out=16'h83e6;
17'h146da:	data_out=16'h71c;
17'h146db:	data_out=16'ha00;
17'h146dc:	data_out=16'h9ff;
17'h146dd:	data_out=16'h990;
17'h146de:	data_out=16'ha00;
17'h146df:	data_out=16'h86a2;
17'h146e0:	data_out=16'h9f6;
17'h146e1:	data_out=16'ha00;
17'h146e2:	data_out=16'h9f4;
17'h146e3:	data_out=16'hc8;
17'h146e4:	data_out=16'h9fb;
17'h146e5:	data_out=16'h810f;
17'h146e6:	data_out=16'h89ee;
17'h146e7:	data_out=16'hd6;
17'h146e8:	data_out=16'ha00;
17'h146e9:	data_out=16'h163;
17'h146ea:	data_out=16'ha00;
17'h146eb:	data_out=16'h88dd;
17'h146ec:	data_out=16'h989;
17'h146ed:	data_out=16'h45;
17'h146ee:	data_out=16'ha00;
17'h146ef:	data_out=16'h89fa;
17'h146f0:	data_out=16'ha00;
17'h146f1:	data_out=16'h482;
17'h146f2:	data_out=16'h868;
17'h146f3:	data_out=16'ha00;
17'h146f4:	data_out=16'h804f;
17'h146f5:	data_out=16'h760;
17'h146f6:	data_out=16'h667;
17'h146f7:	data_out=16'h89ff;
17'h146f8:	data_out=16'h891e;
17'h146f9:	data_out=16'h80b0;
17'h146fa:	data_out=16'h5e7;
17'h146fb:	data_out=16'ha00;
17'h146fc:	data_out=16'h89fe;
17'h146fd:	data_out=16'h89f8;
17'h146fe:	data_out=16'h9fa;
17'h146ff:	data_out=16'h8a00;
17'h14700:	data_out=16'h68c;
17'h14701:	data_out=16'ha00;
17'h14702:	data_out=16'h9fa;
17'h14703:	data_out=16'h89fc;
17'h14704:	data_out=16'h882e;
17'h14705:	data_out=16'h45c;
17'h14706:	data_out=16'h8a00;
17'h14707:	data_out=16'h8a00;
17'h14708:	data_out=16'h9f2;
17'h14709:	data_out=16'h89fa;
17'h1470a:	data_out=16'h8fa;
17'h1470b:	data_out=16'h9f6;
17'h1470c:	data_out=16'h89d9;
17'h1470d:	data_out=16'h8a00;
17'h1470e:	data_out=16'ha00;
17'h1470f:	data_out=16'h9eb;
17'h14710:	data_out=16'h89fa;
17'h14711:	data_out=16'ha00;
17'h14712:	data_out=16'h861a;
17'h14713:	data_out=16'h897f;
17'h14714:	data_out=16'h89be;
17'h14715:	data_out=16'h89f4;
17'h14716:	data_out=16'h89f7;
17'h14717:	data_out=16'h89f3;
17'h14718:	data_out=16'h8a00;
17'h14719:	data_out=16'h88cb;
17'h1471a:	data_out=16'h880c;
17'h1471b:	data_out=16'h9f7;
17'h1471c:	data_out=16'h6c8;
17'h1471d:	data_out=16'ha00;
17'h1471e:	data_out=16'h81df;
17'h1471f:	data_out=16'h87f7;
17'h14720:	data_out=16'h866e;
17'h14721:	data_out=16'ha00;
17'h14722:	data_out=16'h878d;
17'h14723:	data_out=16'h5f7;
17'h14724:	data_out=16'h5ea;
17'h14725:	data_out=16'h8464;
17'h14726:	data_out=16'ha00;
17'h14727:	data_out=16'h9fd;
17'h14728:	data_out=16'ha00;
17'h14729:	data_out=16'ha00;
17'h1472a:	data_out=16'h9f0;
17'h1472b:	data_out=16'h5e5;
17'h1472c:	data_out=16'h89fa;
17'h1472d:	data_out=16'ha00;
17'h1472e:	data_out=16'ha00;
17'h1472f:	data_out=16'h84af;
17'h14730:	data_out=16'hf9;
17'h14731:	data_out=16'ha00;
17'h14732:	data_out=16'ha00;
17'h14733:	data_out=16'h89fc;
17'h14734:	data_out=16'ha00;
17'h14735:	data_out=16'h9fe;
17'h14736:	data_out=16'h9fc;
17'h14737:	data_out=16'ha00;
17'h14738:	data_out=16'ha00;
17'h14739:	data_out=16'h8a00;
17'h1473a:	data_out=16'h89fb;
17'h1473b:	data_out=16'h9fa;
17'h1473c:	data_out=16'ha00;
17'h1473d:	data_out=16'h82f1;
17'h1473e:	data_out=16'ha00;
17'h1473f:	data_out=16'h422;
17'h14740:	data_out=16'h8599;
17'h14741:	data_out=16'h835;
17'h14742:	data_out=16'h9ec;
17'h14743:	data_out=16'h9ec;
17'h14744:	data_out=16'h938;
17'h14745:	data_out=16'h89f4;
17'h14746:	data_out=16'ha00;
17'h14747:	data_out=16'h89fd;
17'h14748:	data_out=16'h89ff;
17'h14749:	data_out=16'h833b;
17'h1474a:	data_out=16'h85fd;
17'h1474b:	data_out=16'h808c;
17'h1474c:	data_out=16'h8941;
17'h1474d:	data_out=16'h895e;
17'h1474e:	data_out=16'h9f6;
17'h1474f:	data_out=16'h8826;
17'h14750:	data_out=16'h8a00;
17'h14751:	data_out=16'h8769;
17'h14752:	data_out=16'hf9;
17'h14753:	data_out=16'ha00;
17'h14754:	data_out=16'h9db;
17'h14755:	data_out=16'h9f9;
17'h14756:	data_out=16'ha00;
17'h14757:	data_out=16'ha00;
17'h14758:	data_out=16'h547;
17'h14759:	data_out=16'h82ec;
17'h1475a:	data_out=16'h90f;
17'h1475b:	data_out=16'h9fe;
17'h1475c:	data_out=16'h9ff;
17'h1475d:	data_out=16'h9de;
17'h1475e:	data_out=16'h85b9;
17'h1475f:	data_out=16'h8957;
17'h14760:	data_out=16'h9fc;
17'h14761:	data_out=16'ha00;
17'h14762:	data_out=16'h9ff;
17'h14763:	data_out=16'h89e3;
17'h14764:	data_out=16'h9f0;
17'h14765:	data_out=16'h829e;
17'h14766:	data_out=16'h8991;
17'h14767:	data_out=16'h17c;
17'h14768:	data_out=16'ha00;
17'h14769:	data_out=16'h9df;
17'h1476a:	data_out=16'ha00;
17'h1476b:	data_out=16'h8997;
17'h1476c:	data_out=16'h9b4;
17'h1476d:	data_out=16'h89e9;
17'h1476e:	data_out=16'ha00;
17'h1476f:	data_out=16'h899a;
17'h14770:	data_out=16'ha00;
17'h14771:	data_out=16'h9ed;
17'h14772:	data_out=16'h842d;
17'h14773:	data_out=16'ha00;
17'h14774:	data_out=16'h2ad;
17'h14775:	data_out=16'h9f9;
17'h14776:	data_out=16'h9f9;
17'h14777:	data_out=16'h89e9;
17'h14778:	data_out=16'h841f;
17'h14779:	data_out=16'h4e8;
17'h1477a:	data_out=16'h85d8;
17'h1477b:	data_out=16'ha00;
17'h1477c:	data_out=16'h89fe;
17'h1477d:	data_out=16'h89f4;
17'h1477e:	data_out=16'ha00;
17'h1477f:	data_out=16'h8a00;
17'h14780:	data_out=16'h830b;
17'h14781:	data_out=16'ha00;
17'h14782:	data_out=16'ha00;
17'h14783:	data_out=16'h89f4;
17'h14784:	data_out=16'h8871;
17'h14785:	data_out=16'h87bb;
17'h14786:	data_out=16'h8a00;
17'h14787:	data_out=16'h873a;
17'h14788:	data_out=16'h9fc;
17'h14789:	data_out=16'h89f9;
17'h1478a:	data_out=16'h9ff;
17'h1478b:	data_out=16'h9f9;
17'h1478c:	data_out=16'h88bc;
17'h1478d:	data_out=16'h8a00;
17'h1478e:	data_out=16'ha00;
17'h1478f:	data_out=16'ha00;
17'h14790:	data_out=16'h89f5;
17'h14791:	data_out=16'ha00;
17'h14792:	data_out=16'h89f6;
17'h14793:	data_out=16'h89e3;
17'h14794:	data_out=16'h89c4;
17'h14795:	data_out=16'h89f5;
17'h14796:	data_out=16'h89f7;
17'h14797:	data_out=16'h89ca;
17'h14798:	data_out=16'h89fe;
17'h14799:	data_out=16'h876c;
17'h1479a:	data_out=16'h8751;
17'h1479b:	data_out=16'h9fc;
17'h1479c:	data_out=16'h86f6;
17'h1479d:	data_out=16'ha00;
17'h1479e:	data_out=16'h88da;
17'h1479f:	data_out=16'h86e4;
17'h147a0:	data_out=16'h897e;
17'h147a1:	data_out=16'ha00;
17'h147a2:	data_out=16'h88a3;
17'h147a3:	data_out=16'h9f3;
17'h147a4:	data_out=16'h9f3;
17'h147a5:	data_out=16'h8439;
17'h147a6:	data_out=16'ha00;
17'h147a7:	data_out=16'h9ff;
17'h147a8:	data_out=16'ha00;
17'h147a9:	data_out=16'ha00;
17'h147aa:	data_out=16'ha00;
17'h147ab:	data_out=16'h8268;
17'h147ac:	data_out=16'h89fc;
17'h147ad:	data_out=16'ha00;
17'h147ae:	data_out=16'ha00;
17'h147af:	data_out=16'h8918;
17'h147b0:	data_out=16'h790;
17'h147b1:	data_out=16'ha00;
17'h147b2:	data_out=16'ha00;
17'h147b3:	data_out=16'h89ec;
17'h147b4:	data_out=16'ha00;
17'h147b5:	data_out=16'h9fe;
17'h147b6:	data_out=16'ha00;
17'h147b7:	data_out=16'ha00;
17'h147b8:	data_out=16'h9ff;
17'h147b9:	data_out=16'h89f6;
17'h147ba:	data_out=16'h89fa;
17'h147bb:	data_out=16'h9fa;
17'h147bc:	data_out=16'ha00;
17'h147bd:	data_out=16'h867d;
17'h147be:	data_out=16'ha00;
17'h147bf:	data_out=16'h87c1;
17'h147c0:	data_out=16'h8401;
17'h147c1:	data_out=16'h8fb;
17'h147c2:	data_out=16'h9f3;
17'h147c3:	data_out=16'h9f6;
17'h147c4:	data_out=16'h9fb;
17'h147c5:	data_out=16'h89f5;
17'h147c6:	data_out=16'ha00;
17'h147c7:	data_out=16'h89e7;
17'h147c8:	data_out=16'h89ff;
17'h147c9:	data_out=16'h82c2;
17'h147ca:	data_out=16'h8307;
17'h147cb:	data_out=16'h6b2;
17'h147cc:	data_out=16'h88f9;
17'h147cd:	data_out=16'h89d0;
17'h147ce:	data_out=16'h9fb;
17'h147cf:	data_out=16'h8713;
17'h147d0:	data_out=16'h89ff;
17'h147d1:	data_out=16'h89ff;
17'h147d2:	data_out=16'h9f4;
17'h147d3:	data_out=16'ha00;
17'h147d4:	data_out=16'h8740;
17'h147d5:	data_out=16'h519;
17'h147d6:	data_out=16'h9ff;
17'h147d7:	data_out=16'ha00;
17'h147d8:	data_out=16'h801;
17'h147d9:	data_out=16'h826f;
17'h147da:	data_out=16'h968;
17'h147db:	data_out=16'h9fd;
17'h147dc:	data_out=16'h9fe;
17'h147dd:	data_out=16'h2a4;
17'h147de:	data_out=16'h8770;
17'h147df:	data_out=16'h89ac;
17'h147e0:	data_out=16'h9ff;
17'h147e1:	data_out=16'h9ff;
17'h147e2:	data_out=16'h8e3;
17'h147e3:	data_out=16'h89da;
17'h147e4:	data_out=16'h9f1;
17'h147e5:	data_out=16'ha00;
17'h147e6:	data_out=16'h8999;
17'h147e7:	data_out=16'h9da;
17'h147e8:	data_out=16'ha00;
17'h147e9:	data_out=16'h9b3;
17'h147ea:	data_out=16'ha00;
17'h147eb:	data_out=16'h8982;
17'h147ec:	data_out=16'h4b9;
17'h147ed:	data_out=16'h89db;
17'h147ee:	data_out=16'ha00;
17'h147ef:	data_out=16'h8970;
17'h147f0:	data_out=16'ha00;
17'h147f1:	data_out=16'h9ff;
17'h147f2:	data_out=16'h8445;
17'h147f3:	data_out=16'ha00;
17'h147f4:	data_out=16'h87e;
17'h147f5:	data_out=16'h9dc;
17'h147f6:	data_out=16'h9fa;
17'h147f7:	data_out=16'h89bc;
17'h147f8:	data_out=16'h52b;
17'h147f9:	data_out=16'h705;
17'h147fa:	data_out=16'h89b2;
17'h147fb:	data_out=16'ha00;
17'h147fc:	data_out=16'h89fa;
17'h147fd:	data_out=16'h89e4;
17'h147fe:	data_out=16'ha00;
17'h147ff:	data_out=16'h8a00;
17'h14800:	data_out=16'h640;
17'h14801:	data_out=16'ha00;
17'h14802:	data_out=16'ha00;
17'h14803:	data_out=16'h89e9;
17'h14804:	data_out=16'h8969;
17'h14805:	data_out=16'h87c4;
17'h14806:	data_out=16'h8a00;
17'h14807:	data_out=16'h233;
17'h14808:	data_out=16'h9f8;
17'h14809:	data_out=16'h89f0;
17'h1480a:	data_out=16'h9ed;
17'h1480b:	data_out=16'h210;
17'h1480c:	data_out=16'h84d5;
17'h1480d:	data_out=16'h8a00;
17'h1480e:	data_out=16'ha00;
17'h1480f:	data_out=16'h9ff;
17'h14810:	data_out=16'h89e9;
17'h14811:	data_out=16'ha00;
17'h14812:	data_out=16'h89d8;
17'h14813:	data_out=16'h89f7;
17'h14814:	data_out=16'h89b3;
17'h14815:	data_out=16'h89f3;
17'h14816:	data_out=16'h89ef;
17'h14817:	data_out=16'h89c2;
17'h14818:	data_out=16'h89f6;
17'h14819:	data_out=16'h14;
17'h1481a:	data_out=16'h88da;
17'h1481b:	data_out=16'h9fc;
17'h1481c:	data_out=16'h89e7;
17'h1481d:	data_out=16'ha00;
17'h1481e:	data_out=16'h8956;
17'h1481f:	data_out=16'h882f;
17'h14820:	data_out=16'h89b0;
17'h14821:	data_out=16'ha00;
17'h14822:	data_out=16'h8952;
17'h14823:	data_out=16'h9e7;
17'h14824:	data_out=16'h9e7;
17'h14825:	data_out=16'h8662;
17'h14826:	data_out=16'ha00;
17'h14827:	data_out=16'h9fd;
17'h14828:	data_out=16'ha00;
17'h14829:	data_out=16'ha00;
17'h1482a:	data_out=16'ha00;
17'h1482b:	data_out=16'h8964;
17'h1482c:	data_out=16'h89f7;
17'h1482d:	data_out=16'ha00;
17'h1482e:	data_out=16'ha00;
17'h1482f:	data_out=16'h89bb;
17'h14830:	data_out=16'h9c8;
17'h14831:	data_out=16'h9fd;
17'h14832:	data_out=16'h9e0;
17'h14833:	data_out=16'h89ca;
17'h14834:	data_out=16'ha00;
17'h14835:	data_out=16'h9fd;
17'h14836:	data_out=16'h9fd;
17'h14837:	data_out=16'ha00;
17'h14838:	data_out=16'h818b;
17'h14839:	data_out=16'h89d2;
17'h1483a:	data_out=16'h89e3;
17'h1483b:	data_out=16'h9c4;
17'h1483c:	data_out=16'h9fd;
17'h1483d:	data_out=16'h88e1;
17'h1483e:	data_out=16'ha00;
17'h1483f:	data_out=16'h87c5;
17'h14840:	data_out=16'h8618;
17'h14841:	data_out=16'h9b1;
17'h14842:	data_out=16'h9e7;
17'h14843:	data_out=16'ha00;
17'h14844:	data_out=16'h9ee;
17'h14845:	data_out=16'h89f5;
17'h14846:	data_out=16'h9ff;
17'h14847:	data_out=16'h89ca;
17'h14848:	data_out=16'h8a00;
17'h14849:	data_out=16'h858b;
17'h1484a:	data_out=16'h859b;
17'h1484b:	data_out=16'h86c6;
17'h1484c:	data_out=16'h8850;
17'h1484d:	data_out=16'h89e9;
17'h1484e:	data_out=16'h9fb;
17'h1484f:	data_out=16'h8702;
17'h14850:	data_out=16'h8a00;
17'h14851:	data_out=16'h89d8;
17'h14852:	data_out=16'h9e1;
17'h14853:	data_out=16'h9fe;
17'h14854:	data_out=16'h8996;
17'h14855:	data_out=16'h81ec;
17'h14856:	data_out=16'h9fc;
17'h14857:	data_out=16'h9ff;
17'h14858:	data_out=16'h6c8;
17'h14859:	data_out=16'h3aa;
17'h1485a:	data_out=16'h98f;
17'h1485b:	data_out=16'h9fb;
17'h1485c:	data_out=16'h9fd;
17'h1485d:	data_out=16'h82eb;
17'h1485e:	data_out=16'h87e4;
17'h1485f:	data_out=16'h89ba;
17'h14860:	data_out=16'ha00;
17'h14861:	data_out=16'h9e0;
17'h14862:	data_out=16'h83ae;
17'h14863:	data_out=16'h89c2;
17'h14864:	data_out=16'h9ef;
17'h14865:	data_out=16'h814a;
17'h14866:	data_out=16'h8999;
17'h14867:	data_out=16'ha00;
17'h14868:	data_out=16'ha00;
17'h14869:	data_out=16'h9b0;
17'h1486a:	data_out=16'ha00;
17'h1486b:	data_out=16'h89b6;
17'h1486c:	data_out=16'h9ee;
17'h1486d:	data_out=16'h89c3;
17'h1486e:	data_out=16'ha00;
17'h1486f:	data_out=16'h8937;
17'h14870:	data_out=16'ha00;
17'h14871:	data_out=16'h9fe;
17'h14872:	data_out=16'h819a;
17'h14873:	data_out=16'h9ea;
17'h14874:	data_out=16'h9c2;
17'h14875:	data_out=16'h9a8;
17'h14876:	data_out=16'h9fd;
17'h14877:	data_out=16'h89ce;
17'h14878:	data_out=16'h9d4;
17'h14879:	data_out=16'h611;
17'h1487a:	data_out=16'h89b4;
17'h1487b:	data_out=16'ha00;
17'h1487c:	data_out=16'h89f7;
17'h1487d:	data_out=16'h89d4;
17'h1487e:	data_out=16'h37b;
17'h1487f:	data_out=16'h8a00;
17'h14880:	data_out=16'h32a;
17'h14881:	data_out=16'ha00;
17'h14882:	data_out=16'h9fe;
17'h14883:	data_out=16'h89ce;
17'h14884:	data_out=16'h8a00;
17'h14885:	data_out=16'h8760;
17'h14886:	data_out=16'h8a00;
17'h14887:	data_out=16'h6f0;
17'h14888:	data_out=16'h9e2;
17'h14889:	data_out=16'h89c6;
17'h1488a:	data_out=16'h9b5;
17'h1488b:	data_out=16'h8688;
17'h1488c:	data_out=16'h9b7;
17'h1488d:	data_out=16'h8a00;
17'h1488e:	data_out=16'ha00;
17'h1488f:	data_out=16'h9fe;
17'h14890:	data_out=16'h8a00;
17'h14891:	data_out=16'ha00;
17'h14892:	data_out=16'h89aa;
17'h14893:	data_out=16'h8a00;
17'h14894:	data_out=16'h897d;
17'h14895:	data_out=16'h89fe;
17'h14896:	data_out=16'h89f2;
17'h14897:	data_out=16'h8977;
17'h14898:	data_out=16'h89f4;
17'h14899:	data_out=16'h9ca;
17'h1489a:	data_out=16'h89c6;
17'h1489b:	data_out=16'h8844;
17'h1489c:	data_out=16'h89eb;
17'h1489d:	data_out=16'ha00;
17'h1489e:	data_out=16'h8999;
17'h1489f:	data_out=16'h88c7;
17'h148a0:	data_out=16'h89db;
17'h148a1:	data_out=16'ha00;
17'h148a2:	data_out=16'h89db;
17'h148a3:	data_out=16'h8c4;
17'h148a4:	data_out=16'h8ab;
17'h148a5:	data_out=16'h8960;
17'h148a6:	data_out=16'h9fe;
17'h148a7:	data_out=16'h9d0;
17'h148a8:	data_out=16'ha00;
17'h148a9:	data_out=16'ha00;
17'h148aa:	data_out=16'ha00;
17'h148ab:	data_out=16'h89c6;
17'h148ac:	data_out=16'h89fa;
17'h148ad:	data_out=16'ha00;
17'h148ae:	data_out=16'ha00;
17'h148af:	data_out=16'h89da;
17'h148b0:	data_out=16'h9d0;
17'h148b1:	data_out=16'h9cf;
17'h148b2:	data_out=16'h9a5;
17'h148b3:	data_out=16'h89ad;
17'h148b4:	data_out=16'ha00;
17'h148b5:	data_out=16'h9f3;
17'h148b6:	data_out=16'h81e5;
17'h148b7:	data_out=16'ha00;
17'h148b8:	data_out=16'h89f8;
17'h148b9:	data_out=16'h89c1;
17'h148ba:	data_out=16'h89e2;
17'h148bb:	data_out=16'h714;
17'h148bc:	data_out=16'h9f8;
17'h148bd:	data_out=16'h89e2;
17'h148be:	data_out=16'ha00;
17'h148bf:	data_out=16'h8746;
17'h148c0:	data_out=16'h89d3;
17'h148c1:	data_out=16'h8306;
17'h148c2:	data_out=16'h9cb;
17'h148c3:	data_out=16'ha00;
17'h148c4:	data_out=16'h96d;
17'h148c5:	data_out=16'h89fd;
17'h148c6:	data_out=16'ha00;
17'h148c7:	data_out=16'h89b3;
17'h148c8:	data_out=16'h8a00;
17'h148c9:	data_out=16'h8970;
17'h148ca:	data_out=16'h82a8;
17'h148cb:	data_out=16'h8471;
17'h148cc:	data_out=16'h895d;
17'h148cd:	data_out=16'h89fe;
17'h148ce:	data_out=16'h662;
17'h148cf:	data_out=16'h8909;
17'h148d0:	data_out=16'h8a00;
17'h148d1:	data_out=16'h89a1;
17'h148d2:	data_out=16'h9be;
17'h148d3:	data_out=16'h9ff;
17'h148d4:	data_out=16'h89c2;
17'h148d5:	data_out=16'h84e3;
17'h148d6:	data_out=16'h9dd;
17'h148d7:	data_out=16'h255;
17'h148d8:	data_out=16'h28d;
17'h148d9:	data_out=16'h89ce;
17'h148da:	data_out=16'h9f2;
17'h148db:	data_out=16'h804;
17'h148dc:	data_out=16'h9f8;
17'h148dd:	data_out=16'h8955;
17'h148de:	data_out=16'h8973;
17'h148df:	data_out=16'h89ed;
17'h148e0:	data_out=16'h9ff;
17'h148e1:	data_out=16'h9ad;
17'h148e2:	data_out=16'h84f1;
17'h148e3:	data_out=16'h89a3;
17'h148e4:	data_out=16'h98e;
17'h148e5:	data_out=16'h84aa;
17'h148e6:	data_out=16'h916;
17'h148e7:	data_out=16'ha00;
17'h148e8:	data_out=16'ha00;
17'h148e9:	data_out=16'h818f;
17'h148ea:	data_out=16'ha00;
17'h148eb:	data_out=16'h89f6;
17'h148ec:	data_out=16'h9dd;
17'h148ed:	data_out=16'h89a6;
17'h148ee:	data_out=16'ha00;
17'h148ef:	data_out=16'h87fc;
17'h148f0:	data_out=16'ha00;
17'h148f1:	data_out=16'h80ff;
17'h148f2:	data_out=16'h877a;
17'h148f3:	data_out=16'h9b7;
17'h148f4:	data_out=16'h9be;
17'h148f5:	data_out=16'h996;
17'h148f6:	data_out=16'h475;
17'h148f7:	data_out=16'h89c5;
17'h148f8:	data_out=16'h9bc;
17'h148f9:	data_out=16'h82e6;
17'h148fa:	data_out=16'h8993;
17'h148fb:	data_out=16'ha00;
17'h148fc:	data_out=16'h89f5;
17'h148fd:	data_out=16'h89d5;
17'h148fe:	data_out=16'h849e;
17'h148ff:	data_out=16'h8a00;
17'h14900:	data_out=16'h9d2;
17'h14901:	data_out=16'ha00;
17'h14902:	data_out=16'h9fa;
17'h14903:	data_out=16'h89c5;
17'h14904:	data_out=16'h8a00;
17'h14905:	data_out=16'h89dc;
17'h14906:	data_out=16'h8a00;
17'h14907:	data_out=16'h9eb;
17'h14908:	data_out=16'h9a7;
17'h14909:	data_out=16'h89ba;
17'h1490a:	data_out=16'h9a6;
17'h1490b:	data_out=16'h88ef;
17'h1490c:	data_out=16'h9c2;
17'h1490d:	data_out=16'h89d5;
17'h1490e:	data_out=16'h9ff;
17'h1490f:	data_out=16'h9fe;
17'h14910:	data_out=16'h8a00;
17'h14911:	data_out=16'h635;
17'h14912:	data_out=16'h8968;
17'h14913:	data_out=16'h8a00;
17'h14914:	data_out=16'h8965;
17'h14915:	data_out=16'h89e9;
17'h14916:	data_out=16'h89c0;
17'h14917:	data_out=16'h8946;
17'h14918:	data_out=16'h89e2;
17'h14919:	data_out=16'h72d;
17'h1491a:	data_out=16'h89fb;
17'h1491b:	data_out=16'h8944;
17'h1491c:	data_out=16'h89e9;
17'h1491d:	data_out=16'h9ff;
17'h1491e:	data_out=16'h896b;
17'h1491f:	data_out=16'h88f1;
17'h14920:	data_out=16'h89cd;
17'h14921:	data_out=16'h9fe;
17'h14922:	data_out=16'h8a00;
17'h14923:	data_out=16'h4d1;
17'h14924:	data_out=16'h4b1;
17'h14925:	data_out=16'h89df;
17'h14926:	data_out=16'h9d9;
17'h14927:	data_out=16'h15a;
17'h14928:	data_out=16'h9fe;
17'h14929:	data_out=16'ha00;
17'h1492a:	data_out=16'ha00;
17'h1492b:	data_out=16'h89fd;
17'h1492c:	data_out=16'h89c6;
17'h1492d:	data_out=16'ha00;
17'h1492e:	data_out=16'ha00;
17'h1492f:	data_out=16'h89e6;
17'h14930:	data_out=16'h9be;
17'h14931:	data_out=16'h9c4;
17'h14932:	data_out=16'hcf;
17'h14933:	data_out=16'h8999;
17'h14934:	data_out=16'ha00;
17'h14935:	data_out=16'h89b4;
17'h14936:	data_out=16'h84a2;
17'h14937:	data_out=16'ha00;
17'h14938:	data_out=16'h8a00;
17'h14939:	data_out=16'h89af;
17'h1493a:	data_out=16'h89d4;
17'h1493b:	data_out=16'h8317;
17'h1493c:	data_out=16'h9ad;
17'h1493d:	data_out=16'h89cc;
17'h1493e:	data_out=16'h9fe;
17'h1493f:	data_out=16'h89dc;
17'h14940:	data_out=16'h8a00;
17'h14941:	data_out=16'h82ee;
17'h14942:	data_out=16'h9a0;
17'h14943:	data_out=16'ha00;
17'h14944:	data_out=16'h4f8;
17'h14945:	data_out=16'h89e7;
17'h14946:	data_out=16'h9d8;
17'h14947:	data_out=16'h8985;
17'h14948:	data_out=16'h89e6;
17'h14949:	data_out=16'h89f8;
17'h1494a:	data_out=16'h4f5;
17'h1494b:	data_out=16'h8232;
17'h1494c:	data_out=16'h89df;
17'h1494d:	data_out=16'h8a00;
17'h1494e:	data_out=16'h61f;
17'h1494f:	data_out=16'h89ce;
17'h14950:	data_out=16'h8a00;
17'h14951:	data_out=16'h88dc;
17'h14952:	data_out=16'h715;
17'h14953:	data_out=16'h8782;
17'h14954:	data_out=16'h89b4;
17'h14955:	data_out=16'h8627;
17'h14956:	data_out=16'h28a;
17'h14957:	data_out=16'h898a;
17'h14958:	data_out=16'hd4;
17'h14959:	data_out=16'h8a00;
17'h1495a:	data_out=16'h8ac;
17'h1495b:	data_out=16'h8234;
17'h1495c:	data_out=16'h8829;
17'h1495d:	data_out=16'h8988;
17'h1495e:	data_out=16'h89b0;
17'h1495f:	data_out=16'h89df;
17'h14960:	data_out=16'h9e6;
17'h14961:	data_out=16'h656;
17'h14962:	data_out=16'h86a1;
17'h14963:	data_out=16'h897e;
17'h14964:	data_out=16'h840a;
17'h14965:	data_out=16'h89b4;
17'h14966:	data_out=16'h9eb;
17'h14967:	data_out=16'ha00;
17'h14968:	data_out=16'h9fe;
17'h14969:	data_out=16'h8576;
17'h1496a:	data_out=16'h9ff;
17'h1496b:	data_out=16'h89dd;
17'h1496c:	data_out=16'h9fa;
17'h1496d:	data_out=16'h8985;
17'h1496e:	data_out=16'h9ff;
17'h1496f:	data_out=16'h8914;
17'h14970:	data_out=16'h9ff;
17'h14971:	data_out=16'h9ff;
17'h14972:	data_out=16'h89e7;
17'h14973:	data_out=16'h42f;
17'h14974:	data_out=16'h99d;
17'h14975:	data_out=16'h43f;
17'h14976:	data_out=16'h126;
17'h14977:	data_out=16'h89da;
17'h14978:	data_out=16'h54b;
17'h14979:	data_out=16'h5bb;
17'h1497a:	data_out=16'h896b;
17'h1497b:	data_out=16'h9fe;
17'h1497c:	data_out=16'h89e6;
17'h1497d:	data_out=16'h89b1;
17'h1497e:	data_out=16'h8829;
17'h1497f:	data_out=16'h8a00;
17'h14980:	data_out=16'h9f3;
17'h14981:	data_out=16'ha00;
17'h14982:	data_out=16'h9f0;
17'h14983:	data_out=16'h899a;
17'h14984:	data_out=16'h89f1;
17'h14985:	data_out=16'h8569;
17'h14986:	data_out=16'h8a00;
17'h14987:	data_out=16'h9b6;
17'h14988:	data_out=16'h12;
17'h14989:	data_out=16'h89cd;
17'h1498a:	data_out=16'h9c3;
17'h1498b:	data_out=16'h89d7;
17'h1498c:	data_out=16'h97c;
17'h1498d:	data_out=16'h89ad;
17'h1498e:	data_out=16'h9fd;
17'h1498f:	data_out=16'h780;
17'h14990:	data_out=16'h8a00;
17'h14991:	data_out=16'h8a00;
17'h14992:	data_out=16'h87ff;
17'h14993:	data_out=16'h89f0;
17'h14994:	data_out=16'h8966;
17'h14995:	data_out=16'h88f6;
17'h14996:	data_out=16'h8112;
17'h14997:	data_out=16'h88f9;
17'h14998:	data_out=16'h890e;
17'h14999:	data_out=16'h80a4;
17'h1499a:	data_out=16'h8987;
17'h1499b:	data_out=16'h8990;
17'h1499c:	data_out=16'h89a6;
17'h1499d:	data_out=16'ha00;
17'h1499e:	data_out=16'h88ae;
17'h1499f:	data_out=16'h881f;
17'h149a0:	data_out=16'h897d;
17'h149a1:	data_out=16'h9fd;
17'h149a2:	data_out=16'h8a00;
17'h149a3:	data_out=16'h8a00;
17'h149a4:	data_out=16'h8a00;
17'h149a5:	data_out=16'h8a00;
17'h149a6:	data_out=16'h8a5;
17'h149a7:	data_out=16'h8674;
17'h149a8:	data_out=16'h9fc;
17'h149a9:	data_out=16'ha00;
17'h149aa:	data_out=16'ha00;
17'h149ab:	data_out=16'h8a00;
17'h149ac:	data_out=16'h83f8;
17'h149ad:	data_out=16'h9fb;
17'h149ae:	data_out=16'ha00;
17'h149af:	data_out=16'h8998;
17'h149b0:	data_out=16'h9ce;
17'h149b1:	data_out=16'h9ef;
17'h149b2:	data_out=16'h63;
17'h149b3:	data_out=16'h8976;
17'h149b4:	data_out=16'ha00;
17'h149b5:	data_out=16'h89b0;
17'h149b6:	data_out=16'h8723;
17'h149b7:	data_out=16'h9fb;
17'h149b8:	data_out=16'h89da;
17'h149b9:	data_out=16'h899b;
17'h149ba:	data_out=16'h89dd;
17'h149bb:	data_out=16'h85ce;
17'h149bc:	data_out=16'h62c;
17'h149bd:	data_out=16'h8963;
17'h149be:	data_out=16'h9fc;
17'h149bf:	data_out=16'h8524;
17'h149c0:	data_out=16'h89f4;
17'h149c1:	data_out=16'h81d5;
17'h149c2:	data_out=16'h88cc;
17'h149c3:	data_out=16'h5dd;
17'h149c4:	data_out=16'h866;
17'h149c5:	data_out=16'h88aa;
17'h149c6:	data_out=16'h9af;
17'h149c7:	data_out=16'h898c;
17'h149c8:	data_out=16'h89b2;
17'h149c9:	data_out=16'h8a00;
17'h149ca:	data_out=16'h5cf;
17'h149cb:	data_out=16'h89b4;
17'h149cc:	data_out=16'h89e4;
17'h149cd:	data_out=16'h8a00;
17'h149ce:	data_out=16'h651;
17'h149cf:	data_out=16'h89f7;
17'h149d0:	data_out=16'h89d4;
17'h149d1:	data_out=16'h8756;
17'h149d2:	data_out=16'h8a00;
17'h149d3:	data_out=16'h8886;
17'h149d4:	data_out=16'h8961;
17'h149d5:	data_out=16'h86f3;
17'h149d6:	data_out=16'h8a00;
17'h149d7:	data_out=16'h89ad;
17'h149d8:	data_out=16'h34;
17'h149d9:	data_out=16'h89fe;
17'h149da:	data_out=16'h4ca;
17'h149db:	data_out=16'h89f7;
17'h149dc:	data_out=16'h886a;
17'h149dd:	data_out=16'h277;
17'h149de:	data_out=16'h8907;
17'h149df:	data_out=16'h8977;
17'h149e0:	data_out=16'h9bd;
17'h149e1:	data_out=16'h8b2;
17'h149e2:	data_out=16'h8812;
17'h149e3:	data_out=16'h895c;
17'h149e4:	data_out=16'h86ec;
17'h149e5:	data_out=16'h89fb;
17'h149e6:	data_out=16'h9fb;
17'h149e7:	data_out=16'ha00;
17'h149e8:	data_out=16'h9fc;
17'h149e9:	data_out=16'h89e5;
17'h149ea:	data_out=16'h9fd;
17'h149eb:	data_out=16'h8963;
17'h149ec:	data_out=16'h9fd;
17'h149ed:	data_out=16'h8963;
17'h149ee:	data_out=16'h9fd;
17'h149ef:	data_out=16'h84f4;
17'h149f0:	data_out=16'h9fd;
17'h149f1:	data_out=16'ha00;
17'h149f2:	data_out=16'h884f;
17'h149f3:	data_out=16'h9e4;
17'h149f4:	data_out=16'h9a5;
17'h149f5:	data_out=16'h708;
17'h149f6:	data_out=16'h86df;
17'h149f7:	data_out=16'h89d6;
17'h149f8:	data_out=16'h5c3;
17'h149f9:	data_out=16'h740;
17'h149fa:	data_out=16'h892f;
17'h149fb:	data_out=16'h9fc;
17'h149fc:	data_out=16'h884d;
17'h149fd:	data_out=16'h8991;
17'h149fe:	data_out=16'h896c;
17'h149ff:	data_out=16'h8a00;
17'h14a00:	data_out=16'h9f9;
17'h14a01:	data_out=16'ha00;
17'h14a02:	data_out=16'h761;
17'h14a03:	data_out=16'h8981;
17'h14a04:	data_out=16'h890a;
17'h14a05:	data_out=16'h9e7;
17'h14a06:	data_out=16'h89fb;
17'h14a07:	data_out=16'h89f8;
17'h14a08:	data_out=16'h89ec;
17'h14a09:	data_out=16'h89fc;
17'h14a0a:	data_out=16'h9e8;
17'h14a0b:	data_out=16'h89f0;
17'h14a0c:	data_out=16'h89fc;
17'h14a0d:	data_out=16'h89b7;
17'h14a0e:	data_out=16'h9ff;
17'h14a0f:	data_out=16'h1c;
17'h14a10:	data_out=16'h8a00;
17'h14a11:	data_out=16'h8a00;
17'h14a12:	data_out=16'h879d;
17'h14a13:	data_out=16'h89eb;
17'h14a14:	data_out=16'h89b1;
17'h14a15:	data_out=16'h9f7;
17'h14a16:	data_out=16'h9bf;
17'h14a17:	data_out=16'h896d;
17'h14a18:	data_out=16'h6c2;
17'h14a19:	data_out=16'h83fe;
17'h14a1a:	data_out=16'h41e;
17'h14a1b:	data_out=16'h89ef;
17'h14a1c:	data_out=16'h8991;
17'h14a1d:	data_out=16'h9ee;
17'h14a1e:	data_out=16'h87b4;
17'h14a1f:	data_out=16'h87fb;
17'h14a20:	data_out=16'h879d;
17'h14a21:	data_out=16'h9ff;
17'h14a22:	data_out=16'h89db;
17'h14a23:	data_out=16'h8a00;
17'h14a24:	data_out=16'h8a00;
17'h14a25:	data_out=16'h89f9;
17'h14a26:	data_out=16'h856f;
17'h14a27:	data_out=16'h89eb;
17'h14a28:	data_out=16'h9ff;
17'h14a29:	data_out=16'ha00;
17'h14a2a:	data_out=16'h80d8;
17'h14a2b:	data_out=16'h8a00;
17'h14a2c:	data_out=16'h9ee;
17'h14a2d:	data_out=16'h2a1;
17'h14a2e:	data_out=16'h8061;
17'h14a2f:	data_out=16'h8840;
17'h14a30:	data_out=16'h9cf;
17'h14a31:	data_out=16'h9e9;
17'h14a32:	data_out=16'h1ff;
17'h14a33:	data_out=16'h8989;
17'h14a34:	data_out=16'h9ff;
17'h14a35:	data_out=16'h8610;
17'h14a36:	data_out=16'h8892;
17'h14a37:	data_out=16'h6ad;
17'h14a38:	data_out=16'h89da;
17'h14a39:	data_out=16'h89a5;
17'h14a3a:	data_out=16'h89f5;
17'h14a3b:	data_out=16'h89dd;
17'h14a3c:	data_out=16'h9df;
17'h14a3d:	data_out=16'h8652;
17'h14a3e:	data_out=16'h9ff;
17'h14a3f:	data_out=16'h9e7;
17'h14a40:	data_out=16'h89b9;
17'h14a41:	data_out=16'h8489;
17'h14a42:	data_out=16'h8a00;
17'h14a43:	data_out=16'h8675;
17'h14a44:	data_out=16'h9d0;
17'h14a45:	data_out=16'h9f7;
17'h14a46:	data_out=16'h9cc;
17'h14a47:	data_out=16'h89ce;
17'h14a48:	data_out=16'h89da;
17'h14a49:	data_out=16'h8a00;
17'h14a4a:	data_out=16'h89ed;
17'h14a4b:	data_out=16'h89fc;
17'h14a4c:	data_out=16'h89dd;
17'h14a4d:	data_out=16'h89de;
17'h14a4e:	data_out=16'h4b9;
17'h14a4f:	data_out=16'h89fb;
17'h14a50:	data_out=16'h8989;
17'h14a51:	data_out=16'h9ed;
17'h14a52:	data_out=16'h8a00;
17'h14a53:	data_out=16'h8960;
17'h14a54:	data_out=16'h87a3;
17'h14a55:	data_out=16'h88b6;
17'h14a56:	data_out=16'h82b3;
17'h14a57:	data_out=16'h89ad;
17'h14a58:	data_out=16'h690;
17'h14a59:	data_out=16'h89a5;
17'h14a5a:	data_out=16'h87a4;
17'h14a5b:	data_out=16'hd6;
17'h14a5c:	data_out=16'h1d3;
17'h14a5d:	data_out=16'ha00;
17'h14a5e:	data_out=16'h883c;
17'h14a5f:	data_out=16'h83f9;
17'h14a60:	data_out=16'h689;
17'h14a61:	data_out=16'h9e5;
17'h14a62:	data_out=16'h8962;
17'h14a63:	data_out=16'h8904;
17'h14a64:	data_out=16'h89c5;
17'h14a65:	data_out=16'h89f5;
17'h14a66:	data_out=16'h9f7;
17'h14a67:	data_out=16'ha00;
17'h14a68:	data_out=16'h9ff;
17'h14a69:	data_out=16'h89fd;
17'h14a6a:	data_out=16'h9ff;
17'h14a6b:	data_out=16'h855a;
17'h14a6c:	data_out=16'h9ff;
17'h14a6d:	data_out=16'h8918;
17'h14a6e:	data_out=16'h9ff;
17'h14a6f:	data_out=16'h81fb;
17'h14a70:	data_out=16'h9ff;
17'h14a71:	data_out=16'ha00;
17'h14a72:	data_out=16'h804;
17'h14a73:	data_out=16'h9f2;
17'h14a74:	data_out=16'h973;
17'h14a75:	data_out=16'h9d9;
17'h14a76:	data_out=16'h8005;
17'h14a77:	data_out=16'h89f0;
17'h14a78:	data_out=16'h89fe;
17'h14a79:	data_out=16'h8b2;
17'h14a7a:	data_out=16'h8926;
17'h14a7b:	data_out=16'h9ff;
17'h14a7c:	data_out=16'h97f;
17'h14a7d:	data_out=16'h86ad;
17'h14a7e:	data_out=16'h89d0;
17'h14a7f:	data_out=16'h81d7;
17'h14a80:	data_out=16'h276;
17'h14a81:	data_out=16'ha00;
17'h14a82:	data_out=16'h3eb;
17'h14a83:	data_out=16'h899f;
17'h14a84:	data_out=16'h842b;
17'h14a85:	data_out=16'h9fa;
17'h14a86:	data_out=16'h89f9;
17'h14a87:	data_out=16'h89ff;
17'h14a88:	data_out=16'h89ee;
17'h14a89:	data_out=16'h89fc;
17'h14a8a:	data_out=16'h9fc;
17'h14a8b:	data_out=16'h89e2;
17'h14a8c:	data_out=16'h8a00;
17'h14a8d:	data_out=16'h89e4;
17'h14a8e:	data_out=16'h9ff;
17'h14a8f:	data_out=16'h8859;
17'h14a90:	data_out=16'h89db;
17'h14a91:	data_out=16'h89d8;
17'h14a92:	data_out=16'h880f;
17'h14a93:	data_out=16'h89db;
17'h14a94:	data_out=16'h86cb;
17'h14a95:	data_out=16'h9fe;
17'h14a96:	data_out=16'h9f4;
17'h14a97:	data_out=16'h8792;
17'h14a98:	data_out=16'h9fa;
17'h14a99:	data_out=16'hb2;
17'h14a9a:	data_out=16'h323;
17'h14a9b:	data_out=16'h89d9;
17'h14a9c:	data_out=16'h898b;
17'h14a9d:	data_out=16'h8419;
17'h14a9e:	data_out=16'h8325;
17'h14a9f:	data_out=16'h8195;
17'h14aa0:	data_out=16'h8531;
17'h14aa1:	data_out=16'h9ff;
17'h14aa2:	data_out=16'h89a1;
17'h14aa3:	data_out=16'h8a00;
17'h14aa4:	data_out=16'h8a00;
17'h14aa5:	data_out=16'h89fa;
17'h14aa6:	data_out=16'h8a00;
17'h14aa7:	data_out=16'h88e6;
17'h14aa8:	data_out=16'h9fe;
17'h14aa9:	data_out=16'ha00;
17'h14aaa:	data_out=16'h87b4;
17'h14aab:	data_out=16'h89f2;
17'h14aac:	data_out=16'h9f9;
17'h14aad:	data_out=16'h8812;
17'h14aae:	data_out=16'h869c;
17'h14aaf:	data_out=16'h86c5;
17'h14ab0:	data_out=16'h5c6;
17'h14ab1:	data_out=16'h9f8;
17'h14ab2:	data_out=16'h89db;
17'h14ab3:	data_out=16'h8717;
17'h14ab4:	data_out=16'h9fe;
17'h14ab5:	data_out=16'h80b6;
17'h14ab6:	data_out=16'h8921;
17'h14ab7:	data_out=16'h4a3;
17'h14ab8:	data_out=16'h8920;
17'h14ab9:	data_out=16'h87d9;
17'h14aba:	data_out=16'h89f6;
17'h14abb:	data_out=16'h89fa;
17'h14abc:	data_out=16'ha00;
17'h14abd:	data_out=16'h8310;
17'h14abe:	data_out=16'h9fe;
17'h14abf:	data_out=16'h9fa;
17'h14ac0:	data_out=16'h88f0;
17'h14ac1:	data_out=16'h8867;
17'h14ac2:	data_out=16'h89ff;
17'h14ac3:	data_out=16'h872a;
17'h14ac4:	data_out=16'h9f3;
17'h14ac5:	data_out=16'h9fe;
17'h14ac6:	data_out=16'h9ea;
17'h14ac7:	data_out=16'h89f2;
17'h14ac8:	data_out=16'h8979;
17'h14ac9:	data_out=16'h89f0;
17'h14aca:	data_out=16'h88cd;
17'h14acb:	data_out=16'h89fe;
17'h14acc:	data_out=16'h89f0;
17'h14acd:	data_out=16'h8948;
17'h14ace:	data_out=16'h89c6;
17'h14acf:	data_out=16'h89ff;
17'h14ad0:	data_out=16'h8884;
17'h14ad1:	data_out=16'h9e1;
17'h14ad2:	data_out=16'h8a00;
17'h14ad3:	data_out=16'h8758;
17'h14ad4:	data_out=16'h85d6;
17'h14ad5:	data_out=16'h403;
17'h14ad6:	data_out=16'h501;
17'h14ad7:	data_out=16'h65d;
17'h14ad8:	data_out=16'h8fa;
17'h14ad9:	data_out=16'h8889;
17'h14ada:	data_out=16'h870e;
17'h14adb:	data_out=16'h8f;
17'h14adc:	data_out=16'h399;
17'h14add:	data_out=16'h8548;
17'h14ade:	data_out=16'h8711;
17'h14adf:	data_out=16'h88e3;
17'h14ae0:	data_out=16'h8a00;
17'h14ae1:	data_out=16'h9f9;
17'h14ae2:	data_out=16'h89b7;
17'h14ae3:	data_out=16'h86c3;
17'h14ae4:	data_out=16'h89ad;
17'h14ae5:	data_out=16'h8905;
17'h14ae6:	data_out=16'ha00;
17'h14ae7:	data_out=16'ha00;
17'h14ae8:	data_out=16'h9ff;
17'h14ae9:	data_out=16'h8a00;
17'h14aea:	data_out=16'h9ff;
17'h14aeb:	data_out=16'h16d;
17'h14aec:	data_out=16'h9fe;
17'h14aed:	data_out=16'h86d7;
17'h14aee:	data_out=16'h9ff;
17'h14aef:	data_out=16'h8281;
17'h14af0:	data_out=16'h9ff;
17'h14af1:	data_out=16'h94e;
17'h14af2:	data_out=16'h9f9;
17'h14af3:	data_out=16'ha00;
17'h14af4:	data_out=16'h4fc;
17'h14af5:	data_out=16'h9f4;
17'h14af6:	data_out=16'h9f8;
17'h14af7:	data_out=16'h89f4;
17'h14af8:	data_out=16'h89f4;
17'h14af9:	data_out=16'h19d;
17'h14afa:	data_out=16'h8760;
17'h14afb:	data_out=16'h9fe;
17'h14afc:	data_out=16'h9fb;
17'h14afd:	data_out=16'h3c;
17'h14afe:	data_out=16'h89df;
17'h14aff:	data_out=16'h627;
17'h14b00:	data_out=16'h8994;
17'h14b01:	data_out=16'h85cf;
17'h14b02:	data_out=16'h89de;
17'h14b03:	data_out=16'h89df;
17'h14b04:	data_out=16'h29c;
17'h14b05:	data_out=16'h218;
17'h14b06:	data_out=16'h895a;
17'h14b07:	data_out=16'h89fe;
17'h14b08:	data_out=16'h89f6;
17'h14b09:	data_out=16'h89ee;
17'h14b0a:	data_out=16'h9ee;
17'h14b0b:	data_out=16'h89de;
17'h14b0c:	data_out=16'h8a00;
17'h14b0d:	data_out=16'h89e9;
17'h14b0e:	data_out=16'h9ff;
17'h14b0f:	data_out=16'h897b;
17'h14b10:	data_out=16'h89da;
17'h14b11:	data_out=16'h89f7;
17'h14b12:	data_out=16'h8966;
17'h14b13:	data_out=16'h89d1;
17'h14b14:	data_out=16'h88ee;
17'h14b15:	data_out=16'h491;
17'h14b16:	data_out=16'h89b0;
17'h14b17:	data_out=16'h8966;
17'h14b18:	data_out=16'h9fd;
17'h14b19:	data_out=16'h9f9;
17'h14b1a:	data_out=16'h15b;
17'h14b1b:	data_out=16'h89b8;
17'h14b1c:	data_out=16'h89dc;
17'h14b1d:	data_out=16'h89fa;
17'h14b1e:	data_out=16'h8867;
17'h14b1f:	data_out=16'h87e;
17'h14b20:	data_out=16'h86c9;
17'h14b21:	data_out=16'h9ff;
17'h14b22:	data_out=16'h82b0;
17'h14b23:	data_out=16'h8988;
17'h14b24:	data_out=16'h89ae;
17'h14b25:	data_out=16'h89df;
17'h14b26:	data_out=16'h89ff;
17'h14b27:	data_out=16'h89b9;
17'h14b28:	data_out=16'ha00;
17'h14b29:	data_out=16'h8070;
17'h14b2a:	data_out=16'h89cc;
17'h14b2b:	data_out=16'h9ac;
17'h14b2c:	data_out=16'h8940;
17'h14b2d:	data_out=16'h89e2;
17'h14b2e:	data_out=16'h8968;
17'h14b2f:	data_out=16'h8976;
17'h14b30:	data_out=16'h802f;
17'h14b31:	data_out=16'h838d;
17'h14b32:	data_out=16'h89fc;
17'h14b33:	data_out=16'h8789;
17'h14b34:	data_out=16'h88b6;
17'h14b35:	data_out=16'h8588;
17'h14b36:	data_out=16'h89dd;
17'h14b37:	data_out=16'h89de;
17'h14b38:	data_out=16'h897a;
17'h14b39:	data_out=16'h87bc;
17'h14b3a:	data_out=16'h897c;
17'h14b3b:	data_out=16'h89fd;
17'h14b3c:	data_out=16'h81f8;
17'h14b3d:	data_out=16'h84ab;
17'h14b3e:	data_out=16'ha00;
17'h14b3f:	data_out=16'h252;
17'h14b40:	data_out=16'h886d;
17'h14b41:	data_out=16'h89d9;
17'h14b42:	data_out=16'h8a00;
17'h14b43:	data_out=16'h860d;
17'h14b44:	data_out=16'h8192;
17'h14b45:	data_out=16'h37d;
17'h14b46:	data_out=16'h8875;
17'h14b47:	data_out=16'h89ab;
17'h14b48:	data_out=16'h898e;
17'h14b49:	data_out=16'h89e2;
17'h14b4a:	data_out=16'h89c3;
17'h14b4b:	data_out=16'h89ff;
17'h14b4c:	data_out=16'h89eb;
17'h14b4d:	data_out=16'h543;
17'h14b4e:	data_out=16'h89d7;
17'h14b4f:	data_out=16'h89fd;
17'h14b50:	data_out=16'h8912;
17'h14b51:	data_out=16'h9ef;
17'h14b52:	data_out=16'h85f5;
17'h14b53:	data_out=16'h8933;
17'h14b54:	data_out=16'h8847;
17'h14b55:	data_out=16'h470;
17'h14b56:	data_out=16'h8a3;
17'h14b57:	data_out=16'h9ff;
17'h14b58:	data_out=16'h850;
17'h14b59:	data_out=16'h8488;
17'h14b5a:	data_out=16'h8906;
17'h14b5b:	data_out=16'h51;
17'h14b5c:	data_out=16'h88a2;
17'h14b5d:	data_out=16'h88b7;
17'h14b5e:	data_out=16'h899b;
17'h14b5f:	data_out=16'h898e;
17'h14b60:	data_out=16'h8a00;
17'h14b61:	data_out=16'h9ee;
17'h14b62:	data_out=16'h89fa;
17'h14b63:	data_out=16'h87c7;
17'h14b64:	data_out=16'h89f4;
17'h14b65:	data_out=16'h89ec;
17'h14b66:	data_out=16'ha00;
17'h14b67:	data_out=16'ha00;
17'h14b68:	data_out=16'ha00;
17'h14b69:	data_out=16'h89fd;
17'h14b6a:	data_out=16'h9ff;
17'h14b6b:	data_out=16'h8336;
17'h14b6c:	data_out=16'h8884;
17'h14b6d:	data_out=16'h87c1;
17'h14b6e:	data_out=16'h9ff;
17'h14b6f:	data_out=16'h8713;
17'h14b70:	data_out=16'h9ff;
17'h14b71:	data_out=16'h873f;
17'h14b72:	data_out=16'h616;
17'h14b73:	data_out=16'h9f9;
17'h14b74:	data_out=16'h812c;
17'h14b75:	data_out=16'h9d6;
17'h14b76:	data_out=16'ha00;
17'h14b77:	data_out=16'h89f6;
17'h14b78:	data_out=16'h89f6;
17'h14b79:	data_out=16'h849e;
17'h14b7a:	data_out=16'h887c;
17'h14b7b:	data_out=16'ha00;
17'h14b7c:	data_out=16'h9fc;
17'h14b7d:	data_out=16'ha00;
17'h14b7e:	data_out=16'h89ea;
17'h14b7f:	data_out=16'ha00;
17'h14b80:	data_out=16'h8999;
17'h14b81:	data_out=16'h89ff;
17'h14b82:	data_out=16'h89f7;
17'h14b83:	data_out=16'h89f3;
17'h14b84:	data_out=16'h726;
17'h14b85:	data_out=16'h8689;
17'h14b86:	data_out=16'h89fa;
17'h14b87:	data_out=16'h89fd;
17'h14b88:	data_out=16'h89fa;
17'h14b89:	data_out=16'h89f5;
17'h14b8a:	data_out=16'haa;
17'h14b8b:	data_out=16'h89f6;
17'h14b8c:	data_out=16'h89fe;
17'h14b8d:	data_out=16'h89c6;
17'h14b8e:	data_out=16'ha00;
17'h14b8f:	data_out=16'h89f8;
17'h14b90:	data_out=16'h89b6;
17'h14b91:	data_out=16'h89fb;
17'h14b92:	data_out=16'h89d8;
17'h14b93:	data_out=16'h8979;
17'h14b94:	data_out=16'h8994;
17'h14b95:	data_out=16'h954;
17'h14b96:	data_out=16'h89c0;
17'h14b97:	data_out=16'h89f7;
17'h14b98:	data_out=16'ha00;
17'h14b99:	data_out=16'h9f8;
17'h14b9a:	data_out=16'h847a;
17'h14b9b:	data_out=16'h89da;
17'h14b9c:	data_out=16'h8988;
17'h14b9d:	data_out=16'h8a00;
17'h14b9e:	data_out=16'h8991;
17'h14b9f:	data_out=16'h76a;
17'h14ba0:	data_out=16'h8793;
17'h14ba1:	data_out=16'ha00;
17'h14ba2:	data_out=16'ha00;
17'h14ba3:	data_out=16'h8388;
17'h14ba4:	data_out=16'h839e;
17'h14ba5:	data_out=16'h82e7;
17'h14ba6:	data_out=16'h89f9;
17'h14ba7:	data_out=16'h89f5;
17'h14ba8:	data_out=16'ha00;
17'h14ba9:	data_out=16'h85b1;
17'h14baa:	data_out=16'h89fb;
17'h14bab:	data_out=16'h9e3;
17'h14bac:	data_out=16'h8991;
17'h14bad:	data_out=16'h8a00;
17'h14bae:	data_out=16'h89fc;
17'h14baf:	data_out=16'h89f8;
17'h14bb0:	data_out=16'h83a7;
17'h14bb1:	data_out=16'h896a;
17'h14bb2:	data_out=16'h8a00;
17'h14bb3:	data_out=16'h8698;
17'h14bb4:	data_out=16'h8a00;
17'h14bb5:	data_out=16'h874f;
17'h14bb6:	data_out=16'h89f9;
17'h14bb7:	data_out=16'h89f7;
17'h14bb8:	data_out=16'h89fd;
17'h14bb9:	data_out=16'h855e;
17'h14bba:	data_out=16'h8949;
17'h14bbb:	data_out=16'h89fe;
17'h14bbc:	data_out=16'h857a;
17'h14bbd:	data_out=16'h81e3;
17'h14bbe:	data_out=16'ha00;
17'h14bbf:	data_out=16'h8651;
17'h14bc0:	data_out=16'h8778;
17'h14bc1:	data_out=16'h89ef;
17'h14bc2:	data_out=16'h8a00;
17'h14bc3:	data_out=16'h84b9;
17'h14bc4:	data_out=16'h8698;
17'h14bc5:	data_out=16'h873;
17'h14bc6:	data_out=16'h8934;
17'h14bc7:	data_out=16'h89eb;
17'h14bc8:	data_out=16'h89f8;
17'h14bc9:	data_out=16'hb5;
17'h14bca:	data_out=16'h89fc;
17'h14bcb:	data_out=16'h89ff;
17'h14bcc:	data_out=16'h89e9;
17'h14bcd:	data_out=16'ha00;
17'h14bce:	data_out=16'h89fa;
17'h14bcf:	data_out=16'h89fa;
17'h14bd0:	data_out=16'h8265;
17'h14bd1:	data_out=16'h9eb;
17'h14bd2:	data_out=16'h4fa;
17'h14bd3:	data_out=16'h89f8;
17'h14bd4:	data_out=16'h89bc;
17'h14bd5:	data_out=16'h440;
17'h14bd6:	data_out=16'h9ce;
17'h14bd7:	data_out=16'ha00;
17'h14bd8:	data_out=16'h9c6;
17'h14bd9:	data_out=16'h447;
17'h14bda:	data_out=16'h89f8;
17'h14bdb:	data_out=16'h8338;
17'h14bdc:	data_out=16'h89f7;
17'h14bdd:	data_out=16'h89bf;
17'h14bde:	data_out=16'h89fa;
17'h14bdf:	data_out=16'h89ef;
17'h14be0:	data_out=16'h89ff;
17'h14be1:	data_out=16'h82cf;
17'h14be2:	data_out=16'h89f9;
17'h14be3:	data_out=16'h898f;
17'h14be4:	data_out=16'h8a00;
17'h14be5:	data_out=16'h89ff;
17'h14be6:	data_out=16'ha00;
17'h14be7:	data_out=16'ha00;
17'h14be8:	data_out=16'ha00;
17'h14be9:	data_out=16'h89fa;
17'h14bea:	data_out=16'ha00;
17'h14beb:	data_out=16'h857a;
17'h14bec:	data_out=16'h8993;
17'h14bed:	data_out=16'h896f;
17'h14bee:	data_out=16'ha00;
17'h14bef:	data_out=16'h89fb;
17'h14bf0:	data_out=16'ha00;
17'h14bf1:	data_out=16'h89f9;
17'h14bf2:	data_out=16'h43b;
17'h14bf3:	data_out=16'h8279;
17'h14bf4:	data_out=16'h8452;
17'h14bf5:	data_out=16'h9de;
17'h14bf6:	data_out=16'h9fc;
17'h14bf7:	data_out=16'h89f6;
17'h14bf8:	data_out=16'h89fb;
17'h14bf9:	data_out=16'h8668;
17'h14bfa:	data_out=16'h89dd;
17'h14bfb:	data_out=16'ha00;
17'h14bfc:	data_out=16'h8c4;
17'h14bfd:	data_out=16'ha00;
17'h14bfe:	data_out=16'h89ee;
17'h14bff:	data_out=16'ha00;
17'h14c00:	data_out=16'h89b8;
17'h14c01:	data_out=16'h8a00;
17'h14c02:	data_out=16'h8952;
17'h14c03:	data_out=16'h89c5;
17'h14c04:	data_out=16'h213;
17'h14c05:	data_out=16'h8995;
17'h14c06:	data_out=16'h89fe;
17'h14c07:	data_out=16'h89fe;
17'h14c08:	data_out=16'h89f8;
17'h14c09:	data_out=16'h82fc;
17'h14c0a:	data_out=16'h8518;
17'h14c0b:	data_out=16'h89f7;
17'h14c0c:	data_out=16'h8a00;
17'h14c0d:	data_out=16'h88e9;
17'h14c0e:	data_out=16'ha00;
17'h14c0f:	data_out=16'h89fb;
17'h14c10:	data_out=16'h8957;
17'h14c11:	data_out=16'h8a00;
17'h14c12:	data_out=16'h89f9;
17'h14c13:	data_out=16'h88ec;
17'h14c14:	data_out=16'h72e;
17'h14c15:	data_out=16'ha00;
17'h14c16:	data_out=16'h89ce;
17'h14c17:	data_out=16'h89f8;
17'h14c18:	data_out=16'ha00;
17'h14c19:	data_out=16'h85b1;
17'h14c1a:	data_out=16'h8829;
17'h14c1b:	data_out=16'h89a4;
17'h14c1c:	data_out=16'h8345;
17'h14c1d:	data_out=16'h8a00;
17'h14c1e:	data_out=16'h89bc;
17'h14c1f:	data_out=16'h9f2;
17'h14c20:	data_out=16'h8995;
17'h14c21:	data_out=16'ha00;
17'h14c22:	data_out=16'ha00;
17'h14c23:	data_out=16'h9e0;
17'h14c24:	data_out=16'h9f5;
17'h14c25:	data_out=16'h760;
17'h14c26:	data_out=16'h89cd;
17'h14c27:	data_out=16'h89fd;
17'h14c28:	data_out=16'ha00;
17'h14c29:	data_out=16'had;
17'h14c2a:	data_out=16'h89fe;
17'h14c2b:	data_out=16'h9ce;
17'h14c2c:	data_out=16'h87ec;
17'h14c2d:	data_out=16'h8a00;
17'h14c2e:	data_out=16'h89ff;
17'h14c2f:	data_out=16'h89fe;
17'h14c30:	data_out=16'h87e6;
17'h14c31:	data_out=16'h8a00;
17'h14c32:	data_out=16'h8a00;
17'h14c33:	data_out=16'h724;
17'h14c34:	data_out=16'h8a00;
17'h14c35:	data_out=16'h892c;
17'h14c36:	data_out=16'h89fa;
17'h14c37:	data_out=16'h89f3;
17'h14c38:	data_out=16'h8a00;
17'h14c39:	data_out=16'h935;
17'h14c3a:	data_out=16'h89ab;
17'h14c3b:	data_out=16'h89fc;
17'h14c3c:	data_out=16'h86ed;
17'h14c3d:	data_out=16'h93f;
17'h14c3e:	data_out=16'ha00;
17'h14c3f:	data_out=16'h8969;
17'h14c40:	data_out=16'h89e0;
17'h14c41:	data_out=16'h89e6;
17'h14c42:	data_out=16'h89ff;
17'h14c43:	data_out=16'h8114;
17'h14c44:	data_out=16'h886e;
17'h14c45:	data_out=16'ha00;
17'h14c46:	data_out=16'h88e8;
17'h14c47:	data_out=16'h89fc;
17'h14c48:	data_out=16'h89fe;
17'h14c49:	data_out=16'ha00;
17'h14c4a:	data_out=16'h8a00;
17'h14c4b:	data_out=16'h8a00;
17'h14c4c:	data_out=16'h89d9;
17'h14c4d:	data_out=16'ha00;
17'h14c4e:	data_out=16'h89fb;
17'h14c4f:	data_out=16'h89ed;
17'h14c50:	data_out=16'h516;
17'h14c51:	data_out=16'ha00;
17'h14c52:	data_out=16'h9dc;
17'h14c53:	data_out=16'h89ff;
17'h14c54:	data_out=16'h89fd;
17'h14c55:	data_out=16'h89f;
17'h14c56:	data_out=16'ha00;
17'h14c57:	data_out=16'ha00;
17'h14c58:	data_out=16'ha00;
17'h14c59:	data_out=16'h6cc;
17'h14c5a:	data_out=16'h89ef;
17'h14c5b:	data_out=16'h82b2;
17'h14c5c:	data_out=16'h89f8;
17'h14c5d:	data_out=16'h89ff;
17'h14c5e:	data_out=16'h89fe;
17'h14c5f:	data_out=16'h8a00;
17'h14c60:	data_out=16'h89fc;
17'h14c61:	data_out=16'h86f5;
17'h14c62:	data_out=16'h89fa;
17'h14c63:	data_out=16'h126;
17'h14c64:	data_out=16'h8a00;
17'h14c65:	data_out=16'h8a00;
17'h14c66:	data_out=16'h8239;
17'h14c67:	data_out=16'h838d;
17'h14c68:	data_out=16'ha00;
17'h14c69:	data_out=16'h89f5;
17'h14c6a:	data_out=16'ha00;
17'h14c6b:	data_out=16'h87f7;
17'h14c6c:	data_out=16'h89e4;
17'h14c6d:	data_out=16'h22f;
17'h14c6e:	data_out=16'ha00;
17'h14c6f:	data_out=16'h89ff;
17'h14c70:	data_out=16'ha00;
17'h14c71:	data_out=16'h89fd;
17'h14c72:	data_out=16'h7ac;
17'h14c73:	data_out=16'h86ab;
17'h14c74:	data_out=16'h8868;
17'h14c75:	data_out=16'h9fa;
17'h14c76:	data_out=16'h9f8;
17'h14c77:	data_out=16'h8290;
17'h14c78:	data_out=16'h8917;
17'h14c79:	data_out=16'h8599;
17'h14c7a:	data_out=16'h81a8;
17'h14c7b:	data_out=16'ha00;
17'h14c7c:	data_out=16'h7f6;
17'h14c7d:	data_out=16'ha00;
17'h14c7e:	data_out=16'h89cc;
17'h14c7f:	data_out=16'ha00;
17'h14c80:	data_out=16'h89cd;
17'h14c81:	data_out=16'h8a00;
17'h14c82:	data_out=16'h89fb;
17'h14c83:	data_out=16'h898b;
17'h14c84:	data_out=16'h80de;
17'h14c85:	data_out=16'h89f2;
17'h14c86:	data_out=16'h857c;
17'h14c87:	data_out=16'h89ff;
17'h14c88:	data_out=16'h89fd;
17'h14c89:	data_out=16'h502;
17'h14c8a:	data_out=16'h85ea;
17'h14c8b:	data_out=16'h89d0;
17'h14c8c:	data_out=16'h89ff;
17'h14c8d:	data_out=16'h89d4;
17'h14c8e:	data_out=16'ha00;
17'h14c8f:	data_out=16'h89fe;
17'h14c90:	data_out=16'h59b;
17'h14c91:	data_out=16'h8955;
17'h14c92:	data_out=16'h89fd;
17'h14c93:	data_out=16'h8857;
17'h14c94:	data_out=16'h999;
17'h14c95:	data_out=16'h9ff;
17'h14c96:	data_out=16'h89e4;
17'h14c97:	data_out=16'h89fa;
17'h14c98:	data_out=16'h9e6;
17'h14c99:	data_out=16'h4b4;
17'h14c9a:	data_out=16'h8993;
17'h14c9b:	data_out=16'h8973;
17'h14c9c:	data_out=16'h30f;
17'h14c9d:	data_out=16'h8a00;
17'h14c9e:	data_out=16'h881e;
17'h14c9f:	data_out=16'h99f;
17'h14ca0:	data_out=16'h89ca;
17'h14ca1:	data_out=16'ha00;
17'h14ca2:	data_out=16'ha00;
17'h14ca3:	data_out=16'h339;
17'h14ca4:	data_out=16'h349;
17'h14ca5:	data_out=16'ha00;
17'h14ca6:	data_out=16'h86ac;
17'h14ca7:	data_out=16'h89fe;
17'h14ca8:	data_out=16'ha00;
17'h14ca9:	data_out=16'h5f;
17'h14caa:	data_out=16'h89ff;
17'h14cab:	data_out=16'h9f4;
17'h14cac:	data_out=16'h89cf;
17'h14cad:	data_out=16'h8a00;
17'h14cae:	data_out=16'h8a00;
17'h14caf:	data_out=16'h8a00;
17'h14cb0:	data_out=16'h890c;
17'h14cb1:	data_out=16'h89fc;
17'h14cb2:	data_out=16'h8a00;
17'h14cb3:	data_out=16'h98d;
17'h14cb4:	data_out=16'h8a00;
17'h14cb5:	data_out=16'h8891;
17'h14cb6:	data_out=16'h89fe;
17'h14cb7:	data_out=16'h89fb;
17'h14cb8:	data_out=16'h8a00;
17'h14cb9:	data_out=16'h9fd;
17'h14cba:	data_out=16'h865a;
17'h14cbb:	data_out=16'h89ff;
17'h14cbc:	data_out=16'h864a;
17'h14cbd:	data_out=16'h9ee;
17'h14cbe:	data_out=16'ha00;
17'h14cbf:	data_out=16'h89f1;
17'h14cc0:	data_out=16'h8322;
17'h14cc1:	data_out=16'h89b8;
17'h14cc2:	data_out=16'h89fd;
17'h14cc3:	data_out=16'h973;
17'h14cc4:	data_out=16'h8948;
17'h14cc5:	data_out=16'h9fe;
17'h14cc6:	data_out=16'h8173;
17'h14cc7:	data_out=16'h89fe;
17'h14cc8:	data_out=16'h8a00;
17'h14cc9:	data_out=16'ha00;
17'h14cca:	data_out=16'h8a00;
17'h14ccb:	data_out=16'h89fe;
17'h14ccc:	data_out=16'h89e5;
17'h14ccd:	data_out=16'ha00;
17'h14cce:	data_out=16'h89fc;
17'h14ccf:	data_out=16'h8783;
17'h14cd0:	data_out=16'h8de;
17'h14cd1:	data_out=16'ha00;
17'h14cd2:	data_out=16'h9fa;
17'h14cd3:	data_out=16'h8a00;
17'h14cd4:	data_out=16'h8a00;
17'h14cd5:	data_out=16'h98b;
17'h14cd6:	data_out=16'ha00;
17'h14cd7:	data_out=16'ha00;
17'h14cd8:	data_out=16'ha00;
17'h14cd9:	data_out=16'h9d8;
17'h14cda:	data_out=16'h89f2;
17'h14cdb:	data_out=16'h7c1;
17'h14cdc:	data_out=16'h89ff;
17'h14cdd:	data_out=16'h8a00;
17'h14cde:	data_out=16'h8a00;
17'h14cdf:	data_out=16'h8a00;
17'h14ce0:	data_out=16'h89d8;
17'h14ce1:	data_out=16'h8794;
17'h14ce2:	data_out=16'h89fa;
17'h14ce3:	data_out=16'h64b;
17'h14ce4:	data_out=16'h89fa;
17'h14ce5:	data_out=16'h8a00;
17'h14ce6:	data_out=16'h803;
17'h14ce7:	data_out=16'hdf;
17'h14ce8:	data_out=16'ha00;
17'h14ce9:	data_out=16'h89f7;
17'h14cea:	data_out=16'ha00;
17'h14ceb:	data_out=16'h86e6;
17'h14cec:	data_out=16'h89f4;
17'h14ced:	data_out=16'h6d6;
17'h14cee:	data_out=16'ha00;
17'h14cef:	data_out=16'h8a00;
17'h14cf0:	data_out=16'ha00;
17'h14cf1:	data_out=16'h89ff;
17'h14cf2:	data_out=16'h559;
17'h14cf3:	data_out=16'h86ed;
17'h14cf4:	data_out=16'h8939;
17'h14cf5:	data_out=16'h974;
17'h14cf6:	data_out=16'ha00;
17'h14cf7:	data_out=16'h4e1;
17'h14cf8:	data_out=16'h14d;
17'h14cf9:	data_out=16'h87d2;
17'h14cfa:	data_out=16'h64a;
17'h14cfb:	data_out=16'ha00;
17'h14cfc:	data_out=16'h8014;
17'h14cfd:	data_out=16'h9ff;
17'h14cfe:	data_out=16'h881;
17'h14cff:	data_out=16'h9ff;
17'h14d00:	data_out=16'h4aa;
17'h14d01:	data_out=16'h8a00;
17'h14d02:	data_out=16'h89fd;
17'h14d03:	data_out=16'h8292;
17'h14d04:	data_out=16'h8376;
17'h14d05:	data_out=16'h89f9;
17'h14d06:	data_out=16'h80c6;
17'h14d07:	data_out=16'h8a00;
17'h14d08:	data_out=16'h89ef;
17'h14d09:	data_out=16'h7c0;
17'h14d0a:	data_out=16'h8924;
17'h14d0b:	data_out=16'h8560;
17'h14d0c:	data_out=16'h89ff;
17'h14d0d:	data_out=16'h89f9;
17'h14d0e:	data_out=16'h5b7;
17'h14d0f:	data_out=16'h8a00;
17'h14d10:	data_out=16'h9fc;
17'h14d11:	data_out=16'h88cf;
17'h14d12:	data_out=16'h8a00;
17'h14d13:	data_out=16'h88a2;
17'h14d14:	data_out=16'h9fa;
17'h14d15:	data_out=16'ha00;
17'h14d16:	data_out=16'h89ef;
17'h14d17:	data_out=16'h86e9;
17'h14d18:	data_out=16'h7fd;
17'h14d19:	data_out=16'h93;
17'h14d1a:	data_out=16'h89d5;
17'h14d1b:	data_out=16'h8983;
17'h14d1c:	data_out=16'h51f;
17'h14d1d:	data_out=16'h8a00;
17'h14d1e:	data_out=16'h86d3;
17'h14d1f:	data_out=16'h6b9;
17'h14d20:	data_out=16'h88d;
17'h14d21:	data_out=16'h586;
17'h14d22:	data_out=16'ha00;
17'h14d23:	data_out=16'h6f3;
17'h14d24:	data_out=16'h6ff;
17'h14d25:	data_out=16'ha00;
17'h14d26:	data_out=16'ha00;
17'h14d27:	data_out=16'h89cd;
17'h14d28:	data_out=16'h569;
17'h14d29:	data_out=16'h8183;
17'h14d2a:	data_out=16'h89ff;
17'h14d2b:	data_out=16'h9fd;
17'h14d2c:	data_out=16'h849c;
17'h14d2d:	data_out=16'h8987;
17'h14d2e:	data_out=16'h8a00;
17'h14d2f:	data_out=16'h89ff;
17'h14d30:	data_out=16'h89ab;
17'h14d31:	data_out=16'h89f0;
17'h14d32:	data_out=16'h89ff;
17'h14d33:	data_out=16'h9f7;
17'h14d34:	data_out=16'h8a00;
17'h14d35:	data_out=16'h8810;
17'h14d36:	data_out=16'h89fb;
17'h14d37:	data_out=16'h89fe;
17'h14d38:	data_out=16'h82f8;
17'h14d39:	data_out=16'h9fb;
17'h14d3a:	data_out=16'h8145;
17'h14d3b:	data_out=16'h89fe;
17'h14d3c:	data_out=16'h85fb;
17'h14d3d:	data_out=16'h9fa;
17'h14d3e:	data_out=16'h567;
17'h14d3f:	data_out=16'h89f7;
17'h14d40:	data_out=16'h5a8;
17'h14d41:	data_out=16'h8955;
17'h14d42:	data_out=16'h89fd;
17'h14d43:	data_out=16'h944;
17'h14d44:	data_out=16'h2a4;
17'h14d45:	data_out=16'h9ff;
17'h14d46:	data_out=16'ha00;
17'h14d47:	data_out=16'h885a;
17'h14d48:	data_out=16'h8a00;
17'h14d49:	data_out=16'ha00;
17'h14d4a:	data_out=16'h8a00;
17'h14d4b:	data_out=16'h89fe;
17'h14d4c:	data_out=16'h89f7;
17'h14d4d:	data_out=16'ha00;
17'h14d4e:	data_out=16'h89fc;
17'h14d4f:	data_out=16'h8542;
17'h14d50:	data_out=16'h9a8;
17'h14d51:	data_out=16'h9ea;
17'h14d52:	data_out=16'ha00;
17'h14d53:	data_out=16'h8a00;
17'h14d54:	data_out=16'h89e4;
17'h14d55:	data_out=16'h917;
17'h14d56:	data_out=16'ha00;
17'h14d57:	data_out=16'ha00;
17'h14d58:	data_out=16'ha00;
17'h14d59:	data_out=16'h9f6;
17'h14d5a:	data_out=16'h89f9;
17'h14d5b:	data_out=16'h4cc;
17'h14d5c:	data_out=16'h89fb;
17'h14d5d:	data_out=16'h89f7;
17'h14d5e:	data_out=16'h89ff;
17'h14d5f:	data_out=16'h8a00;
17'h14d60:	data_out=16'h89dc;
17'h14d61:	data_out=16'h80ee;
17'h14d62:	data_out=16'h89fa;
17'h14d63:	data_out=16'h8a4;
17'h14d64:	data_out=16'h2d9;
17'h14d65:	data_out=16'h8a00;
17'h14d66:	data_out=16'h23f;
17'h14d67:	data_out=16'hcd;
17'h14d68:	data_out=16'h581;
17'h14d69:	data_out=16'h89f4;
17'h14d6a:	data_out=16'h5ea;
17'h14d6b:	data_out=16'h8342;
17'h14d6c:	data_out=16'h89d3;
17'h14d6d:	data_out=16'h900;
17'h14d6e:	data_out=16'h5e8;
17'h14d6f:	data_out=16'h8a00;
17'h14d70:	data_out=16'h5ca;
17'h14d71:	data_out=16'h8a00;
17'h14d72:	data_out=16'h84c6;
17'h14d73:	data_out=16'h31d;
17'h14d74:	data_out=16'h89b3;
17'h14d75:	data_out=16'h8958;
17'h14d76:	data_out=16'ha00;
17'h14d77:	data_out=16'h876;
17'h14d78:	data_out=16'h282;
17'h14d79:	data_out=16'h8858;
17'h14d7a:	data_out=16'h8be;
17'h14d7b:	data_out=16'h563;
17'h14d7c:	data_out=16'h8358;
17'h14d7d:	data_out=16'h2ec;
17'h14d7e:	data_out=16'h9a9;
17'h14d7f:	data_out=16'h9ff;
17'h14d80:	data_out=16'h9fd;
17'h14d81:	data_out=16'h89fd;
17'h14d82:	data_out=16'h8597;
17'h14d83:	data_out=16'h19c;
17'h14d84:	data_out=16'h82dd;
17'h14d85:	data_out=16'h8805;
17'h14d86:	data_out=16'h97;
17'h14d87:	data_out=16'h8a00;
17'h14d88:	data_out=16'h607;
17'h14d89:	data_out=16'h951;
17'h14d8a:	data_out=16'h895b;
17'h14d8b:	data_out=16'h819;
17'h14d8c:	data_out=16'h8a00;
17'h14d8d:	data_out=16'h89de;
17'h14d8e:	data_out=16'h2c1;
17'h14d8f:	data_out=16'h8a00;
17'h14d90:	data_out=16'ha00;
17'h14d91:	data_out=16'h8863;
17'h14d92:	data_out=16'h8a00;
17'h14d93:	data_out=16'h854d;
17'h14d94:	data_out=16'h838;
17'h14d95:	data_out=16'h9ff;
17'h14d96:	data_out=16'h843a;
17'h14d97:	data_out=16'h8301;
17'h14d98:	data_out=16'h3f9;
17'h14d99:	data_out=16'h8036;
17'h14d9a:	data_out=16'h89e3;
17'h14d9b:	data_out=16'h8844;
17'h14d9c:	data_out=16'h578;
17'h14d9d:	data_out=16'h8a00;
17'h14d9e:	data_out=16'h8449;
17'h14d9f:	data_out=16'h702;
17'h14da0:	data_out=16'h7e3;
17'h14da1:	data_out=16'h2ab;
17'h14da2:	data_out=16'ha00;
17'h14da3:	data_out=16'h8043;
17'h14da4:	data_out=16'h8039;
17'h14da5:	data_out=16'h951;
17'h14da6:	data_out=16'ha00;
17'h14da7:	data_out=16'h89c2;
17'h14da8:	data_out=16'h2ad;
17'h14da9:	data_out=16'h420;
17'h14daa:	data_out=16'h8a00;
17'h14dab:	data_out=16'ha00;
17'h14dac:	data_out=16'h103;
17'h14dad:	data_out=16'h5a3;
17'h14dae:	data_out=16'h8a00;
17'h14daf:	data_out=16'h8a00;
17'h14db0:	data_out=16'h8996;
17'h14db1:	data_out=16'h89fa;
17'h14db2:	data_out=16'h89fa;
17'h14db3:	data_out=16'h9ee;
17'h14db4:	data_out=16'h8a00;
17'h14db5:	data_out=16'h86a3;
17'h14db6:	data_out=16'h8570;
17'h14db7:	data_out=16'h8637;
17'h14db8:	data_out=16'h831b;
17'h14db9:	data_out=16'h7a0;
17'h14dba:	data_out=16'h34a;
17'h14dbb:	data_out=16'h852f;
17'h14dbc:	data_out=16'h85ba;
17'h14dbd:	data_out=16'h9fb;
17'h14dbe:	data_out=16'h2ac;
17'h14dbf:	data_out=16'h87c4;
17'h14dc0:	data_out=16'h860;
17'h14dc1:	data_out=16'h4e3;
17'h14dc2:	data_out=16'h89ed;
17'h14dc3:	data_out=16'h6ba;
17'h14dc4:	data_out=16'h54c;
17'h14dc5:	data_out=16'h9f6;
17'h14dc6:	data_out=16'ha00;
17'h14dc7:	data_out=16'h8339;
17'h14dc8:	data_out=16'h8a00;
17'h14dc9:	data_out=16'ha00;
17'h14dca:	data_out=16'h8a00;
17'h14dcb:	data_out=16'h89ff;
17'h14dcc:	data_out=16'h89db;
17'h14dcd:	data_out=16'ha00;
17'h14dce:	data_out=16'h89fd;
17'h14dcf:	data_out=16'h852b;
17'h14dd0:	data_out=16'h9c3;
17'h14dd1:	data_out=16'h9fb;
17'h14dd2:	data_out=16'h359;
17'h14dd3:	data_out=16'h8a00;
17'h14dd4:	data_out=16'h8093;
17'h14dd5:	data_out=16'h9b7;
17'h14dd6:	data_out=16'ha00;
17'h14dd7:	data_out=16'ha00;
17'h14dd8:	data_out=16'ha00;
17'h14dd9:	data_out=16'h9f9;
17'h14dda:	data_out=16'h89f9;
17'h14ddb:	data_out=16'h243;
17'h14ddc:	data_out=16'h89f9;
17'h14ddd:	data_out=16'h89f5;
17'h14dde:	data_out=16'h8a00;
17'h14ddf:	data_out=16'h8809;
17'h14de0:	data_out=16'h4b8;
17'h14de1:	data_out=16'hd0;
17'h14de2:	data_out=16'h89f1;
17'h14de3:	data_out=16'h893;
17'h14de4:	data_out=16'h61f;
17'h14de5:	data_out=16'h89ff;
17'h14de6:	data_out=16'h810e;
17'h14de7:	data_out=16'h60;
17'h14de8:	data_out=16'h2ae;
17'h14de9:	data_out=16'h3f6;
17'h14dea:	data_out=16'h2da;
17'h14deb:	data_out=16'h8087;
17'h14dec:	data_out=16'h8973;
17'h14ded:	data_out=16'h8c0;
17'h14dee:	data_out=16'h2d9;
17'h14def:	data_out=16'h8a00;
17'h14df0:	data_out=16'h2cb;
17'h14df1:	data_out=16'h8a00;
17'h14df2:	data_out=16'h859b;
17'h14df3:	data_out=16'h1d3;
17'h14df4:	data_out=16'h8985;
17'h14df5:	data_out=16'h89c4;
17'h14df6:	data_out=16'ha00;
17'h14df7:	data_out=16'h9d2;
17'h14df8:	data_out=16'ha5;
17'h14df9:	data_out=16'h88ef;
17'h14dfa:	data_out=16'h789;
17'h14dfb:	data_out=16'h2aa;
17'h14dfc:	data_out=16'h8321;
17'h14dfd:	data_out=16'h82bd;
17'h14dfe:	data_out=16'ha00;
17'h14dff:	data_out=16'h9ff;
17'h14e00:	data_out=16'h930;
17'h14e01:	data_out=16'h8a00;
17'h14e02:	data_out=16'h801f;
17'h14e03:	data_out=16'h80eb;
17'h14e04:	data_out=16'h84cb;
17'h14e05:	data_out=16'h8850;
17'h14e06:	data_out=16'h8504;
17'h14e07:	data_out=16'h867c;
17'h14e08:	data_out=16'h804;
17'h14e09:	data_out=16'h9cb;
17'h14e0a:	data_out=16'h8a00;
17'h14e0b:	data_out=16'h5ef;
17'h14e0c:	data_out=16'h8a00;
17'h14e0d:	data_out=16'h85d7;
17'h14e0e:	data_out=16'h76;
17'h14e0f:	data_out=16'h84ec;
17'h14e10:	data_out=16'ha00;
17'h14e11:	data_out=16'h88fb;
17'h14e12:	data_out=16'h8a00;
17'h14e13:	data_out=16'h82f2;
17'h14e14:	data_out=16'h4a1;
17'h14e15:	data_out=16'h3d8;
17'h14e16:	data_out=16'h8230;
17'h14e17:	data_out=16'h8091;
17'h14e18:	data_out=16'h3ac;
17'h14e19:	data_out=16'h8407;
17'h14e1a:	data_out=16'h8942;
17'h14e1b:	data_out=16'h8833;
17'h14e1c:	data_out=16'h81a7;
17'h14e1d:	data_out=16'h8894;
17'h14e1e:	data_out=16'h813b;
17'h14e1f:	data_out=16'h400;
17'h14e20:	data_out=16'h577;
17'h14e21:	data_out=16'h75;
17'h14e22:	data_out=16'ha00;
17'h14e23:	data_out=16'h8327;
17'h14e24:	data_out=16'h8321;
17'h14e25:	data_out=16'h3af;
17'h14e26:	data_out=16'h9fa;
17'h14e27:	data_out=16'h85ff;
17'h14e28:	data_out=16'h81;
17'h14e29:	data_out=16'h4c8;
17'h14e2a:	data_out=16'h8936;
17'h14e2b:	data_out=16'h6d4;
17'h14e2c:	data_out=16'h80ed;
17'h14e2d:	data_out=16'h829f;
17'h14e2e:	data_out=16'h8317;
17'h14e2f:	data_out=16'h83d9;
17'h14e30:	data_out=16'h89fe;
17'h14e31:	data_out=16'h8a00;
17'h14e32:	data_out=16'h8a00;
17'h14e33:	data_out=16'h63b;
17'h14e34:	data_out=16'h88b6;
17'h14e35:	data_out=16'h8775;
17'h14e36:	data_out=16'h3e9;
17'h14e37:	data_out=16'h81a7;
17'h14e38:	data_out=16'h8904;
17'h14e39:	data_out=16'h580;
17'h14e3a:	data_out=16'h36;
17'h14e3b:	data_out=16'h8452;
17'h14e3c:	data_out=16'h8144;
17'h14e3d:	data_out=16'h9ff;
17'h14e3e:	data_out=16'h81;
17'h14e3f:	data_out=16'h8832;
17'h14e40:	data_out=16'h8122;
17'h14e41:	data_out=16'h819;
17'h14e42:	data_out=16'h8a00;
17'h14e43:	data_out=16'h80ae;
17'h14e44:	data_out=16'h5e;
17'h14e45:	data_out=16'h446;
17'h14e46:	data_out=16'h6da;
17'h14e47:	data_out=16'h82e3;
17'h14e48:	data_out=16'h879e;
17'h14e49:	data_out=16'h496;
17'h14e4a:	data_out=16'h8a00;
17'h14e4b:	data_out=16'h8a00;
17'h14e4c:	data_out=16'h88fd;
17'h14e4d:	data_out=16'ha00;
17'h14e4e:	data_out=16'h89fc;
17'h14e4f:	data_out=16'h8764;
17'h14e50:	data_out=16'h6a8;
17'h14e51:	data_out=16'h4ba;
17'h14e52:	data_out=16'h82c3;
17'h14e53:	data_out=16'h8a00;
17'h14e54:	data_out=16'h206;
17'h14e55:	data_out=16'h9ae;
17'h14e56:	data_out=16'h795;
17'h14e57:	data_out=16'h83e;
17'h14e58:	data_out=16'ha00;
17'h14e59:	data_out=16'h81cd;
17'h14e5a:	data_out=16'h87e2;
17'h14e5b:	data_out=16'h8349;
17'h14e5c:	data_out=16'h895c;
17'h14e5d:	data_out=16'h8974;
17'h14e5e:	data_out=16'h843e;
17'h14e5f:	data_out=16'h81a7;
17'h14e60:	data_out=16'h8307;
17'h14e61:	data_out=16'h83b7;
17'h14e62:	data_out=16'h857f;
17'h14e63:	data_out=16'h598;
17'h14e64:	data_out=16'h80c5;
17'h14e65:	data_out=16'h8a00;
17'h14e66:	data_out=16'h8337;
17'h14e67:	data_out=16'h8071;
17'h14e68:	data_out=16'h7b;
17'h14e69:	data_out=16'h58f;
17'h14e6a:	data_out=16'h7c;
17'h14e6b:	data_out=16'h8442;
17'h14e6c:	data_out=16'h89bf;
17'h14e6d:	data_out=16'h59a;
17'h14e6e:	data_out=16'h7c;
17'h14e6f:	data_out=16'h8a00;
17'h14e70:	data_out=16'h78;
17'h14e71:	data_out=16'h8a00;
17'h14e72:	data_out=16'h89fc;
17'h14e73:	data_out=16'h8753;
17'h14e74:	data_out=16'h89fd;
17'h14e75:	data_out=16'h89fe;
17'h14e76:	data_out=16'h3b9;
17'h14e77:	data_out=16'h9e6;
17'h14e78:	data_out=16'h852a;
17'h14e79:	data_out=16'h8624;
17'h14e7a:	data_out=16'h4c3;
17'h14e7b:	data_out=16'h80;
17'h14e7c:	data_out=16'hd5;
17'h14e7d:	data_out=16'h8573;
17'h14e7e:	data_out=16'ha00;
17'h14e7f:	data_out=16'h189;
17'h14e80:	data_out=16'h944;
17'h14e81:	data_out=16'h55;
17'h14e82:	data_out=16'h836b;
17'h14e83:	data_out=16'h8241;
17'h14e84:	data_out=16'h36d;
17'h14e85:	data_out=16'ha2;
17'h14e86:	data_out=16'h842e;
17'h14e87:	data_out=16'h8021;
17'h14e88:	data_out=16'h211;
17'h14e89:	data_out=16'h556;
17'h14e8a:	data_out=16'h8002;
17'h14e8b:	data_out=16'h8831;
17'h14e8c:	data_out=16'h8568;
17'h14e8d:	data_out=16'h82ab;
17'h14e8e:	data_out=16'h80c8;
17'h14e8f:	data_out=16'h829f;
17'h14e90:	data_out=16'h29e;
17'h14e91:	data_out=16'h2b3;
17'h14e92:	data_out=16'h883f;
17'h14e93:	data_out=16'h83be;
17'h14e94:	data_out=16'h8308;
17'h14e95:	data_out=16'h388;
17'h14e96:	data_out=16'h146;
17'h14e97:	data_out=16'h8651;
17'h14e98:	data_out=16'h141;
17'h14e99:	data_out=16'he7;
17'h14e9a:	data_out=16'h181;
17'h14e9b:	data_out=16'h86fa;
17'h14e9c:	data_out=16'h171;
17'h14e9d:	data_out=16'h87;
17'h14e9e:	data_out=16'h831c;
17'h14e9f:	data_out=16'h14a;
17'h14ea0:	data_out=16'h6d1;
17'h14ea1:	data_out=16'h80c4;
17'h14ea2:	data_out=16'h34a;
17'h14ea3:	data_out=16'h80ca;
17'h14ea4:	data_out=16'h80c7;
17'h14ea5:	data_out=16'h92;
17'h14ea6:	data_out=16'h80f7;
17'h14ea7:	data_out=16'h152;
17'h14ea8:	data_out=16'h80c1;
17'h14ea9:	data_out=16'h81b0;
17'h14eaa:	data_out=16'h8761;
17'h14eab:	data_out=16'h21f;
17'h14eac:	data_out=16'h1df;
17'h14ead:	data_out=16'h8494;
17'h14eae:	data_out=16'h8527;
17'h14eaf:	data_out=16'h809b;
17'h14eb0:	data_out=16'h8550;
17'h14eb1:	data_out=16'h25;
17'h14eb2:	data_out=16'h8585;
17'h14eb3:	data_out=16'h811f;
17'h14eb4:	data_out=16'h10c;
17'h14eb5:	data_out=16'h28;
17'h14eb6:	data_out=16'h3;
17'h14eb7:	data_out=16'h8411;
17'h14eb8:	data_out=16'h392;
17'h14eb9:	data_out=16'h8078;
17'h14eba:	data_out=16'hfd;
17'h14ebb:	data_out=16'h380;
17'h14ebc:	data_out=16'h867c;
17'h14ebd:	data_out=16'h9bf;
17'h14ebe:	data_out=16'h80c4;
17'h14ebf:	data_out=16'h106;
17'h14ec0:	data_out=16'h159;
17'h14ec1:	data_out=16'h81da;
17'h14ec2:	data_out=16'h88c7;
17'h14ec3:	data_out=16'h828d;
17'h14ec4:	data_out=16'h3ce;
17'h14ec5:	data_out=16'h37d;
17'h14ec6:	data_out=16'h81e0;
17'h14ec7:	data_out=16'h8121;
17'h14ec8:	data_out=16'h8494;
17'h14ec9:	data_out=16'h140;
17'h14eca:	data_out=16'h813a;
17'h14ecb:	data_out=16'h8a00;
17'h14ecc:	data_out=16'h839e;
17'h14ecd:	data_out=16'h3b7;
17'h14ece:	data_out=16'h85fe;
17'h14ecf:	data_out=16'h8227;
17'h14ed0:	data_out=16'h1cd;
17'h14ed1:	data_out=16'h51;
17'h14ed2:	data_out=16'h805a;
17'h14ed3:	data_out=16'h8439;
17'h14ed4:	data_out=16'h2c8;
17'h14ed5:	data_out=16'h8269;
17'h14ed6:	data_out=16'h50;
17'h14ed7:	data_out=16'h117;
17'h14ed8:	data_out=16'h816f;
17'h14ed9:	data_out=16'h191;
17'h14eda:	data_out=16'h8a00;
17'h14edb:	data_out=16'h37f;
17'h14edc:	data_out=16'h2a;
17'h14edd:	data_out=16'h8291;
17'h14ede:	data_out=16'h8142;
17'h14edf:	data_out=16'h77;
17'h14ee0:	data_out=16'h8410;
17'h14ee1:	data_out=16'h4a5;
17'h14ee2:	data_out=16'h88e5;
17'h14ee3:	data_out=16'h817d;
17'h14ee4:	data_out=16'h355;
17'h14ee5:	data_out=16'h8111;
17'h14ee6:	data_out=16'h144;
17'h14ee7:	data_out=16'h8379;
17'h14ee8:	data_out=16'h80c2;
17'h14ee9:	data_out=16'h8097;
17'h14eea:	data_out=16'h80cb;
17'h14eeb:	data_out=16'h518;
17'h14eec:	data_out=16'h828b;
17'h14eed:	data_out=16'h815e;
17'h14eee:	data_out=16'h80d6;
17'h14eef:	data_out=16'h84de;
17'h14ef0:	data_out=16'h80c4;
17'h14ef1:	data_out=16'h82eb;
17'h14ef2:	data_out=16'h8050;
17'h14ef3:	data_out=16'h19f;
17'h14ef4:	data_out=16'h8566;
17'h14ef5:	data_out=16'h8863;
17'h14ef6:	data_out=16'h19d;
17'h14ef7:	data_out=16'h193;
17'h14ef8:	data_out=16'h820c;
17'h14ef9:	data_out=16'h8523;
17'h14efa:	data_out=16'h8267;
17'h14efb:	data_out=16'h80c0;
17'h14efc:	data_out=16'h76;
17'h14efd:	data_out=16'h82f9;
17'h14efe:	data_out=16'h45b;
17'h14eff:	data_out=16'h39f;
17'h14f00:	data_out=16'h8d;
17'h14f01:	data_out=16'hdd;
17'h14f02:	data_out=16'h804a;
17'h14f03:	data_out=16'h66;
17'h14f04:	data_out=16'h91;
17'h14f05:	data_out=16'hbf;
17'h14f06:	data_out=16'h39;
17'h14f07:	data_out=16'hde;
17'h14f08:	data_out=16'h61;
17'h14f09:	data_out=16'h10;
17'h14f0a:	data_out=16'h8021;
17'h14f0b:	data_out=16'h8044;
17'h14f0c:	data_out=16'h8026;
17'h14f0d:	data_out=16'h103;
17'h14f0e:	data_out=16'h801e;
17'h14f0f:	data_out=16'h9c;
17'h14f10:	data_out=16'h8043;
17'h14f11:	data_out=16'h1b;
17'h14f12:	data_out=16'h8099;
17'h14f13:	data_out=16'h66;
17'h14f14:	data_out=16'haa;
17'h14f15:	data_out=16'hd5;
17'h14f16:	data_out=16'h14c;
17'h14f17:	data_out=16'h5f;
17'h14f18:	data_out=16'h21;
17'h14f19:	data_out=16'h80e5;
17'h14f1a:	data_out=16'h51;
17'h14f1b:	data_out=16'h8038;
17'h14f1c:	data_out=16'hac;
17'h14f1d:	data_out=16'h16;
17'h14f1e:	data_out=16'h32;
17'h14f1f:	data_out=16'he4;
17'h14f20:	data_out=16'h159;
17'h14f21:	data_out=16'h8018;
17'h14f22:	data_out=16'h8072;
17'h14f23:	data_out=16'h8073;
17'h14f24:	data_out=16'h8074;
17'h14f25:	data_out=16'h8025;
17'h14f26:	data_out=16'h8084;
17'h14f27:	data_out=16'h3b;
17'h14f28:	data_out=16'h801a;
17'h14f29:	data_out=16'h3;
17'h14f2a:	data_out=16'h809a;
17'h14f2b:	data_out=16'h8043;
17'h14f2c:	data_out=16'h12a;
17'h14f2d:	data_out=16'h8154;
17'h14f2e:	data_out=16'h8063;
17'h14f2f:	data_out=16'hc5;
17'h14f30:	data_out=16'ha4;
17'h14f31:	data_out=16'h8036;
17'h14f32:	data_out=16'h8a;
17'h14f33:	data_out=16'hc9;
17'h14f34:	data_out=16'h80c0;
17'h14f35:	data_out=16'h90;
17'h14f36:	data_out=16'h148;
17'h14f37:	data_out=16'h800c;
17'h14f38:	data_out=16'h16;
17'h14f39:	data_out=16'ha6;
17'h14f3a:	data_out=16'h2b;
17'h14f3b:	data_out=16'hcc;
17'h14f3c:	data_out=16'h80a9;
17'h14f3d:	data_out=16'hcc;
17'h14f3e:	data_out=16'h8010;
17'h14f3f:	data_out=16'h79;
17'h14f40:	data_out=16'h2b;
17'h14f41:	data_out=16'h86;
17'h14f42:	data_out=16'h80de;
17'h14f43:	data_out=16'h3e;
17'h14f44:	data_out=16'hc2;
17'h14f45:	data_out=16'h12f;
17'h14f46:	data_out=16'h80df;
17'h14f47:	data_out=16'h20;
17'h14f48:	data_out=16'h80d8;
17'h14f49:	data_out=16'h8004;
17'h14f4a:	data_out=16'h5b;
17'h14f4b:	data_out=16'h80d6;
17'h14f4c:	data_out=16'h8078;
17'h14f4d:	data_out=16'h801d;
17'h14f4e:	data_out=16'h8023;
17'h14f4f:	data_out=16'h8056;
17'h14f50:	data_out=16'h5f;
17'h14f51:	data_out=16'h119;
17'h14f52:	data_out=16'h8042;
17'h14f53:	data_out=16'h43;
17'h14f54:	data_out=16'h13d;
17'h14f55:	data_out=16'h71;
17'h14f56:	data_out=16'h60;
17'h14f57:	data_out=16'h8045;
17'h14f58:	data_out=16'h8019;
17'h14f59:	data_out=16'h801e;
17'h14f5a:	data_out=16'h814a;
17'h14f5b:	data_out=16'h1e1;
17'h14f5c:	data_out=16'ha6;
17'h14f5d:	data_out=16'h801e;
17'h14f5e:	data_out=16'hb8;
17'h14f5f:	data_out=16'h1a;
17'h14f60:	data_out=16'h80fd;
17'h14f61:	data_out=16'h179;
17'h14f62:	data_out=16'h3c;
17'h14f63:	data_out=16'hb8;
17'h14f64:	data_out=16'h808d;
17'h14f65:	data_out=16'h808f;
17'h14f66:	data_out=16'h8099;
17'h14f67:	data_out=16'h80b6;
17'h14f68:	data_out=16'h8011;
17'h14f69:	data_out=16'h8f;
17'h14f6a:	data_out=16'h8024;
17'h14f6b:	data_out=16'h97;
17'h14f6c:	data_out=16'h8009;
17'h14f6d:	data_out=16'hbb;
17'h14f6e:	data_out=16'h801d;
17'h14f6f:	data_out=16'h801f;
17'h14f70:	data_out=16'h801e;
17'h14f71:	data_out=16'h4e;
17'h14f72:	data_out=16'h801f;
17'h14f73:	data_out=16'ha7;
17'h14f74:	data_out=16'ha0;
17'h14f75:	data_out=16'h8003;
17'h14f76:	data_out=16'h8031;
17'h14f77:	data_out=16'h1f;
17'h14f78:	data_out=16'h44;
17'h14f79:	data_out=16'ha;
17'h14f7a:	data_out=16'hbe;
17'h14f7b:	data_out=16'h8017;
17'h14f7c:	data_out=16'ha7;
17'h14f7d:	data_out=16'h11e;
17'h14f7e:	data_out=16'h8013;
17'h14f7f:	data_out=16'h56;
17'h14f80:	data_out=16'h5;
17'h14f81:	data_out=16'h8009;
17'h14f82:	data_out=16'h8001;
17'h14f83:	data_out=16'h1;
17'h14f84:	data_out=16'h8008;
17'h14f85:	data_out=16'h8006;
17'h14f86:	data_out=16'h8001;
17'h14f87:	data_out=16'h8008;
17'h14f88:	data_out=16'h8005;
17'h14f89:	data_out=16'h5;
17'h14f8a:	data_out=16'h8000;
17'h14f8b:	data_out=16'h8008;
17'h14f8c:	data_out=16'h5;
17'h14f8d:	data_out=16'h8006;
17'h14f8e:	data_out=16'h5;
17'h14f8f:	data_out=16'h8004;
17'h14f90:	data_out=16'h5;
17'h14f91:	data_out=16'h6;
17'h14f92:	data_out=16'h8007;
17'h14f93:	data_out=16'h8000;
17'h14f94:	data_out=16'h8004;
17'h14f95:	data_out=16'h8005;
17'h14f96:	data_out=16'h8001;
17'h14f97:	data_out=16'h6;
17'h14f98:	data_out=16'h4;
17'h14f99:	data_out=16'h3;
17'h14f9a:	data_out=16'h8005;
17'h14f9b:	data_out=16'h8001;
17'h14f9c:	data_out=16'h9;
17'h14f9d:	data_out=16'h8009;
17'h14f9e:	data_out=16'h8000;
17'h14f9f:	data_out=16'h4;
17'h14fa0:	data_out=16'h8008;
17'h14fa1:	data_out=16'h8;
17'h14fa2:	data_out=16'h8003;
17'h14fa3:	data_out=16'h8007;
17'h14fa4:	data_out=16'h8006;
17'h14fa5:	data_out=16'h5;
17'h14fa6:	data_out=16'h8005;
17'h14fa7:	data_out=16'h8003;
17'h14fa8:	data_out=16'h1;
17'h14fa9:	data_out=16'h4;
17'h14faa:	data_out=16'h8001;
17'h14fab:	data_out=16'h8003;
17'h14fac:	data_out=16'h6;
17'h14fad:	data_out=16'h8006;
17'h14fae:	data_out=16'h1;
17'h14faf:	data_out=16'h2;
17'h14fb0:	data_out=16'h9;
17'h14fb1:	data_out=16'h4;
17'h14fb2:	data_out=16'h8007;
17'h14fb3:	data_out=16'h8004;
17'h14fb4:	data_out=16'h8;
17'h14fb5:	data_out=16'h1;
17'h14fb6:	data_out=16'h8007;
17'h14fb7:	data_out=16'h3;
17'h14fb8:	data_out=16'h8004;
17'h14fb9:	data_out=16'h8002;
17'h14fba:	data_out=16'h8008;
17'h14fbb:	data_out=16'h8005;
17'h14fbc:	data_out=16'h8002;
17'h14fbd:	data_out=16'h1;
17'h14fbe:	data_out=16'h9;
17'h14fbf:	data_out=16'h8001;
17'h14fc0:	data_out=16'h0;
17'h14fc1:	data_out=16'h8003;
17'h14fc2:	data_out=16'h1;
17'h14fc3:	data_out=16'h3;
17'h14fc4:	data_out=16'h8008;
17'h14fc5:	data_out=16'h5;
17'h14fc6:	data_out=16'h8009;
17'h14fc7:	data_out=16'h2;
17'h14fc8:	data_out=16'h8000;
17'h14fc9:	data_out=16'h8001;
17'h14fca:	data_out=16'h8;
17'h14fcb:	data_out=16'h8003;
17'h14fcc:	data_out=16'h3;
17'h14fcd:	data_out=16'h8000;
17'h14fce:	data_out=16'h8;
17'h14fcf:	data_out=16'h3;
17'h14fd0:	data_out=16'h8006;
17'h14fd1:	data_out=16'h8008;
17'h14fd2:	data_out=16'h8;
17'h14fd3:	data_out=16'h8007;
17'h14fd4:	data_out=16'h3;
17'h14fd5:	data_out=16'h8008;
17'h14fd6:	data_out=16'h5;
17'h14fd7:	data_out=16'h7;
17'h14fd8:	data_out=16'h8001;
17'h14fd9:	data_out=16'h6;
17'h14fda:	data_out=16'h8006;
17'h14fdb:	data_out=16'h6;
17'h14fdc:	data_out=16'h8002;
17'h14fdd:	data_out=16'h8007;
17'h14fde:	data_out=16'h8004;
17'h14fdf:	data_out=16'h8;
17'h14fe0:	data_out=16'h8001;
17'h14fe1:	data_out=16'h7;
17'h14fe2:	data_out=16'h2;
17'h14fe3:	data_out=16'h0;
17'h14fe4:	data_out=16'h2;
17'h14fe5:	data_out=16'h2;
17'h14fe6:	data_out=16'h8007;
17'h14fe7:	data_out=16'h8007;
17'h14fe8:	data_out=16'h8008;
17'h14fe9:	data_out=16'h8008;
17'h14fea:	data_out=16'h8001;
17'h14feb:	data_out=16'h4;
17'h14fec:	data_out=16'h0;
17'h14fed:	data_out=16'h8002;
17'h14fee:	data_out=16'h8003;
17'h14fef:	data_out=16'h4;
17'h14ff0:	data_out=16'h8001;
17'h14ff1:	data_out=16'h8004;
17'h14ff2:	data_out=16'h6;
17'h14ff3:	data_out=16'h8007;
17'h14ff4:	data_out=16'h8002;
17'h14ff5:	data_out=16'h1;
17'h14ff6:	data_out=16'h8009;
17'h14ff7:	data_out=16'h6;
17'h14ff8:	data_out=16'h8002;
17'h14ff9:	data_out=16'h8006;
17'h14ffa:	data_out=16'h3;
17'h14ffb:	data_out=16'h5;
17'h14ffc:	data_out=16'h8004;
17'h14ffd:	data_out=16'h8;
17'h14ffe:	data_out=16'h4;
17'h14fff:	data_out=16'h5;
17'h15000:	data_out=16'h6;
17'h15001:	data_out=16'h8004;
17'h15002:	data_out=16'h8004;
17'h15003:	data_out=16'h8001;
17'h15004:	data_out=16'h8;
17'h15005:	data_out=16'h8002;
17'h15006:	data_out=16'h1;
17'h15007:	data_out=16'h9;
17'h15008:	data_out=16'h8001;
17'h15009:	data_out=16'h9;
17'h1500a:	data_out=16'h4;
17'h1500b:	data_out=16'h8;
17'h1500c:	data_out=16'h8003;
17'h1500d:	data_out=16'h8008;
17'h1500e:	data_out=16'h3;
17'h1500f:	data_out=16'h6;
17'h15010:	data_out=16'h8003;
17'h15011:	data_out=16'h8000;
17'h15012:	data_out=16'h8;
17'h15013:	data_out=16'h4;
17'h15014:	data_out=16'h8008;
17'h15015:	data_out=16'h8;
17'h15016:	data_out=16'h0;
17'h15017:	data_out=16'h8001;
17'h15018:	data_out=16'h8007;
17'h15019:	data_out=16'h8006;
17'h1501a:	data_out=16'h8004;
17'h1501b:	data_out=16'h8002;
17'h1501c:	data_out=16'h8007;
17'h1501d:	data_out=16'h9;
17'h1501e:	data_out=16'h8007;
17'h1501f:	data_out=16'h8;
17'h15020:	data_out=16'h8004;
17'h15021:	data_out=16'h8002;
17'h15022:	data_out=16'h8002;
17'h15023:	data_out=16'h8006;
17'h15024:	data_out=16'h6;
17'h15025:	data_out=16'h8;
17'h15026:	data_out=16'h8006;
17'h15027:	data_out=16'h8005;
17'h15028:	data_out=16'h7;
17'h15029:	data_out=16'h7;
17'h1502a:	data_out=16'h8005;
17'h1502b:	data_out=16'h8004;
17'h1502c:	data_out=16'h8;
17'h1502d:	data_out=16'h7;
17'h1502e:	data_out=16'h8008;
17'h1502f:	data_out=16'h8004;
17'h15030:	data_out=16'h8003;
17'h15031:	data_out=16'h9;
17'h15032:	data_out=16'h9;
17'h15033:	data_out=16'h8001;
17'h15034:	data_out=16'h8;
17'h15035:	data_out=16'h0;
17'h15036:	data_out=16'h7;
17'h15037:	data_out=16'h8009;
17'h15038:	data_out=16'h3;
17'h15039:	data_out=16'h8006;
17'h1503a:	data_out=16'h8002;
17'h1503b:	data_out=16'h6;
17'h1503c:	data_out=16'h8007;
17'h1503d:	data_out=16'h1;
17'h1503e:	data_out=16'h5;
17'h1503f:	data_out=16'h8002;
17'h15040:	data_out=16'h8;
17'h15041:	data_out=16'h8006;
17'h15042:	data_out=16'h1;
17'h15043:	data_out=16'h5;
17'h15044:	data_out=16'h8008;
17'h15045:	data_out=16'h4;
17'h15046:	data_out=16'h9;
17'h15047:	data_out=16'h9;
17'h15048:	data_out=16'h2;
17'h15049:	data_out=16'h8005;
17'h1504a:	data_out=16'h8005;
17'h1504b:	data_out=16'h0;
17'h1504c:	data_out=16'h8008;
17'h1504d:	data_out=16'h8004;
17'h1504e:	data_out=16'h5;
17'h1504f:	data_out=16'h8001;
17'h15050:	data_out=16'h8004;
17'h15051:	data_out=16'h5;
17'h15052:	data_out=16'h7;
17'h15053:	data_out=16'h8005;
17'h15054:	data_out=16'h8004;
17'h15055:	data_out=16'h5;
17'h15056:	data_out=16'h8005;
17'h15057:	data_out=16'h9;
17'h15058:	data_out=16'h7;
17'h15059:	data_out=16'h3;
17'h1505a:	data_out=16'h6;
17'h1505b:	data_out=16'h8009;
17'h1505c:	data_out=16'h8006;
17'h1505d:	data_out=16'h1;
17'h1505e:	data_out=16'h8002;
17'h1505f:	data_out=16'h8007;
17'h15060:	data_out=16'h4;
17'h15061:	data_out=16'h9;
17'h15062:	data_out=16'h7;
17'h15063:	data_out=16'h5;
17'h15064:	data_out=16'h4;
17'h15065:	data_out=16'h7;
17'h15066:	data_out=16'h5;
17'h15067:	data_out=16'h8003;
17'h15068:	data_out=16'h8007;
17'h15069:	data_out=16'h9;
17'h1506a:	data_out=16'h7;
17'h1506b:	data_out=16'h8006;
17'h1506c:	data_out=16'h8004;
17'h1506d:	data_out=16'h3;
17'h1506e:	data_out=16'h2;
17'h1506f:	data_out=16'h2;
17'h15070:	data_out=16'h8001;
17'h15071:	data_out=16'h8000;
17'h15072:	data_out=16'h6;
17'h15073:	data_out=16'h4;
17'h15074:	data_out=16'h8005;
17'h15075:	data_out=16'h8008;
17'h15076:	data_out=16'h4;
17'h15077:	data_out=16'h8007;
17'h15078:	data_out=16'h4;
17'h15079:	data_out=16'h0;
17'h1507a:	data_out=16'h8006;
17'h1507b:	data_out=16'h8;
17'h1507c:	data_out=16'h8008;
17'h1507d:	data_out=16'h1;
17'h1507e:	data_out=16'h8008;
17'h1507f:	data_out=16'h6;
17'h15080:	data_out=16'h1;
17'h15081:	data_out=16'h8;
17'h15082:	data_out=16'h2;
17'h15083:	data_out=16'h8004;
17'h15084:	data_out=16'h6;
17'h15085:	data_out=16'h8003;
17'h15086:	data_out=16'h2;
17'h15087:	data_out=16'h8;
17'h15088:	data_out=16'h8003;
17'h15089:	data_out=16'h8000;
17'h1508a:	data_out=16'h8007;
17'h1508b:	data_out=16'h2;
17'h1508c:	data_out=16'h8006;
17'h1508d:	data_out=16'h4;
17'h1508e:	data_out=16'h8005;
17'h1508f:	data_out=16'h2;
17'h15090:	data_out=16'h8005;
17'h15091:	data_out=16'h8008;
17'h15092:	data_out=16'h8003;
17'h15093:	data_out=16'h8001;
17'h15094:	data_out=16'h8007;
17'h15095:	data_out=16'h8008;
17'h15096:	data_out=16'h2;
17'h15097:	data_out=16'h7;
17'h15098:	data_out=16'h1;
17'h15099:	data_out=16'h5;
17'h1509a:	data_out=16'h5;
17'h1509b:	data_out=16'h3;
17'h1509c:	data_out=16'h8003;
17'h1509d:	data_out=16'h6;
17'h1509e:	data_out=16'h8001;
17'h1509f:	data_out=16'h7;
17'h150a0:	data_out=16'h5;
17'h150a1:	data_out=16'h8008;
17'h150a2:	data_out=16'h8007;
17'h150a3:	data_out=16'h2;
17'h150a4:	data_out=16'h8002;
17'h150a5:	data_out=16'h5;
17'h150a6:	data_out=16'h1;
17'h150a7:	data_out=16'h4;
17'h150a8:	data_out=16'h8005;
17'h150a9:	data_out=16'h3;
17'h150aa:	data_out=16'h8002;
17'h150ab:	data_out=16'h8002;
17'h150ac:	data_out=16'h8002;
17'h150ad:	data_out=16'h2;
17'h150ae:	data_out=16'h9;
17'h150af:	data_out=16'h2;
17'h150b0:	data_out=16'h3;
17'h150b1:	data_out=16'h8003;
17'h150b2:	data_out=16'h8007;
17'h150b3:	data_out=16'h6;
17'h150b4:	data_out=16'h8003;
17'h150b5:	data_out=16'h4;
17'h150b6:	data_out=16'h3;
17'h150b7:	data_out=16'h8;
17'h150b8:	data_out=16'h8001;
17'h150b9:	data_out=16'h8001;
17'h150ba:	data_out=16'h2;
17'h150bb:	data_out=16'h5;
17'h150bc:	data_out=16'h8004;
17'h150bd:	data_out=16'h8008;
17'h150be:	data_out=16'h2;
17'h150bf:	data_out=16'h8009;
17'h150c0:	data_out=16'h8007;
17'h150c1:	data_out=16'h5;
17'h150c2:	data_out=16'h2;
17'h150c3:	data_out=16'h0;
17'h150c4:	data_out=16'h0;
17'h150c5:	data_out=16'h8006;
17'h150c6:	data_out=16'h8005;
17'h150c7:	data_out=16'h5;
17'h150c8:	data_out=16'h6;
17'h150c9:	data_out=16'h2;
17'h150ca:	data_out=16'h8007;
17'h150cb:	data_out=16'h8005;
17'h150cc:	data_out=16'h8005;
17'h150cd:	data_out=16'h8007;
17'h150ce:	data_out=16'h7;
17'h150cf:	data_out=16'h7;
17'h150d0:	data_out=16'h8001;
17'h150d1:	data_out=16'h9;
17'h150d2:	data_out=16'h4;
17'h150d3:	data_out=16'h5;
17'h150d4:	data_out=16'h3;
17'h150d5:	data_out=16'h8002;
17'h150d6:	data_out=16'h4;
17'h150d7:	data_out=16'h8007;
17'h150d8:	data_out=16'h6;
17'h150d9:	data_out=16'h8004;
17'h150da:	data_out=16'h7;
17'h150db:	data_out=16'h8008;
17'h150dc:	data_out=16'h8003;
17'h150dd:	data_out=16'h1;
17'h150de:	data_out=16'h8007;
17'h150df:	data_out=16'h8001;
17'h150e0:	data_out=16'h8004;
17'h150e1:	data_out=16'h4;
17'h150e2:	data_out=16'h9;
17'h150e3:	data_out=16'h6;
17'h150e4:	data_out=16'h7;
17'h150e5:	data_out=16'h8005;
17'h150e6:	data_out=16'h1;
17'h150e7:	data_out=16'h4;
17'h150e8:	data_out=16'h6;
17'h150e9:	data_out=16'h4;
17'h150ea:	data_out=16'h9;
17'h150eb:	data_out=16'h8008;
17'h150ec:	data_out=16'h6;
17'h150ed:	data_out=16'h6;
17'h150ee:	data_out=16'h8;
17'h150ef:	data_out=16'h8005;
17'h150f0:	data_out=16'h5;
17'h150f1:	data_out=16'h3;
17'h150f2:	data_out=16'h8009;
17'h150f3:	data_out=16'h8000;
17'h150f4:	data_out=16'h8008;
17'h150f5:	data_out=16'h5;
17'h150f6:	data_out=16'h2;
17'h150f7:	data_out=16'h7;
17'h150f8:	data_out=16'h8008;
17'h150f9:	data_out=16'h0;
17'h150fa:	data_out=16'h8;
17'h150fb:	data_out=16'h8002;
17'h150fc:	data_out=16'h8008;
17'h150fd:	data_out=16'h8008;
17'h150fe:	data_out=16'h7;
17'h150ff:	data_out=16'h8003;
17'h15100:	data_out=16'h18;
17'h15101:	data_out=16'h28;
17'h15102:	data_out=16'h87;
17'h15103:	data_out=16'h21;
17'h15104:	data_out=16'h80a4;
17'h15105:	data_out=16'he5;
17'h15106:	data_out=16'h11b;
17'h15107:	data_out=16'h803b;
17'h15108:	data_out=16'h100;
17'h15109:	data_out=16'h57;
17'h1510a:	data_out=16'h8001;
17'h1510b:	data_out=16'h7e;
17'h1510c:	data_out=16'h806c;
17'h1510d:	data_out=16'h8013;
17'h1510e:	data_out=16'h800f;
17'h1510f:	data_out=16'h3b;
17'h15110:	data_out=16'h8036;
17'h15111:	data_out=16'h801f;
17'h15112:	data_out=16'h96;
17'h15113:	data_out=16'h8012;
17'h15114:	data_out=16'he2;
17'h15115:	data_out=16'h80d3;
17'h15116:	data_out=16'h8085;
17'h15117:	data_out=16'hfd;
17'h15118:	data_out=16'h807f;
17'h15119:	data_out=16'h8076;
17'h1511a:	data_out=16'h8098;
17'h1511b:	data_out=16'h74;
17'h1511c:	data_out=16'hdd;
17'h1511d:	data_out=16'h95;
17'h1511e:	data_out=16'h137;
17'h1511f:	data_out=16'hbc;
17'h15120:	data_out=16'h10f;
17'h15121:	data_out=16'h8012;
17'h15122:	data_out=16'h51;
17'h15123:	data_out=16'h80f9;
17'h15124:	data_out=16'h80f9;
17'h15125:	data_out=16'h2d;
17'h15126:	data_out=16'h73;
17'h15127:	data_out=16'hb1;
17'h15128:	data_out=16'h8002;
17'h15129:	data_out=16'h807f;
17'h1512a:	data_out=16'h59;
17'h1512b:	data_out=16'h33;
17'h1512c:	data_out=16'h8032;
17'h1512d:	data_out=16'h80d2;
17'h1512e:	data_out=16'h5a;
17'h1512f:	data_out=16'he9;
17'h15130:	data_out=16'h805a;
17'h15131:	data_out=16'h84;
17'h15132:	data_out=16'h805d;
17'h15133:	data_out=16'hdc;
17'h15134:	data_out=16'h8071;
17'h15135:	data_out=16'h53;
17'h15136:	data_out=16'h1c0;
17'h15137:	data_out=16'ha9;
17'h15138:	data_out=16'hd4;
17'h15139:	data_out=16'h8f;
17'h1513a:	data_out=16'h14;
17'h1513b:	data_out=16'h800e;
17'h1513c:	data_out=16'h16b;
17'h1513d:	data_out=16'h8005;
17'h1513e:	data_out=16'h8008;
17'h1513f:	data_out=16'h15;
17'h15140:	data_out=16'h8010;
17'h15141:	data_out=16'h15a;
17'h15142:	data_out=16'h801f;
17'h15143:	data_out=16'ha0;
17'h15144:	data_out=16'h808c;
17'h15145:	data_out=16'h8105;
17'h15146:	data_out=16'hc9;
17'h15147:	data_out=16'h802f;
17'h15148:	data_out=16'h45;
17'h15149:	data_out=16'h16;
17'h1514a:	data_out=16'h80ca;
17'h1514b:	data_out=16'h801f;
17'h1514c:	data_out=16'h803c;
17'h1514d:	data_out=16'h5d;
17'h1514e:	data_out=16'h69;
17'h1514f:	data_out=16'h8071;
17'h15150:	data_out=16'h805d;
17'h15151:	data_out=16'h8019;
17'h15152:	data_out=16'h80d0;
17'h15153:	data_out=16'hd1;
17'h15154:	data_out=16'he4;
17'h15155:	data_out=16'h12e;
17'h15156:	data_out=16'h74;
17'h15157:	data_out=16'h43;
17'h15158:	data_out=16'ha1;
17'h15159:	data_out=16'h28;
17'h1515a:	data_out=16'hb0;
17'h1515b:	data_out=16'h12b;
17'h1515c:	data_out=16'h5f;
17'h1515d:	data_out=16'h1d;
17'h1515e:	data_out=16'h122;
17'h1515f:	data_out=16'h9;
17'h15160:	data_out=16'h8065;
17'h15161:	data_out=16'h803d;
17'h15162:	data_out=16'h1d1;
17'h15163:	data_out=16'hbc;
17'h15164:	data_out=16'h80a2;
17'h15165:	data_out=16'h8077;
17'h15166:	data_out=16'h8083;
17'h15167:	data_out=16'h3c;
17'h15168:	data_out=16'h800d;
17'h15169:	data_out=16'hf6;
17'h1516a:	data_out=16'h8006;
17'h1516b:	data_out=16'h52;
17'h1516c:	data_out=16'h5b;
17'h1516d:	data_out=16'hdf;
17'h1516e:	data_out=16'h8016;
17'h1516f:	data_out=16'h48;
17'h15170:	data_out=16'h8012;
17'h15171:	data_out=16'h8019;
17'h15172:	data_out=16'h8055;
17'h15173:	data_out=16'h10;
17'h15174:	data_out=16'h8055;
17'h15175:	data_out=16'ha0;
17'h15176:	data_out=16'h6c;
17'h15177:	data_out=16'h80e3;
17'h15178:	data_out=16'h63;
17'h15179:	data_out=16'h96;
17'h1517a:	data_out=16'hf2;
17'h1517b:	data_out=16'h800f;
17'h1517c:	data_out=16'h41;
17'h1517d:	data_out=16'h14b;
17'h1517e:	data_out=16'h7b;
17'h1517f:	data_out=16'h80eb;
17'h15180:	data_out=16'h89fb;
17'h15181:	data_out=16'h28f;
17'h15182:	data_out=16'h129;
17'h15183:	data_out=16'h8588;
17'h15184:	data_out=16'h836b;
17'h15185:	data_out=16'h677;
17'h15186:	data_out=16'h8007;
17'h15187:	data_out=16'h8537;
17'h15188:	data_out=16'h2e2;
17'h15189:	data_out=16'h8a00;
17'h1518a:	data_out=16'h8482;
17'h1518b:	data_out=16'h77d;
17'h1518c:	data_out=16'h9fb;
17'h1518d:	data_out=16'h8034;
17'h1518e:	data_out=16'h8192;
17'h1518f:	data_out=16'hb7;
17'h15190:	data_out=16'h8618;
17'h15191:	data_out=16'h54c;
17'h15192:	data_out=16'h8262;
17'h15193:	data_out=16'h860f;
17'h15194:	data_out=16'h283;
17'h15195:	data_out=16'h839f;
17'h15196:	data_out=16'h8564;
17'h15197:	data_out=16'h2ad;
17'h15198:	data_out=16'h816e;
17'h15199:	data_out=16'h786;
17'h1519a:	data_out=16'h820b;
17'h1519b:	data_out=16'ha00;
17'h1519c:	data_out=16'h2ed;
17'h1519d:	data_out=16'h48f;
17'h1519e:	data_out=16'h22f;
17'h1519f:	data_out=16'h82c4;
17'h151a0:	data_out=16'h5f3;
17'h151a1:	data_out=16'h817e;
17'h151a2:	data_out=16'h8a00;
17'h151a3:	data_out=16'h836c;
17'h151a4:	data_out=16'h8369;
17'h151a5:	data_out=16'h88b2;
17'h151a6:	data_out=16'h88f4;
17'h151a7:	data_out=16'h907;
17'h151a8:	data_out=16'h8129;
17'h151a9:	data_out=16'h85b8;
17'h151aa:	data_out=16'h87c8;
17'h151ab:	data_out=16'ha00;
17'h151ac:	data_out=16'h850c;
17'h151ad:	data_out=16'h8a00;
17'h151ae:	data_out=16'h81c8;
17'h151af:	data_out=16'h3e5;
17'h151b0:	data_out=16'h8186;
17'h151b1:	data_out=16'h5d5;
17'h151b2:	data_out=16'h82a4;
17'h151b3:	data_out=16'h2c2;
17'h151b4:	data_out=16'h811f;
17'h151b5:	data_out=16'h9fd;
17'h151b6:	data_out=16'h481;
17'h151b7:	data_out=16'h204;
17'h151b8:	data_out=16'h20f;
17'h151b9:	data_out=16'h318;
17'h151ba:	data_out=16'h8a00;
17'h151bb:	data_out=16'h371;
17'h151bc:	data_out=16'h631;
17'h151bd:	data_out=16'h89b0;
17'h151be:	data_out=16'h8123;
17'h151bf:	data_out=16'h685;
17'h151c0:	data_out=16'h89ff;
17'h151c1:	data_out=16'ha00;
17'h151c2:	data_out=16'h8915;
17'h151c3:	data_out=16'h10a;
17'h151c4:	data_out=16'h2ec;
17'h151c5:	data_out=16'h83bd;
17'h151c6:	data_out=16'h1bd;
17'h151c7:	data_out=16'h8a00;
17'h151c8:	data_out=16'h804c;
17'h151c9:	data_out=16'h88a7;
17'h151ca:	data_out=16'h80f4;
17'h151cb:	data_out=16'h3a2;
17'h151cc:	data_out=16'h8a00;
17'h151cd:	data_out=16'h8a00;
17'h151ce:	data_out=16'h80db;
17'h151cf:	data_out=16'h8a00;
17'h151d0:	data_out=16'h8a00;
17'h151d1:	data_out=16'h4d7;
17'h151d2:	data_out=16'h873a;
17'h151d3:	data_out=16'ha00;
17'h151d4:	data_out=16'h289;
17'h151d5:	data_out=16'h5ee;
17'h151d6:	data_out=16'h8a00;
17'h151d7:	data_out=16'h89fe;
17'h151d8:	data_out=16'h3b2;
17'h151d9:	data_out=16'h8a00;
17'h151da:	data_out=16'ha00;
17'h151db:	data_out=16'h8c3;
17'h151dc:	data_out=16'ha00;
17'h151dd:	data_out=16'h8533;
17'h151de:	data_out=16'h2c5;
17'h151df:	data_out=16'h8042;
17'h151e0:	data_out=16'h8a00;
17'h151e1:	data_out=16'h523;
17'h151e2:	data_out=16'h6d6;
17'h151e3:	data_out=16'h3cf;
17'h151e4:	data_out=16'h4f;
17'h151e5:	data_out=16'hfb;
17'h151e6:	data_out=16'h7db;
17'h151e7:	data_out=16'h85d4;
17'h151e8:	data_out=16'h8160;
17'h151e9:	data_out=16'h219;
17'h151ea:	data_out=16'h81a2;
17'h151eb:	data_out=16'h80b4;
17'h151ec:	data_out=16'h89fc;
17'h151ed:	data_out=16'h36c;
17'h151ee:	data_out=16'h81a2;
17'h151ef:	data_out=16'h849e;
17'h151f0:	data_out=16'h8198;
17'h151f1:	data_out=16'h101;
17'h151f2:	data_out=16'h8a00;
17'h151f3:	data_out=16'h8669;
17'h151f4:	data_out=16'h816d;
17'h151f5:	data_out=16'h9ff;
17'h151f6:	data_out=16'h7a0;
17'h151f7:	data_out=16'h8a00;
17'h151f8:	data_out=16'h4;
17'h151f9:	data_out=16'h8112;
17'h151fa:	data_out=16'h34e;
17'h151fb:	data_out=16'h8116;
17'h151fc:	data_out=16'h1;
17'h151fd:	data_out=16'h4a9;
17'h151fe:	data_out=16'h8a00;
17'h151ff:	data_out=16'h89ff;
17'h15200:	data_out=16'h89f7;
17'h15201:	data_out=16'h308;
17'h15202:	data_out=16'h347;
17'h15203:	data_out=16'h8a00;
17'h15204:	data_out=16'h8a00;
17'h15205:	data_out=16'h86b6;
17'h15206:	data_out=16'h8a00;
17'h15207:	data_out=16'h89de;
17'h15208:	data_out=16'ha00;
17'h15209:	data_out=16'h8a00;
17'h1520a:	data_out=16'h8a00;
17'h1520b:	data_out=16'h9fe;
17'h1520c:	data_out=16'h71a;
17'h1520d:	data_out=16'h26f;
17'h1520e:	data_out=16'h8600;
17'h1520f:	data_out=16'h81b7;
17'h15210:	data_out=16'hb6;
17'h15211:	data_out=16'h89fa;
17'h15212:	data_out=16'h4a;
17'h15213:	data_out=16'h8a00;
17'h15214:	data_out=16'h9f4;
17'h15215:	data_out=16'h8a00;
17'h15216:	data_out=16'h8a00;
17'h15217:	data_out=16'h9f8;
17'h15218:	data_out=16'h8313;
17'h15219:	data_out=16'h9ff;
17'h1521a:	data_out=16'h89fb;
17'h1521b:	data_out=16'ha00;
17'h1521c:	data_out=16'h8933;
17'h1521d:	data_out=16'h438;
17'h1521e:	data_out=16'h7b4;
17'h1521f:	data_out=16'h8750;
17'h15220:	data_out=16'ha00;
17'h15221:	data_out=16'h85b7;
17'h15222:	data_out=16'h8a00;
17'h15223:	data_out=16'h8a00;
17'h15224:	data_out=16'h8a00;
17'h15225:	data_out=16'h8a00;
17'h15226:	data_out=16'h8a00;
17'h15227:	data_out=16'h9ff;
17'h15228:	data_out=16'h853e;
17'h15229:	data_out=16'hf2;
17'h1522a:	data_out=16'h89f4;
17'h1522b:	data_out=16'ha00;
17'h1522c:	data_out=16'h8a00;
17'h1522d:	data_out=16'h8a00;
17'h1522e:	data_out=16'h74b;
17'h1522f:	data_out=16'ha00;
17'h15230:	data_out=16'h8a00;
17'h15231:	data_out=16'h993;
17'h15232:	data_out=16'h8a00;
17'h15233:	data_out=16'ha00;
17'h15234:	data_out=16'h89fd;
17'h15235:	data_out=16'h83c;
17'h15236:	data_out=16'ha00;
17'h15237:	data_out=16'h414;
17'h15238:	data_out=16'h8923;
17'h15239:	data_out=16'ha00;
17'h1523a:	data_out=16'h8a00;
17'h1523b:	data_out=16'h8899;
17'h1523c:	data_out=16'h9fe;
17'h1523d:	data_out=16'h8a00;
17'h1523e:	data_out=16'h853a;
17'h1523f:	data_out=16'h86ef;
17'h15240:	data_out=16'h8a00;
17'h15241:	data_out=16'ha00;
17'h15242:	data_out=16'h898f;
17'h15243:	data_out=16'h880a;
17'h15244:	data_out=16'h8759;
17'h15245:	data_out=16'h8a00;
17'h15246:	data_out=16'ha00;
17'h15247:	data_out=16'h8a00;
17'h15248:	data_out=16'h9ed;
17'h15249:	data_out=16'h8a00;
17'h1524a:	data_out=16'h5ad;
17'h1524b:	data_out=16'h8bf;
17'h1524c:	data_out=16'h8a00;
17'h1524d:	data_out=16'h8a00;
17'h1524e:	data_out=16'h1d9;
17'h1524f:	data_out=16'h8a00;
17'h15250:	data_out=16'h8a00;
17'h15251:	data_out=16'h8261;
17'h15252:	data_out=16'h8a00;
17'h15253:	data_out=16'ha00;
17'h15254:	data_out=16'ha00;
17'h15255:	data_out=16'h72e;
17'h15256:	data_out=16'h8a00;
17'h15257:	data_out=16'h8a00;
17'h15258:	data_out=16'ha00;
17'h15259:	data_out=16'h8a00;
17'h1525a:	data_out=16'ha00;
17'h1525b:	data_out=16'h8344;
17'h1525c:	data_out=16'ha00;
17'h1525d:	data_out=16'h878f;
17'h1525e:	data_out=16'h9f5;
17'h1525f:	data_out=16'h1f3;
17'h15260:	data_out=16'h8a00;
17'h15261:	data_out=16'h8a00;
17'h15262:	data_out=16'h9d8;
17'h15263:	data_out=16'ha00;
17'h15264:	data_out=16'h8411;
17'h15265:	data_out=16'h85a4;
17'h15266:	data_out=16'h9f6;
17'h15267:	data_out=16'h85ef;
17'h15268:	data_out=16'h858b;
17'h15269:	data_out=16'ha00;
17'h1526a:	data_out=16'h8639;
17'h1526b:	data_out=16'h8a00;
17'h1526c:	data_out=16'h89fb;
17'h1526d:	data_out=16'ha00;
17'h1526e:	data_out=16'h8638;
17'h1526f:	data_out=16'h8a00;
17'h15270:	data_out=16'h8618;
17'h15271:	data_out=16'h824d;
17'h15272:	data_out=16'h8a00;
17'h15273:	data_out=16'h8a00;
17'h15274:	data_out=16'h8a00;
17'h15275:	data_out=16'ha00;
17'h15276:	data_out=16'h9f7;
17'h15277:	data_out=16'h8a00;
17'h15278:	data_out=16'h89f8;
17'h15279:	data_out=16'h4d5;
17'h1527a:	data_out=16'h9ff;
17'h1527b:	data_out=16'h8539;
17'h1527c:	data_out=16'h1d6;
17'h1527d:	data_out=16'h862f;
17'h1527e:	data_out=16'h8a00;
17'h1527f:	data_out=16'h8a00;
17'h15280:	data_out=16'h809e;
17'h15281:	data_out=16'hd5;
17'h15282:	data_out=16'h8315;
17'h15283:	data_out=16'h8213;
17'h15284:	data_out=16'h8a00;
17'h15285:	data_out=16'h89ff;
17'h15286:	data_out=16'h8a00;
17'h15287:	data_out=16'h8a00;
17'h15288:	data_out=16'ha00;
17'h15289:	data_out=16'h8a00;
17'h1528a:	data_out=16'h8a00;
17'h1528b:	data_out=16'h9fd;
17'h1528c:	data_out=16'h87e0;
17'h1528d:	data_out=16'ha00;
17'h1528e:	data_out=16'h8a00;
17'h1528f:	data_out=16'h87c4;
17'h15290:	data_out=16'h3f2;
17'h15291:	data_out=16'h8a00;
17'h15292:	data_out=16'h148;
17'h15293:	data_out=16'h8a00;
17'h15294:	data_out=16'h9ea;
17'h15295:	data_out=16'h8a00;
17'h15296:	data_out=16'h8a00;
17'h15297:	data_out=16'h9f0;
17'h15298:	data_out=16'h8411;
17'h15299:	data_out=16'h87ed;
17'h1529a:	data_out=16'h8a00;
17'h1529b:	data_out=16'ha00;
17'h1529c:	data_out=16'h854f;
17'h1529d:	data_out=16'h8650;
17'h1529e:	data_out=16'h98c;
17'h1529f:	data_out=16'h8a00;
17'h152a0:	data_out=16'ha00;
17'h152a1:	data_out=16'h8a00;
17'h152a2:	data_out=16'h8a00;
17'h152a3:	data_out=16'h8a00;
17'h152a4:	data_out=16'h8a00;
17'h152a5:	data_out=16'h8a00;
17'h152a6:	data_out=16'h8a00;
17'h152a7:	data_out=16'h9d5;
17'h152a8:	data_out=16'h8a00;
17'h152a9:	data_out=16'h9e0;
17'h152aa:	data_out=16'h8197;
17'h152ab:	data_out=16'ha00;
17'h152ac:	data_out=16'h8a00;
17'h152ad:	data_out=16'h8a00;
17'h152ae:	data_out=16'h8ae;
17'h152af:	data_out=16'ha00;
17'h152b0:	data_out=16'h8a00;
17'h152b1:	data_out=16'h81a5;
17'h152b2:	data_out=16'h8a00;
17'h152b3:	data_out=16'ha00;
17'h152b4:	data_out=16'h8a00;
17'h152b5:	data_out=16'h8a00;
17'h152b6:	data_out=16'ha00;
17'h152b7:	data_out=16'h8309;
17'h152b8:	data_out=16'h89a2;
17'h152b9:	data_out=16'ha00;
17'h152ba:	data_out=16'h8a00;
17'h152bb:	data_out=16'h89ff;
17'h152bc:	data_out=16'h9bf;
17'h152bd:	data_out=16'h8a00;
17'h152be:	data_out=16'h8a00;
17'h152bf:	data_out=16'h89ff;
17'h152c0:	data_out=16'h8a00;
17'h152c1:	data_out=16'ha00;
17'h152c2:	data_out=16'h8a00;
17'h152c3:	data_out=16'h89ff;
17'h152c4:	data_out=16'h89fe;
17'h152c5:	data_out=16'h8a00;
17'h152c6:	data_out=16'h9f2;
17'h152c7:	data_out=16'h8a00;
17'h152c8:	data_out=16'h973;
17'h152c9:	data_out=16'h8a00;
17'h152ca:	data_out=16'ha00;
17'h152cb:	data_out=16'h83f;
17'h152cc:	data_out=16'h8a00;
17'h152cd:	data_out=16'h8a00;
17'h152ce:	data_out=16'h410;
17'h152cf:	data_out=16'h8a00;
17'h152d0:	data_out=16'h8a00;
17'h152d1:	data_out=16'h89fc;
17'h152d2:	data_out=16'h8a00;
17'h152d3:	data_out=16'h9ff;
17'h152d4:	data_out=16'h9ff;
17'h152d5:	data_out=16'h28c;
17'h152d6:	data_out=16'h89f9;
17'h152d7:	data_out=16'h8a00;
17'h152d8:	data_out=16'ha00;
17'h152d9:	data_out=16'h8a00;
17'h152da:	data_out=16'ha00;
17'h152db:	data_out=16'h8a00;
17'h152dc:	data_out=16'h9fe;
17'h152dd:	data_out=16'h8448;
17'h152de:	data_out=16'h9fa;
17'h152df:	data_out=16'h838;
17'h152e0:	data_out=16'h8a00;
17'h152e1:	data_out=16'h8a00;
17'h152e2:	data_out=16'h9db;
17'h152e3:	data_out=16'ha00;
17'h152e4:	data_out=16'h89f8;
17'h152e5:	data_out=16'h8a00;
17'h152e6:	data_out=16'h896b;
17'h152e7:	data_out=16'h87ec;
17'h152e8:	data_out=16'h8a00;
17'h152e9:	data_out=16'ha00;
17'h152ea:	data_out=16'h8a00;
17'h152eb:	data_out=16'h8a00;
17'h152ec:	data_out=16'h89d3;
17'h152ed:	data_out=16'ha00;
17'h152ee:	data_out=16'h8a00;
17'h152ef:	data_out=16'h8a00;
17'h152f0:	data_out=16'h8a00;
17'h152f1:	data_out=16'h414;
17'h152f2:	data_out=16'h8a00;
17'h152f3:	data_out=16'h8a00;
17'h152f4:	data_out=16'h8a00;
17'h152f5:	data_out=16'h1fd;
17'h152f6:	data_out=16'h3e2;
17'h152f7:	data_out=16'h8a00;
17'h152f8:	data_out=16'h89fd;
17'h152f9:	data_out=16'ha00;
17'h152fa:	data_out=16'h9fb;
17'h152fb:	data_out=16'h8a00;
17'h152fc:	data_out=16'h442;
17'h152fd:	data_out=16'h89ff;
17'h152fe:	data_out=16'h8a00;
17'h152ff:	data_out=16'h89fd;
17'h15300:	data_out=16'h8069;
17'h15301:	data_out=16'h89fd;
17'h15302:	data_out=16'h8a00;
17'h15303:	data_out=16'h446;
17'h15304:	data_out=16'h8a00;
17'h15305:	data_out=16'h89fd;
17'h15306:	data_out=16'h8a00;
17'h15307:	data_out=16'h8a00;
17'h15308:	data_out=16'ha00;
17'h15309:	data_out=16'h8a00;
17'h1530a:	data_out=16'h8a00;
17'h1530b:	data_out=16'h9ff;
17'h1530c:	data_out=16'h8a00;
17'h1530d:	data_out=16'h9f7;
17'h1530e:	data_out=16'h8a00;
17'h1530f:	data_out=16'h8a00;
17'h15310:	data_out=16'h8247;
17'h15311:	data_out=16'h89ac;
17'h15312:	data_out=16'h451;
17'h15313:	data_out=16'h8a00;
17'h15314:	data_out=16'h9f1;
17'h15315:	data_out=16'h8a00;
17'h15316:	data_out=16'h8a00;
17'h15317:	data_out=16'h9ed;
17'h15318:	data_out=16'h8743;
17'h15319:	data_out=16'h89ec;
17'h1531a:	data_out=16'h8a00;
17'h1531b:	data_out=16'h9fb;
17'h1531c:	data_out=16'h80e5;
17'h1531d:	data_out=16'h8a00;
17'h1531e:	data_out=16'h858;
17'h1531f:	data_out=16'h8a00;
17'h15320:	data_out=16'ha00;
17'h15321:	data_out=16'h8a00;
17'h15322:	data_out=16'h8a00;
17'h15323:	data_out=16'h8a00;
17'h15324:	data_out=16'h8a00;
17'h15325:	data_out=16'h8a00;
17'h15326:	data_out=16'h8a00;
17'h15327:	data_out=16'h421;
17'h15328:	data_out=16'h8a00;
17'h15329:	data_out=16'h9d0;
17'h1532a:	data_out=16'h879d;
17'h1532b:	data_out=16'ha00;
17'h1532c:	data_out=16'h8a00;
17'h1532d:	data_out=16'h8a00;
17'h1532e:	data_out=16'h722;
17'h1532f:	data_out=16'ha00;
17'h15330:	data_out=16'h8a00;
17'h15331:	data_out=16'h8020;
17'h15332:	data_out=16'h8a00;
17'h15333:	data_out=16'ha00;
17'h15334:	data_out=16'h8a00;
17'h15335:	data_out=16'h8a00;
17'h15336:	data_out=16'h9ff;
17'h15337:	data_out=16'h8a00;
17'h15338:	data_out=16'h873e;
17'h15339:	data_out=16'ha00;
17'h1533a:	data_out=16'h8a00;
17'h1533b:	data_out=16'h8a00;
17'h1533c:	data_out=16'ha00;
17'h1533d:	data_out=16'h89fd;
17'h1533e:	data_out=16'h8a00;
17'h1533f:	data_out=16'h89fd;
17'h15340:	data_out=16'h8a00;
17'h15341:	data_out=16'ha00;
17'h15342:	data_out=16'h8a00;
17'h15343:	data_out=16'h84b8;
17'h15344:	data_out=16'h89e3;
17'h15345:	data_out=16'h8a00;
17'h15346:	data_out=16'h93d;
17'h15347:	data_out=16'h8a00;
17'h15348:	data_out=16'h7ca;
17'h15349:	data_out=16'h8a00;
17'h1534a:	data_out=16'h9ff;
17'h1534b:	data_out=16'h51f;
17'h1534c:	data_out=16'h8a00;
17'h1534d:	data_out=16'h8a00;
17'h1534e:	data_out=16'h8138;
17'h1534f:	data_out=16'h8a00;
17'h15350:	data_out=16'h8a00;
17'h15351:	data_out=16'h89fb;
17'h15352:	data_out=16'h8a00;
17'h15353:	data_out=16'h9ff;
17'h15354:	data_out=16'h9ff;
17'h15355:	data_out=16'h8151;
17'h15356:	data_out=16'h89ff;
17'h15357:	data_out=16'h8a00;
17'h15358:	data_out=16'h3d4;
17'h15359:	data_out=16'h8a00;
17'h1535a:	data_out=16'ha00;
17'h1535b:	data_out=16'h89fe;
17'h1535c:	data_out=16'h9f6;
17'h1535d:	data_out=16'h8a00;
17'h1535e:	data_out=16'h9fa;
17'h1535f:	data_out=16'h48e;
17'h15360:	data_out=16'h8a00;
17'h15361:	data_out=16'h8a00;
17'h15362:	data_out=16'h9dc;
17'h15363:	data_out=16'ha00;
17'h15364:	data_out=16'h89f7;
17'h15365:	data_out=16'h8a00;
17'h15366:	data_out=16'h8a00;
17'h15367:	data_out=16'h89fc;
17'h15368:	data_out=16'h8a00;
17'h15369:	data_out=16'ha00;
17'h1536a:	data_out=16'h8a00;
17'h1536b:	data_out=16'h8a00;
17'h1536c:	data_out=16'h89f3;
17'h1536d:	data_out=16'ha00;
17'h1536e:	data_out=16'h8a00;
17'h1536f:	data_out=16'h8a00;
17'h15370:	data_out=16'h8a00;
17'h15371:	data_out=16'h8e1;
17'h15372:	data_out=16'h8a00;
17'h15373:	data_out=16'h8a00;
17'h15374:	data_out=16'h8a00;
17'h15375:	data_out=16'h805d;
17'h15376:	data_out=16'h8c7;
17'h15377:	data_out=16'h8a00;
17'h15378:	data_out=16'h89e5;
17'h15379:	data_out=16'ha00;
17'h1537a:	data_out=16'h9fb;
17'h1537b:	data_out=16'h8a00;
17'h1537c:	data_out=16'h1aa;
17'h1537d:	data_out=16'h89dc;
17'h1537e:	data_out=16'h89ff;
17'h1537f:	data_out=16'h89fc;
17'h15380:	data_out=16'h2e1;
17'h15381:	data_out=16'h89f9;
17'h15382:	data_out=16'h89b2;
17'h15383:	data_out=16'h580;
17'h15384:	data_out=16'h8a00;
17'h15385:	data_out=16'h89de;
17'h15386:	data_out=16'h8a00;
17'h15387:	data_out=16'h8a00;
17'h15388:	data_out=16'h9ff;
17'h15389:	data_out=16'h8a00;
17'h1538a:	data_out=16'h8a00;
17'h1538b:	data_out=16'h9f9;
17'h1538c:	data_out=16'h8a00;
17'h1538d:	data_out=16'h9ea;
17'h1538e:	data_out=16'h89ff;
17'h1538f:	data_out=16'h8a00;
17'h15390:	data_out=16'h89ff;
17'h15391:	data_out=16'h870c;
17'h15392:	data_out=16'h51c;
17'h15393:	data_out=16'h8a00;
17'h15394:	data_out=16'h9d7;
17'h15395:	data_out=16'h8a00;
17'h15396:	data_out=16'h8a00;
17'h15397:	data_out=16'h9cf;
17'h15398:	data_out=16'h859e;
17'h15399:	data_out=16'h89f6;
17'h1539a:	data_out=16'h89fb;
17'h1539b:	data_out=16'h9f6;
17'h1539c:	data_out=16'h932;
17'h1539d:	data_out=16'h89ff;
17'h1539e:	data_out=16'h60c;
17'h1539f:	data_out=16'h880f;
17'h153a0:	data_out=16'h9d6;
17'h153a1:	data_out=16'h89ff;
17'h153a2:	data_out=16'h8a00;
17'h153a3:	data_out=16'h89f9;
17'h153a4:	data_out=16'h89f9;
17'h153a5:	data_out=16'h8a00;
17'h153a6:	data_out=16'h89ff;
17'h153a7:	data_out=16'h5b5;
17'h153a8:	data_out=16'h89ff;
17'h153a9:	data_out=16'h9e9;
17'h153aa:	data_out=16'h8a00;
17'h153ab:	data_out=16'h9ef;
17'h153ac:	data_out=16'h8a00;
17'h153ad:	data_out=16'h8a00;
17'h153ae:	data_out=16'h61;
17'h153af:	data_out=16'h9e8;
17'h153b0:	data_out=16'h8a00;
17'h153b1:	data_out=16'h74b;
17'h153b2:	data_out=16'h8a00;
17'h153b3:	data_out=16'h9f3;
17'h153b4:	data_out=16'h89fe;
17'h153b5:	data_out=16'h8871;
17'h153b6:	data_out=16'h9f3;
17'h153b7:	data_out=16'h88b2;
17'h153b8:	data_out=16'h8822;
17'h153b9:	data_out=16'h9f9;
17'h153ba:	data_out=16'h8a00;
17'h153bb:	data_out=16'h89ff;
17'h153bc:	data_out=16'ha00;
17'h153bd:	data_out=16'h8a00;
17'h153be:	data_out=16'h89ff;
17'h153bf:	data_out=16'h89e1;
17'h153c0:	data_out=16'h8a00;
17'h153c1:	data_out=16'h9fe;
17'h153c2:	data_out=16'h8a00;
17'h153c3:	data_out=16'h2a0;
17'h153c4:	data_out=16'h852e;
17'h153c5:	data_out=16'h8a00;
17'h153c6:	data_out=16'h9f9;
17'h153c7:	data_out=16'h8a00;
17'h153c8:	data_out=16'h8303;
17'h153c9:	data_out=16'h8a00;
17'h153ca:	data_out=16'h9e8;
17'h153cb:	data_out=16'h8461;
17'h153cc:	data_out=16'h8a00;
17'h153cd:	data_out=16'h8a00;
17'h153ce:	data_out=16'h81b7;
17'h153cf:	data_out=16'h8a00;
17'h153d0:	data_out=16'h8a00;
17'h153d1:	data_out=16'h5d1;
17'h153d2:	data_out=16'h8a00;
17'h153d3:	data_out=16'h9fe;
17'h153d4:	data_out=16'h96e;
17'h153d5:	data_out=16'h82a3;
17'h153d6:	data_out=16'h89ee;
17'h153d7:	data_out=16'h8a00;
17'h153d8:	data_out=16'ha00;
17'h153d9:	data_out=16'h8a00;
17'h153da:	data_out=16'h9fc;
17'h153db:	data_out=16'h89fc;
17'h153dc:	data_out=16'h9f9;
17'h153dd:	data_out=16'h8a00;
17'h153de:	data_out=16'h9ca;
17'h153df:	data_out=16'h8625;
17'h153e0:	data_out=16'h8a00;
17'h153e1:	data_out=16'h89fe;
17'h153e2:	data_out=16'h54f;
17'h153e3:	data_out=16'h9f2;
17'h153e4:	data_out=16'h89f2;
17'h153e5:	data_out=16'h8a00;
17'h153e6:	data_out=16'h8a00;
17'h153e7:	data_out=16'h8a00;
17'h153e8:	data_out=16'h89ff;
17'h153e9:	data_out=16'h9fe;
17'h153ea:	data_out=16'h89fe;
17'h153eb:	data_out=16'h89ff;
17'h153ec:	data_out=16'h89f1;
17'h153ed:	data_out=16'h9f2;
17'h153ee:	data_out=16'h89fe;
17'h153ef:	data_out=16'h8a00;
17'h153f0:	data_out=16'h89fe;
17'h153f1:	data_out=16'h4a3;
17'h153f2:	data_out=16'h8a00;
17'h153f3:	data_out=16'h8a00;
17'h153f4:	data_out=16'h8a00;
17'h153f5:	data_out=16'h9dc;
17'h153f6:	data_out=16'h89a0;
17'h153f7:	data_out=16'h8a00;
17'h153f8:	data_out=16'h8941;
17'h153f9:	data_out=16'h9fd;
17'h153fa:	data_out=16'h9e3;
17'h153fb:	data_out=16'h89ff;
17'h153fc:	data_out=16'h35f;
17'h153fd:	data_out=16'h89fc;
17'h153fe:	data_out=16'h89fe;
17'h153ff:	data_out=16'h89f4;
17'h15400:	data_out=16'h85b7;
17'h15401:	data_out=16'h88ae;
17'h15402:	data_out=16'h9bf;
17'h15403:	data_out=16'h571;
17'h15404:	data_out=16'h89f1;
17'h15405:	data_out=16'h8828;
17'h15406:	data_out=16'h8a00;
17'h15407:	data_out=16'h8a00;
17'h15408:	data_out=16'h9f9;
17'h15409:	data_out=16'h8a00;
17'h1540a:	data_out=16'h89f8;
17'h1540b:	data_out=16'h9f5;
17'h1540c:	data_out=16'h8a00;
17'h1540d:	data_out=16'h941;
17'h1540e:	data_out=16'h866f;
17'h1540f:	data_out=16'h2f6;
17'h15410:	data_out=16'h8a00;
17'h15411:	data_out=16'hea;
17'h15412:	data_out=16'h3b7;
17'h15413:	data_out=16'h8a00;
17'h15414:	data_out=16'h9af;
17'h15415:	data_out=16'h89fe;
17'h15416:	data_out=16'h8a00;
17'h15417:	data_out=16'h98a;
17'h15418:	data_out=16'h8794;
17'h15419:	data_out=16'h89c9;
17'h1541a:	data_out=16'h89dd;
17'h1541b:	data_out=16'h9f8;
17'h1541c:	data_out=16'h9ff;
17'h1541d:	data_out=16'h89d9;
17'h1541e:	data_out=16'h683;
17'h1541f:	data_out=16'h86bd;
17'h15420:	data_out=16'h8df;
17'h15421:	data_out=16'h8611;
17'h15422:	data_out=16'h8a00;
17'h15423:	data_out=16'h89ea;
17'h15424:	data_out=16'h89e9;
17'h15425:	data_out=16'h8a00;
17'h15426:	data_out=16'h8968;
17'h15427:	data_out=16'hd6;
17'h15428:	data_out=16'h84ff;
17'h15429:	data_out=16'h9fb;
17'h1542a:	data_out=16'h8a00;
17'h1542b:	data_out=16'h9df;
17'h1542c:	data_out=16'h8a00;
17'h1542d:	data_out=16'h8a00;
17'h1542e:	data_out=16'h285;
17'h1542f:	data_out=16'h9bd;
17'h15430:	data_out=16'h89fe;
17'h15431:	data_out=16'h9f2;
17'h15432:	data_out=16'h89f7;
17'h15433:	data_out=16'h9db;
17'h15434:	data_out=16'h89fa;
17'h15435:	data_out=16'h8374;
17'h15436:	data_out=16'h9ce;
17'h15437:	data_out=16'h9c5;
17'h15438:	data_out=16'h80fa;
17'h15439:	data_out=16'h9e4;
17'h1543a:	data_out=16'h8a00;
17'h1543b:	data_out=16'h884e;
17'h1543c:	data_out=16'ha00;
17'h1543d:	data_out=16'h89fe;
17'h1543e:	data_out=16'h84f3;
17'h1543f:	data_out=16'h8861;
17'h15440:	data_out=16'h89fe;
17'h15441:	data_out=16'h9f9;
17'h15442:	data_out=16'h8a00;
17'h15443:	data_out=16'h9e7;
17'h15444:	data_out=16'h8172;
17'h15445:	data_out=16'h89fe;
17'h15446:	data_out=16'h9fc;
17'h15447:	data_out=16'h8a00;
17'h15448:	data_out=16'h8a00;
17'h15449:	data_out=16'h8a00;
17'h1544a:	data_out=16'h9ce;
17'h1544b:	data_out=16'h83d4;
17'h1544c:	data_out=16'h8a00;
17'h1544d:	data_out=16'h8a00;
17'h1544e:	data_out=16'h3c;
17'h1544f:	data_out=16'h8a00;
17'h15450:	data_out=16'h8a00;
17'h15451:	data_out=16'h9c0;
17'h15452:	data_out=16'h89fd;
17'h15453:	data_out=16'h9fe;
17'h15454:	data_out=16'h266;
17'h15455:	data_out=16'h3ca;
17'h15456:	data_out=16'h8994;
17'h15457:	data_out=16'h89f5;
17'h15458:	data_out=16'ha00;
17'h15459:	data_out=16'h89fe;
17'h1545a:	data_out=16'h9f3;
17'h1545b:	data_out=16'h849d;
17'h1545c:	data_out=16'ha00;
17'h1545d:	data_out=16'h8a00;
17'h1545e:	data_out=16'h33d;
17'h1545f:	data_out=16'h8a00;
17'h15460:	data_out=16'h8a00;
17'h15461:	data_out=16'h89f0;
17'h15462:	data_out=16'h60b;
17'h15463:	data_out=16'h9da;
17'h15464:	data_out=16'h89f0;
17'h15465:	data_out=16'h89fd;
17'h15466:	data_out=16'h89f7;
17'h15467:	data_out=16'h8653;
17'h15468:	data_out=16'h85c9;
17'h15469:	data_out=16'h9f7;
17'h1546a:	data_out=16'h86b6;
17'h1546b:	data_out=16'h89fd;
17'h1546c:	data_out=16'h89f3;
17'h1546d:	data_out=16'h9da;
17'h1546e:	data_out=16'h86b6;
17'h1546f:	data_out=16'h89fe;
17'h15470:	data_out=16'h8685;
17'h15471:	data_out=16'h5cb;
17'h15472:	data_out=16'h89ff;
17'h15473:	data_out=16'h89fe;
17'h15474:	data_out=16'h89fe;
17'h15475:	data_out=16'h9f3;
17'h15476:	data_out=16'h89f2;
17'h15477:	data_out=16'h8a00;
17'h15478:	data_out=16'h856a;
17'h15479:	data_out=16'h9ee;
17'h1547a:	data_out=16'h9c3;
17'h1547b:	data_out=16'h84ed;
17'h1547c:	data_out=16'h81d9;
17'h1547d:	data_out=16'h89fa;
17'h1547e:	data_out=16'h89ff;
17'h1547f:	data_out=16'h89fd;
17'h15480:	data_out=16'h84dc;
17'h15481:	data_out=16'h821c;
17'h15482:	data_out=16'h9cf;
17'h15483:	data_out=16'h8481;
17'h15484:	data_out=16'h8958;
17'h15485:	data_out=16'h8120;
17'h15486:	data_out=16'h8a00;
17'h15487:	data_out=16'h8a00;
17'h15488:	data_out=16'h9f5;
17'h15489:	data_out=16'h8a00;
17'h1548a:	data_out=16'h89e5;
17'h1548b:	data_out=16'h9be;
17'h1548c:	data_out=16'h8a00;
17'h1548d:	data_out=16'h706;
17'h1548e:	data_out=16'ha00;
17'h1548f:	data_out=16'h8f2;
17'h15490:	data_out=16'h8a00;
17'h15491:	data_out=16'ha00;
17'h15492:	data_out=16'h763;
17'h15493:	data_out=16'h8a00;
17'h15494:	data_out=16'h93f;
17'h15495:	data_out=16'h89fa;
17'h15496:	data_out=16'h8a00;
17'h15497:	data_out=16'h8a3;
17'h15498:	data_out=16'h862b;
17'h15499:	data_out=16'h89a2;
17'h1549a:	data_out=16'h87a7;
17'h1549b:	data_out=16'h9f2;
17'h1549c:	data_out=16'h9f2;
17'h1549d:	data_out=16'h881f;
17'h1549e:	data_out=16'h85d;
17'h1549f:	data_out=16'h15e;
17'h154a0:	data_out=16'h14;
17'h154a1:	data_out=16'ha00;
17'h154a2:	data_out=16'h8a00;
17'h154a3:	data_out=16'h818f;
17'h154a4:	data_out=16'h8177;
17'h154a5:	data_out=16'h8a00;
17'h154a6:	data_out=16'h9da;
17'h154a7:	data_out=16'h9fa;
17'h154a8:	data_out=16'ha00;
17'h154a9:	data_out=16'h9f4;
17'h154aa:	data_out=16'h71b;
17'h154ab:	data_out=16'h84ca;
17'h154ac:	data_out=16'h8a00;
17'h154ad:	data_out=16'h8a00;
17'h154ae:	data_out=16'h74b;
17'h154af:	data_out=16'h8f8;
17'h154b0:	data_out=16'h89ef;
17'h154b1:	data_out=16'h900;
17'h154b2:	data_out=16'h8834;
17'h154b3:	data_out=16'h972;
17'h154b4:	data_out=16'h89d2;
17'h154b5:	data_out=16'h9d7;
17'h154b6:	data_out=16'h9cb;
17'h154b7:	data_out=16'h9e3;
17'h154b8:	data_out=16'h63c;
17'h154b9:	data_out=16'h96b;
17'h154ba:	data_out=16'h8a00;
17'h154bb:	data_out=16'h8121;
17'h154bc:	data_out=16'ha00;
17'h154bd:	data_out=16'h89f3;
17'h154be:	data_out=16'ha00;
17'h154bf:	data_out=16'h819e;
17'h154c0:	data_out=16'h89e9;
17'h154c1:	data_out=16'h9d9;
17'h154c2:	data_out=16'h89f6;
17'h154c3:	data_out=16'h9d8;
17'h154c4:	data_out=16'h82f;
17'h154c5:	data_out=16'h89fa;
17'h154c6:	data_out=16'h9fe;
17'h154c7:	data_out=16'h8a00;
17'h154c8:	data_out=16'h8a00;
17'h154c9:	data_out=16'h8a00;
17'h154ca:	data_out=16'h9c1;
17'h154cb:	data_out=16'h8318;
17'h154cc:	data_out=16'h8a00;
17'h154cd:	data_out=16'h8a00;
17'h154ce:	data_out=16'h564;
17'h154cf:	data_out=16'h8a00;
17'h154d0:	data_out=16'h8a00;
17'h154d1:	data_out=16'h9a4;
17'h154d2:	data_out=16'h89f1;
17'h154d3:	data_out=16'ha00;
17'h154d4:	data_out=16'h81cc;
17'h154d5:	data_out=16'h988;
17'h154d6:	data_out=16'h8580;
17'h154d7:	data_out=16'h899e;
17'h154d8:	data_out=16'h9f5;
17'h154d9:	data_out=16'h89ed;
17'h154da:	data_out=16'h9dc;
17'h154db:	data_out=16'ha00;
17'h154dc:	data_out=16'ha00;
17'h154dd:	data_out=16'h8a00;
17'h154de:	data_out=16'h812c;
17'h154df:	data_out=16'h8a00;
17'h154e0:	data_out=16'h89fb;
17'h154e1:	data_out=16'h8640;
17'h154e2:	data_out=16'h44d;
17'h154e3:	data_out=16'h98d;
17'h154e4:	data_out=16'h89ee;
17'h154e5:	data_out=16'h89e5;
17'h154e6:	data_out=16'h89e6;
17'h154e7:	data_out=16'h8533;
17'h154e8:	data_out=16'ha00;
17'h154e9:	data_out=16'h9ef;
17'h154ea:	data_out=16'ha00;
17'h154eb:	data_out=16'h89fd;
17'h154ec:	data_out=16'h89e4;
17'h154ed:	data_out=16'h97d;
17'h154ee:	data_out=16'ha00;
17'h154ef:	data_out=16'h89fd;
17'h154f0:	data_out=16'ha00;
17'h154f1:	data_out=16'h898;
17'h154f2:	data_out=16'h89fc;
17'h154f3:	data_out=16'h89f1;
17'h154f4:	data_out=16'h89e0;
17'h154f5:	data_out=16'ha00;
17'h154f6:	data_out=16'h89d3;
17'h154f7:	data_out=16'h8a00;
17'h154f8:	data_out=16'h875c;
17'h154f9:	data_out=16'h9d2;
17'h154fa:	data_out=16'h970;
17'h154fb:	data_out=16'ha00;
17'h154fc:	data_out=16'h821c;
17'h154fd:	data_out=16'h88ad;
17'h154fe:	data_out=16'h898b;
17'h154ff:	data_out=16'h8a00;
17'h15500:	data_out=16'h89e3;
17'h15501:	data_out=16'hab;
17'h15502:	data_out=16'h9f7;
17'h15503:	data_out=16'h8a00;
17'h15504:	data_out=16'h8890;
17'h15505:	data_out=16'h83ba;
17'h15506:	data_out=16'h8a00;
17'h15507:	data_out=16'h89ff;
17'h15508:	data_out=16'h9fb;
17'h15509:	data_out=16'h8a00;
17'h1550a:	data_out=16'h8982;
17'h1550b:	data_out=16'h9df;
17'h1550c:	data_out=16'h8a00;
17'h1550d:	data_out=16'h8a00;
17'h1550e:	data_out=16'ha00;
17'h1550f:	data_out=16'h94a;
17'h15510:	data_out=16'h8a00;
17'h15511:	data_out=16'ha00;
17'h15512:	data_out=16'h71d;
17'h15513:	data_out=16'h8a00;
17'h15514:	data_out=16'h8ed;
17'h15515:	data_out=16'h89fc;
17'h15516:	data_out=16'h8a00;
17'h15517:	data_out=16'h821;
17'h15518:	data_out=16'h882b;
17'h15519:	data_out=16'h8922;
17'h1551a:	data_out=16'h84c3;
17'h1551b:	data_out=16'h9fd;
17'h1551c:	data_out=16'h9cd;
17'h1551d:	data_out=16'h80f5;
17'h1551e:	data_out=16'h796;
17'h1551f:	data_out=16'h3ce;
17'h15520:	data_out=16'h8912;
17'h15521:	data_out=16'ha00;
17'h15522:	data_out=16'h89eb;
17'h15523:	data_out=16'h8890;
17'h15524:	data_out=16'h886a;
17'h15525:	data_out=16'h89e4;
17'h15526:	data_out=16'h9f9;
17'h15527:	data_out=16'h9fe;
17'h15528:	data_out=16'ha00;
17'h15529:	data_out=16'ha00;
17'h1552a:	data_out=16'h924;
17'h1552b:	data_out=16'h842f;
17'h1552c:	data_out=16'h8a00;
17'h1552d:	data_out=16'h869c;
17'h1552e:	data_out=16'h9b0;
17'h1552f:	data_out=16'h231;
17'h15530:	data_out=16'h884f;
17'h15531:	data_out=16'h8302;
17'h15532:	data_out=16'h81e5;
17'h15533:	data_out=16'h8e2;
17'h15534:	data_out=16'h8884;
17'h15535:	data_out=16'h9b2;
17'h15536:	data_out=16'h9f4;
17'h15537:	data_out=16'ha00;
17'h15538:	data_out=16'h577;
17'h15539:	data_out=16'h885;
17'h1553a:	data_out=16'h8a00;
17'h1553b:	data_out=16'h14c;
17'h1553c:	data_out=16'ha00;
17'h1553d:	data_out=16'h89d7;
17'h1553e:	data_out=16'ha00;
17'h1553f:	data_out=16'h83d1;
17'h15540:	data_out=16'h894c;
17'h15541:	data_out=16'h9a9;
17'h15542:	data_out=16'h89ae;
17'h15543:	data_out=16'h9e8;
17'h15544:	data_out=16'h81f8;
17'h15545:	data_out=16'h89fd;
17'h15546:	data_out=16'ha00;
17'h15547:	data_out=16'h8a00;
17'h15548:	data_out=16'h8a00;
17'h15549:	data_out=16'h89d0;
17'h1554a:	data_out=16'h9f9;
17'h1554b:	data_out=16'h80cc;
17'h1554c:	data_out=16'h8a00;
17'h1554d:	data_out=16'h89e9;
17'h1554e:	data_out=16'ha00;
17'h1554f:	data_out=16'h8a00;
17'h15550:	data_out=16'h8a00;
17'h15551:	data_out=16'h925;
17'h15552:	data_out=16'h89ef;
17'h15553:	data_out=16'ha00;
17'h15554:	data_out=16'h87d3;
17'h15555:	data_out=16'h9b1;
17'h15556:	data_out=16'h9fc;
17'h15557:	data_out=16'h8757;
17'h15558:	data_out=16'h9f5;
17'h15559:	data_out=16'h899e;
17'h1555a:	data_out=16'h9de;
17'h1555b:	data_out=16'h9ff;
17'h1555c:	data_out=16'ha00;
17'h1555d:	data_out=16'h89e1;
17'h1555e:	data_out=16'h864f;
17'h1555f:	data_out=16'h89fb;
17'h15560:	data_out=16'h687;
17'h15561:	data_out=16'hd1;
17'h15562:	data_out=16'h7b6;
17'h15563:	data_out=16'h931;
17'h15564:	data_out=16'h89f7;
17'h15565:	data_out=16'h87a2;
17'h15566:	data_out=16'h89aa;
17'h15567:	data_out=16'h837;
17'h15568:	data_out=16'ha00;
17'h15569:	data_out=16'h9a9;
17'h1556a:	data_out=16'ha00;
17'h1556b:	data_out=16'h89ec;
17'h1556c:	data_out=16'h89dd;
17'h1556d:	data_out=16'h919;
17'h1556e:	data_out=16'ha00;
17'h1556f:	data_out=16'h89e4;
17'h15570:	data_out=16'ha00;
17'h15571:	data_out=16'h8e9;
17'h15572:	data_out=16'h89d5;
17'h15573:	data_out=16'h897c;
17'h15574:	data_out=16'h8789;
17'h15575:	data_out=16'ha00;
17'h15576:	data_out=16'h68c;
17'h15577:	data_out=16'h8a00;
17'h15578:	data_out=16'h231;
17'h15579:	data_out=16'h99b;
17'h1557a:	data_out=16'h938;
17'h1557b:	data_out=16'ha00;
17'h1557c:	data_out=16'h853f;
17'h1557d:	data_out=16'h8980;
17'h1557e:	data_out=16'h8417;
17'h1557f:	data_out=16'h8a00;
17'h15580:	data_out=16'h89db;
17'h15581:	data_out=16'ha00;
17'h15582:	data_out=16'ha00;
17'h15583:	data_out=16'h8a00;
17'h15584:	data_out=16'h8905;
17'h15585:	data_out=16'h83fd;
17'h15586:	data_out=16'h8a00;
17'h15587:	data_out=16'h89ff;
17'h15588:	data_out=16'h9f8;
17'h15589:	data_out=16'h8a00;
17'h1558a:	data_out=16'h893e;
17'h1558b:	data_out=16'h930;
17'h1558c:	data_out=16'h8837;
17'h1558d:	data_out=16'h8a00;
17'h1558e:	data_out=16'ha00;
17'h1558f:	data_out=16'h99e;
17'h15590:	data_out=16'h8a00;
17'h15591:	data_out=16'ha00;
17'h15592:	data_out=16'h729;
17'h15593:	data_out=16'h8a00;
17'h15594:	data_out=16'h466;
17'h15595:	data_out=16'h89f9;
17'h15596:	data_out=16'h8a00;
17'h15597:	data_out=16'h6ac;
17'h15598:	data_out=16'h819b;
17'h15599:	data_out=16'h889d;
17'h1559a:	data_out=16'h84f0;
17'h1559b:	data_out=16'h9ed;
17'h1559c:	data_out=16'h968;
17'h1559d:	data_out=16'ha00;
17'h1559e:	data_out=16'h29e;
17'h1559f:	data_out=16'h91;
17'h155a0:	data_out=16'h89b9;
17'h155a1:	data_out=16'ha00;
17'h155a2:	data_out=16'h89e4;
17'h155a3:	data_out=16'h82d2;
17'h155a4:	data_out=16'h82c3;
17'h155a5:	data_out=16'h89e1;
17'h155a6:	data_out=16'h9ee;
17'h155a7:	data_out=16'h9ff;
17'h155a8:	data_out=16'ha00;
17'h155a9:	data_out=16'ha00;
17'h155aa:	data_out=16'h9bb;
17'h155ab:	data_out=16'h88c3;
17'h155ac:	data_out=16'h8a00;
17'h155ad:	data_out=16'ha00;
17'h155ae:	data_out=16'h9f7;
17'h155af:	data_out=16'h892e;
17'h155b0:	data_out=16'h8436;
17'h155b1:	data_out=16'h84dc;
17'h155b2:	data_out=16'hda;
17'h155b3:	data_out=16'h58a;
17'h155b4:	data_out=16'h8617;
17'h155b5:	data_out=16'h9fb;
17'h155b6:	data_out=16'h9f6;
17'h155b7:	data_out=16'ha00;
17'h155b8:	data_out=16'h412;
17'h155b9:	data_out=16'h221;
17'h155ba:	data_out=16'h8a00;
17'h155bb:	data_out=16'hdc;
17'h155bc:	data_out=16'ha00;
17'h155bd:	data_out=16'h89c7;
17'h155be:	data_out=16'ha00;
17'h155bf:	data_out=16'h8412;
17'h155c0:	data_out=16'h8842;
17'h155c1:	data_out=16'h952;
17'h155c2:	data_out=16'h8313;
17'h155c3:	data_out=16'h9ec;
17'h155c4:	data_out=16'h821e;
17'h155c5:	data_out=16'h89f9;
17'h155c6:	data_out=16'ha00;
17'h155c7:	data_out=16'h8a00;
17'h155c8:	data_out=16'h8a00;
17'h155c9:	data_out=16'h8994;
17'h155ca:	data_out=16'h9fd;
17'h155cb:	data_out=16'h852e;
17'h155cc:	data_out=16'h89f6;
17'h155cd:	data_out=16'h89ea;
17'h155ce:	data_out=16'ha00;
17'h155cf:	data_out=16'h89f8;
17'h155d0:	data_out=16'h8a00;
17'h155d1:	data_out=16'h8bd;
17'h155d2:	data_out=16'h8895;
17'h155d3:	data_out=16'ha00;
17'h155d4:	data_out=16'h899d;
17'h155d5:	data_out=16'h9e2;
17'h155d6:	data_out=16'h9fc;
17'h155d7:	data_out=16'h9d5;
17'h155d8:	data_out=16'h9da;
17'h155d9:	data_out=16'h88ec;
17'h155da:	data_out=16'h9de;
17'h155db:	data_out=16'h9fd;
17'h155dc:	data_out=16'ha00;
17'h155dd:	data_out=16'h89ca;
17'h155de:	data_out=16'h89ca;
17'h155df:	data_out=16'h89ef;
17'h155e0:	data_out=16'h9ef;
17'h155e1:	data_out=16'h9ff;
17'h155e2:	data_out=16'h58f;
17'h155e3:	data_out=16'h8df;
17'h155e4:	data_out=16'h89fb;
17'h155e5:	data_out=16'h86e2;
17'h155e6:	data_out=16'h89eb;
17'h155e7:	data_out=16'h9ff;
17'h155e8:	data_out=16'ha00;
17'h155e9:	data_out=16'h953;
17'h155ea:	data_out=16'ha00;
17'h155eb:	data_out=16'h89dc;
17'h155ec:	data_out=16'h89c8;
17'h155ed:	data_out=16'h8bb;
17'h155ee:	data_out=16'ha00;
17'h155ef:	data_out=16'h89da;
17'h155f0:	data_out=16'ha00;
17'h155f1:	data_out=16'h9b6;
17'h155f2:	data_out=16'h89ab;
17'h155f3:	data_out=16'h878e;
17'h155f4:	data_out=16'h8120;
17'h155f5:	data_out=16'h9fd;
17'h155f6:	data_out=16'h12e;
17'h155f7:	data_out=16'h8a00;
17'h155f8:	data_out=16'h9fa;
17'h155f9:	data_out=16'h982;
17'h155fa:	data_out=16'h8f7;
17'h155fb:	data_out=16'ha00;
17'h155fc:	data_out=16'h8518;
17'h155fd:	data_out=16'h89e1;
17'h155fe:	data_out=16'h82ef;
17'h155ff:	data_out=16'h8a00;
17'h15600:	data_out=16'h8913;
17'h15601:	data_out=16'ha00;
17'h15602:	data_out=16'h9ff;
17'h15603:	data_out=16'h8a00;
17'h15604:	data_out=16'h89c9;
17'h15605:	data_out=16'h8323;
17'h15606:	data_out=16'h8a00;
17'h15607:	data_out=16'h2a7;
17'h15608:	data_out=16'h9c6;
17'h15609:	data_out=16'h8a00;
17'h1560a:	data_out=16'h895d;
17'h1560b:	data_out=16'h9d6;
17'h1560c:	data_out=16'h151;
17'h1560d:	data_out=16'h8a00;
17'h1560e:	data_out=16'ha00;
17'h1560f:	data_out=16'h9ad;
17'h15610:	data_out=16'h89ff;
17'h15611:	data_out=16'ha00;
17'h15612:	data_out=16'h786;
17'h15613:	data_out=16'h8a00;
17'h15614:	data_out=16'h8544;
17'h15615:	data_out=16'h89ff;
17'h15616:	data_out=16'h8a00;
17'h15617:	data_out=16'h84f6;
17'h15618:	data_out=16'h809d;
17'h15619:	data_out=16'h85b;
17'h1561a:	data_out=16'h88bd;
17'h1561b:	data_out=16'h9fc;
17'h1561c:	data_out=16'h86e;
17'h1561d:	data_out=16'ha00;
17'h1561e:	data_out=16'h8646;
17'h1561f:	data_out=16'h899c;
17'h15620:	data_out=16'h89d8;
17'h15621:	data_out=16'ha00;
17'h15622:	data_out=16'h89c9;
17'h15623:	data_out=16'h604;
17'h15624:	data_out=16'h60e;
17'h15625:	data_out=16'h89cd;
17'h15626:	data_out=16'h9ec;
17'h15627:	data_out=16'h9ff;
17'h15628:	data_out=16'ha00;
17'h15629:	data_out=16'ha00;
17'h1562a:	data_out=16'h9c3;
17'h1562b:	data_out=16'h886d;
17'h1562c:	data_out=16'h8a00;
17'h1562d:	data_out=16'ha00;
17'h1562e:	data_out=16'ha00;
17'h1562f:	data_out=16'h8962;
17'h15630:	data_out=16'h9d4;
17'h15631:	data_out=16'h82a6;
17'h15632:	data_out=16'h9f8;
17'h15633:	data_out=16'h87e9;
17'h15634:	data_out=16'h58a;
17'h15635:	data_out=16'h9ee;
17'h15636:	data_out=16'h9d6;
17'h15637:	data_out=16'ha00;
17'h15638:	data_out=16'h82;
17'h15639:	data_out=16'h89f7;
17'h1563a:	data_out=16'h8a00;
17'h1563b:	data_out=16'h9a9;
17'h1563c:	data_out=16'ha00;
17'h1563d:	data_out=16'h89d9;
17'h1563e:	data_out=16'ha00;
17'h1563f:	data_out=16'h83a1;
17'h15640:	data_out=16'h89ce;
17'h15641:	data_out=16'h97d;
17'h15642:	data_out=16'h82fd;
17'h15643:	data_out=16'h838;
17'h15644:	data_out=16'h95e;
17'h15645:	data_out=16'h8a00;
17'h15646:	data_out=16'ha00;
17'h15647:	data_out=16'h89f8;
17'h15648:	data_out=16'h8a00;
17'h15649:	data_out=16'h89ce;
17'h1564a:	data_out=16'h9c8;
17'h1564b:	data_out=16'h857c;
17'h1564c:	data_out=16'h89d9;
17'h1564d:	data_out=16'h89e2;
17'h1564e:	data_out=16'ha00;
17'h1564f:	data_out=16'h89ea;
17'h15650:	data_out=16'h8a00;
17'h15651:	data_out=16'h5a8;
17'h15652:	data_out=16'h650;
17'h15653:	data_out=16'ha00;
17'h15654:	data_out=16'h8742;
17'h15655:	data_out=16'h9cb;
17'h15656:	data_out=16'h9ee;
17'h15657:	data_out=16'h9ef;
17'h15658:	data_out=16'h995;
17'h15659:	data_out=16'h898f;
17'h1565a:	data_out=16'h9da;
17'h1565b:	data_out=16'h9e7;
17'h1565c:	data_out=16'h9fc;
17'h1565d:	data_out=16'h8699;
17'h1565e:	data_out=16'h89ed;
17'h1565f:	data_out=16'h89d4;
17'h15660:	data_out=16'h9f4;
17'h15661:	data_out=16'h9f6;
17'h15662:	data_out=16'h210;
17'h15663:	data_out=16'h1ae;
17'h15664:	data_out=16'h89f3;
17'h15665:	data_out=16'h8792;
17'h15666:	data_out=16'h89e6;
17'h15667:	data_out=16'ha00;
17'h15668:	data_out=16'ha00;
17'h15669:	data_out=16'h959;
17'h1566a:	data_out=16'ha00;
17'h1566b:	data_out=16'h8a00;
17'h1566c:	data_out=16'h85d9;
17'h1566d:	data_out=16'h812d;
17'h1566e:	data_out=16'ha00;
17'h1566f:	data_out=16'h8a00;
17'h15670:	data_out=16'ha00;
17'h15671:	data_out=16'h9bd;
17'h15672:	data_out=16'h89c6;
17'h15673:	data_out=16'h640;
17'h15674:	data_out=16'h9d5;
17'h15675:	data_out=16'h9c8;
17'h15676:	data_out=16'h9fe;
17'h15677:	data_out=16'h8a00;
17'h15678:	data_out=16'h9ec;
17'h15679:	data_out=16'h9b8;
17'h1567a:	data_out=16'h2d2;
17'h1567b:	data_out=16'ha00;
17'h1567c:	data_out=16'h842f;
17'h1567d:	data_out=16'h89e6;
17'h1567e:	data_out=16'h82c0;
17'h1567f:	data_out=16'h8a00;
17'h15680:	data_out=16'h8129;
17'h15681:	data_out=16'h9f2;
17'h15682:	data_out=16'h9ff;
17'h15683:	data_out=16'h8a00;
17'h15684:	data_out=16'h8a00;
17'h15685:	data_out=16'h89f8;
17'h15686:	data_out=16'h8a00;
17'h15687:	data_out=16'hbe;
17'h15688:	data_out=16'h9b7;
17'h15689:	data_out=16'h89e7;
17'h1568a:	data_out=16'h82e7;
17'h1568b:	data_out=16'h575;
17'h1568c:	data_out=16'h82f7;
17'h1568d:	data_out=16'h8a00;
17'h1568e:	data_out=16'ha00;
17'h1568f:	data_out=16'h9dd;
17'h15690:	data_out=16'h89f6;
17'h15691:	data_out=16'h9e9;
17'h15692:	data_out=16'h994;
17'h15693:	data_out=16'h8a00;
17'h15694:	data_out=16'h89e5;
17'h15695:	data_out=16'h8a00;
17'h15696:	data_out=16'h8a00;
17'h15697:	data_out=16'h8955;
17'h15698:	data_out=16'h780;
17'h15699:	data_out=16'h9dd;
17'h1569a:	data_out=16'h89f7;
17'h1569b:	data_out=16'h9f9;
17'h1569c:	data_out=16'h7aa;
17'h1569d:	data_out=16'h9db;
17'h1569e:	data_out=16'h816f;
17'h1569f:	data_out=16'h899a;
17'h156a0:	data_out=16'h89d0;
17'h156a1:	data_out=16'ha00;
17'h156a2:	data_out=16'h89ac;
17'h156a3:	data_out=16'h8538;
17'h156a4:	data_out=16'h8564;
17'h156a5:	data_out=16'h89bd;
17'h156a6:	data_out=16'h9ae;
17'h156a7:	data_out=16'h9c2;
17'h156a8:	data_out=16'ha00;
17'h156a9:	data_out=16'ha00;
17'h156aa:	data_out=16'h9f2;
17'h156ab:	data_out=16'h89d3;
17'h156ac:	data_out=16'h8a00;
17'h156ad:	data_out=16'ha00;
17'h156ae:	data_out=16'ha00;
17'h156af:	data_out=16'hc8;
17'h156b0:	data_out=16'h8d1;
17'h156b1:	data_out=16'h8089;
17'h156b2:	data_out=16'h77f;
17'h156b3:	data_out=16'h8463;
17'h156b4:	data_out=16'h9d6;
17'h156b5:	data_out=16'h609;
17'h156b6:	data_out=16'h9dc;
17'h156b7:	data_out=16'ha00;
17'h156b8:	data_out=16'h3cd;
17'h156b9:	data_out=16'h863f;
17'h156ba:	data_out=16'h89e4;
17'h156bb:	data_out=16'h4bc;
17'h156bc:	data_out=16'h9e0;
17'h156bd:	data_out=16'h89dc;
17'h156be:	data_out=16'ha00;
17'h156bf:	data_out=16'h89f8;
17'h156c0:	data_out=16'h8a00;
17'h156c1:	data_out=16'h9cf;
17'h156c2:	data_out=16'h89bb;
17'h156c3:	data_out=16'h3;
17'h156c4:	data_out=16'h387;
17'h156c5:	data_out=16'h8a00;
17'h156c6:	data_out=16'ha00;
17'h156c7:	data_out=16'h89bd;
17'h156c8:	data_out=16'h89ff;
17'h156c9:	data_out=16'h89c4;
17'h156ca:	data_out=16'h98d;
17'h156cb:	data_out=16'h8970;
17'h156cc:	data_out=16'h89a4;
17'h156cd:	data_out=16'h89c3;
17'h156ce:	data_out=16'ha00;
17'h156cf:	data_out=16'h89c7;
17'h156d0:	data_out=16'h8a00;
17'h156d1:	data_out=16'h1fc;
17'h156d2:	data_out=16'h88c3;
17'h156d3:	data_out=16'h9ef;
17'h156d4:	data_out=16'h858;
17'h156d5:	data_out=16'h758;
17'h156d6:	data_out=16'h808;
17'h156d7:	data_out=16'h5e5;
17'h156d8:	data_out=16'h9b0;
17'h156d9:	data_out=16'h89d1;
17'h156da:	data_out=16'h9f6;
17'h156db:	data_out=16'h607;
17'h156dc:	data_out=16'h9de;
17'h156dd:	data_out=16'h6d1;
17'h156de:	data_out=16'h89d0;
17'h156df:	data_out=16'h606;
17'h156e0:	data_out=16'h9e4;
17'h156e1:	data_out=16'h9bf;
17'h156e2:	data_out=16'h812b;
17'h156e3:	data_out=16'hb3;
17'h156e4:	data_out=16'h8349;
17'h156e5:	data_out=16'h89b2;
17'h156e6:	data_out=16'h89e5;
17'h156e7:	data_out=16'ha00;
17'h156e8:	data_out=16'ha00;
17'h156e9:	data_out=16'h98e;
17'h156ea:	data_out=16'ha00;
17'h156eb:	data_out=16'h8a00;
17'h156ec:	data_out=16'h9d6;
17'h156ed:	data_out=16'h8047;
17'h156ee:	data_out=16'ha00;
17'h156ef:	data_out=16'h8a00;
17'h156f0:	data_out=16'ha00;
17'h156f1:	data_out=16'h9e1;
17'h156f2:	data_out=16'h89fd;
17'h156f3:	data_out=16'h232;
17'h156f4:	data_out=16'h8d6;
17'h156f5:	data_out=16'h996;
17'h156f6:	data_out=16'h9a1;
17'h156f7:	data_out=16'h89de;
17'h156f8:	data_out=16'h947;
17'h156f9:	data_out=16'ha00;
17'h156fa:	data_out=16'h80a5;
17'h156fb:	data_out=16'ha00;
17'h156fc:	data_out=16'h9f3;
17'h156fd:	data_out=16'h89e4;
17'h156fe:	data_out=16'h85e3;
17'h156ff:	data_out=16'h8a00;
17'h15700:	data_out=16'h9ed;
17'h15701:	data_out=16'h9f0;
17'h15702:	data_out=16'h9f9;
17'h15703:	data_out=16'h8a00;
17'h15704:	data_out=16'h8a00;
17'h15705:	data_out=16'h89f9;
17'h15706:	data_out=16'h8a00;
17'h15707:	data_out=16'h87a8;
17'h15708:	data_out=16'h97a;
17'h15709:	data_out=16'h89dc;
17'h1570a:	data_out=16'h393;
17'h1570b:	data_out=16'h89f6;
17'h1570c:	data_out=16'h8a00;
17'h1570d:	data_out=16'h89f4;
17'h1570e:	data_out=16'ha00;
17'h1570f:	data_out=16'h9ed;
17'h15710:	data_out=16'h8a00;
17'h15711:	data_out=16'h62a;
17'h15712:	data_out=16'ha00;
17'h15713:	data_out=16'h8a00;
17'h15714:	data_out=16'h8887;
17'h15715:	data_out=16'h89fe;
17'h15716:	data_out=16'h8a00;
17'h15717:	data_out=16'h85f7;
17'h15718:	data_out=16'ha00;
17'h15719:	data_out=16'h990;
17'h1571a:	data_out=16'h89fc;
17'h1571b:	data_out=16'h96e;
17'h1571c:	data_out=16'h6f2;
17'h1571d:	data_out=16'h9d6;
17'h1571e:	data_out=16'h29e;
17'h1571f:	data_out=16'h8910;
17'h15720:	data_out=16'h8998;
17'h15721:	data_out=16'ha00;
17'h15722:	data_out=16'h89d7;
17'h15723:	data_out=16'h8a00;
17'h15724:	data_out=16'h8a00;
17'h15725:	data_out=16'h89cc;
17'h15726:	data_out=16'h695;
17'h15727:	data_out=16'h923;
17'h15728:	data_out=16'ha00;
17'h15729:	data_out=16'ha00;
17'h1572a:	data_out=16'h9f8;
17'h1572b:	data_out=16'h8a00;
17'h1572c:	data_out=16'h8a00;
17'h1572d:	data_out=16'ha00;
17'h1572e:	data_out=16'ha00;
17'h1572f:	data_out=16'h16e;
17'h15730:	data_out=16'h94e;
17'h15731:	data_out=16'h807d;
17'h15732:	data_out=16'h8073;
17'h15733:	data_out=16'h812a;
17'h15734:	data_out=16'h9e8;
17'h15735:	data_out=16'h2d;
17'h15736:	data_out=16'h9b8;
17'h15737:	data_out=16'ha00;
17'h15738:	data_out=16'h7cc;
17'h15739:	data_out=16'h8189;
17'h1573a:	data_out=16'h89d3;
17'h1573b:	data_out=16'h8a00;
17'h1573c:	data_out=16'h9a1;
17'h1573d:	data_out=16'h89c2;
17'h1573e:	data_out=16'ha00;
17'h1573f:	data_out=16'h89f9;
17'h15740:	data_out=16'h8a00;
17'h15741:	data_out=16'h9b7;
17'h15742:	data_out=16'h8a00;
17'h15743:	data_out=16'h830a;
17'h15744:	data_out=16'h84cf;
17'h15745:	data_out=16'h89ff;
17'h15746:	data_out=16'h9be;
17'h15747:	data_out=16'h8992;
17'h15748:	data_out=16'h89e7;
17'h15749:	data_out=16'h89eb;
17'h1574a:	data_out=16'h77f;
17'h1574b:	data_out=16'h8a00;
17'h1574c:	data_out=16'h89a5;
17'h1574d:	data_out=16'h89e0;
17'h1574e:	data_out=16'ha00;
17'h1574f:	data_out=16'h89cd;
17'h15750:	data_out=16'h8a00;
17'h15751:	data_out=16'h462;
17'h15752:	data_out=16'h8a00;
17'h15753:	data_out=16'h983;
17'h15754:	data_out=16'h9b1;
17'h15755:	data_out=16'h23a;
17'h15756:	data_out=16'h24e;
17'h15757:	data_out=16'h1a3;
17'h15758:	data_out=16'h98d;
17'h15759:	data_out=16'h89e9;
17'h1575a:	data_out=16'h9e0;
17'h1575b:	data_out=16'h54;
17'h1575c:	data_out=16'h9ac;
17'h1575d:	data_out=16'h742;
17'h1575e:	data_out=16'h894c;
17'h1575f:	data_out=16'h9fe;
17'h15760:	data_out=16'h92d;
17'h15761:	data_out=16'h81f;
17'h15762:	data_out=16'h843a;
17'h15763:	data_out=16'h218;
17'h15764:	data_out=16'h87b6;
17'h15765:	data_out=16'h8a00;
17'h15766:	data_out=16'h89fa;
17'h15767:	data_out=16'ha00;
17'h15768:	data_out=16'ha00;
17'h15769:	data_out=16'h891;
17'h1576a:	data_out=16'ha00;
17'h1576b:	data_out=16'h8a00;
17'h1576c:	data_out=16'h9fd;
17'h1576d:	data_out=16'h188;
17'h1576e:	data_out=16'ha00;
17'h1576f:	data_out=16'h8a00;
17'h15770:	data_out=16'ha00;
17'h15771:	data_out=16'h9ff;
17'h15772:	data_out=16'h89c2;
17'h15773:	data_out=16'h2f0;
17'h15774:	data_out=16'h915;
17'h15775:	data_out=16'h574;
17'h15776:	data_out=16'h9ba;
17'h15777:	data_out=16'h89fd;
17'h15778:	data_out=16'h176;
17'h15779:	data_out=16'h9fd;
17'h1577a:	data_out=16'h8053;
17'h1577b:	data_out=16'ha00;
17'h1577c:	data_out=16'ha00;
17'h1577d:	data_out=16'h89a2;
17'h1577e:	data_out=16'h881f;
17'h1577f:	data_out=16'h8a00;
17'h15780:	data_out=16'h7bf;
17'h15781:	data_out=16'h9fa;
17'h15782:	data_out=16'h9c7;
17'h15783:	data_out=16'h8a00;
17'h15784:	data_out=16'h8a00;
17'h15785:	data_out=16'h86d5;
17'h15786:	data_out=16'h8a00;
17'h15787:	data_out=16'h8a00;
17'h15788:	data_out=16'h96b;
17'h15789:	data_out=16'h8a00;
17'h1578a:	data_out=16'h686;
17'h1578b:	data_out=16'h89fc;
17'h1578c:	data_out=16'h8a00;
17'h1578d:	data_out=16'h89fe;
17'h1578e:	data_out=16'ha00;
17'h1578f:	data_out=16'h9dc;
17'h15790:	data_out=16'h8a00;
17'h15791:	data_out=16'h8a00;
17'h15792:	data_out=16'ha00;
17'h15793:	data_out=16'h8a00;
17'h15794:	data_out=16'h318;
17'h15795:	data_out=16'h89ea;
17'h15796:	data_out=16'h89e6;
17'h15797:	data_out=16'h58e;
17'h15798:	data_out=16'h9ff;
17'h15799:	data_out=16'h7e;
17'h1579a:	data_out=16'h89fc;
17'h1579b:	data_out=16'h943;
17'h1579c:	data_out=16'h916;
17'h1579d:	data_out=16'h9ef;
17'h1579e:	data_out=16'h9f6;
17'h1579f:	data_out=16'h882e;
17'h157a0:	data_out=16'h8781;
17'h157a1:	data_out=16'ha00;
17'h157a2:	data_out=16'h89dc;
17'h157a3:	data_out=16'h8a00;
17'h157a4:	data_out=16'h8a00;
17'h157a5:	data_out=16'h8a00;
17'h157a6:	data_out=16'h74e;
17'h157a7:	data_out=16'h508;
17'h157a8:	data_out=16'ha00;
17'h157a9:	data_out=16'ha00;
17'h157aa:	data_out=16'h9d7;
17'h157ab:	data_out=16'h8a00;
17'h157ac:	data_out=16'h89d3;
17'h157ad:	data_out=16'ha00;
17'h157ae:	data_out=16'ha00;
17'h157af:	data_out=16'h8131;
17'h157b0:	data_out=16'h8e5;
17'h157b1:	data_out=16'h188;
17'h157b2:	data_out=16'h8a00;
17'h157b3:	data_out=16'h6c6;
17'h157b4:	data_out=16'h9fb;
17'h157b5:	data_out=16'h89fe;
17'h157b6:	data_out=16'h9b9;
17'h157b7:	data_out=16'h9e5;
17'h157b8:	data_out=16'h8fb;
17'h157b9:	data_out=16'h663;
17'h157ba:	data_out=16'h89fc;
17'h157bb:	data_out=16'h8a00;
17'h157bc:	data_out=16'h9aa;
17'h157bd:	data_out=16'h87db;
17'h157be:	data_out=16'ha00;
17'h157bf:	data_out=16'h86b5;
17'h157c0:	data_out=16'h8a00;
17'h157c1:	data_out=16'h9c0;
17'h157c2:	data_out=16'h8a00;
17'h157c3:	data_out=16'h464;
17'h157c4:	data_out=16'h8a00;
17'h157c5:	data_out=16'h89e8;
17'h157c6:	data_out=16'h9b6;
17'h157c7:	data_out=16'h89bb;
17'h157c8:	data_out=16'h89f0;
17'h157c9:	data_out=16'h8a00;
17'h157ca:	data_out=16'h89fe;
17'h157cb:	data_out=16'h8a00;
17'h157cc:	data_out=16'h89da;
17'h157cd:	data_out=16'h89e4;
17'h157ce:	data_out=16'h9f3;
17'h157cf:	data_out=16'h89f9;
17'h157d0:	data_out=16'h8a00;
17'h157d1:	data_out=16'h9f3;
17'h157d2:	data_out=16'h8a00;
17'h157d3:	data_out=16'h968;
17'h157d4:	data_out=16'h6ec;
17'h157d5:	data_out=16'h745;
17'h157d6:	data_out=16'h281;
17'h157d7:	data_out=16'h8025;
17'h157d8:	data_out=16'h9ba;
17'h157d9:	data_out=16'h89f8;
17'h157da:	data_out=16'h9ed;
17'h157db:	data_out=16'h8469;
17'h157dc:	data_out=16'h9ad;
17'h157dd:	data_out=16'h953;
17'h157de:	data_out=16'h8836;
17'h157df:	data_out=16'h9ff;
17'h157e0:	data_out=16'h820;
17'h157e1:	data_out=16'h895;
17'h157e2:	data_out=16'h1b7;
17'h157e3:	data_out=16'h839;
17'h157e4:	data_out=16'h88f5;
17'h157e5:	data_out=16'h8a00;
17'h157e6:	data_out=16'h8825;
17'h157e7:	data_out=16'ha00;
17'h157e8:	data_out=16'ha00;
17'h157e9:	data_out=16'h60b;
17'h157ea:	data_out=16'ha00;
17'h157eb:	data_out=16'h89cc;
17'h157ec:	data_out=16'h9ff;
17'h157ed:	data_out=16'h7e7;
17'h157ee:	data_out=16'ha00;
17'h157ef:	data_out=16'h8a00;
17'h157f0:	data_out=16'ha00;
17'h157f1:	data_out=16'h9fe;
17'h157f2:	data_out=16'h303;
17'h157f3:	data_out=16'h830;
17'h157f4:	data_out=16'h939;
17'h157f5:	data_out=16'h73f;
17'h157f6:	data_out=16'h95b;
17'h157f7:	data_out=16'h8a00;
17'h157f8:	data_out=16'h403;
17'h157f9:	data_out=16'h9f5;
17'h157fa:	data_out=16'h734;
17'h157fb:	data_out=16'ha00;
17'h157fc:	data_out=16'ha00;
17'h157fd:	data_out=16'h8908;
17'h157fe:	data_out=16'h88ee;
17'h157ff:	data_out=16'h865d;
17'h15800:	data_out=16'h84e2;
17'h15801:	data_out=16'h9fe;
17'h15802:	data_out=16'h9c0;
17'h15803:	data_out=16'h89fd;
17'h15804:	data_out=16'h89f8;
17'h15805:	data_out=16'h84ed;
17'h15806:	data_out=16'h89f4;
17'h15807:	data_out=16'h8a00;
17'h15808:	data_out=16'h841;
17'h15809:	data_out=16'h89fd;
17'h1580a:	data_out=16'h90b;
17'h1580b:	data_out=16'h89fa;
17'h1580c:	data_out=16'h8a00;
17'h1580d:	data_out=16'h89fb;
17'h1580e:	data_out=16'ha00;
17'h1580f:	data_out=16'h9dd;
17'h15810:	data_out=16'h89fe;
17'h15811:	data_out=16'h8a00;
17'h15812:	data_out=16'h9ff;
17'h15813:	data_out=16'h8a00;
17'h15814:	data_out=16'h7ab;
17'h15815:	data_out=16'h89ef;
17'h15816:	data_out=16'h89fb;
17'h15817:	data_out=16'h91b;
17'h15818:	data_out=16'h9fd;
17'h15819:	data_out=16'h9af;
17'h1581a:	data_out=16'h87a3;
17'h1581b:	data_out=16'h91c;
17'h1581c:	data_out=16'h5e9;
17'h1581d:	data_out=16'h2f6;
17'h1581e:	data_out=16'h9f8;
17'h1581f:	data_out=16'h8291;
17'h15820:	data_out=16'h86e8;
17'h15821:	data_out=16'ha00;
17'h15822:	data_out=16'h65a;
17'h15823:	data_out=16'h8a00;
17'h15824:	data_out=16'h8a00;
17'h15825:	data_out=16'h89fc;
17'h15826:	data_out=16'hb4;
17'h15827:	data_out=16'h8700;
17'h15828:	data_out=16'ha00;
17'h15829:	data_out=16'ha00;
17'h1582a:	data_out=16'h9d7;
17'h1582b:	data_out=16'h8a00;
17'h1582c:	data_out=16'h89e5;
17'h1582d:	data_out=16'ha00;
17'h1582e:	data_out=16'h9fe;
17'h1582f:	data_out=16'h874c;
17'h15830:	data_out=16'h968;
17'h15831:	data_out=16'h85c6;
17'h15832:	data_out=16'h8477;
17'h15833:	data_out=16'h9fb;
17'h15834:	data_out=16'h6dc;
17'h15835:	data_out=16'h886f;
17'h15836:	data_out=16'h3ef;
17'h15837:	data_out=16'h9eb;
17'h15838:	data_out=16'h9fe;
17'h15839:	data_out=16'h96f;
17'h1583a:	data_out=16'h89ff;
17'h1583b:	data_out=16'h8a00;
17'h1583c:	data_out=16'h9f2;
17'h1583d:	data_out=16'h8646;
17'h1583e:	data_out=16'ha00;
17'h1583f:	data_out=16'h84e8;
17'h15840:	data_out=16'h89fb;
17'h15841:	data_out=16'h646;
17'h15842:	data_out=16'h8a00;
17'h15843:	data_out=16'h836c;
17'h15844:	data_out=16'h89ea;
17'h15845:	data_out=16'h89ef;
17'h15846:	data_out=16'h9ea;
17'h15847:	data_out=16'h897d;
17'h15848:	data_out=16'h84a7;
17'h15849:	data_out=16'h89fe;
17'h1584a:	data_out=16'h89d2;
17'h1584b:	data_out=16'h8a00;
17'h1584c:	data_out=16'h89f7;
17'h1584d:	data_out=16'h9f8;
17'h1584e:	data_out=16'h9fb;
17'h1584f:	data_out=16'h89fd;
17'h15850:	data_out=16'h89f0;
17'h15851:	data_out=16'h9e6;
17'h15852:	data_out=16'h8a00;
17'h15853:	data_out=16'h9de;
17'h15854:	data_out=16'h8320;
17'h15855:	data_out=16'h6e0;
17'h15856:	data_out=16'h493;
17'h15857:	data_out=16'h635;
17'h15858:	data_out=16'h9c3;
17'h15859:	data_out=16'h88da;
17'h1585a:	data_out=16'h9fe;
17'h1585b:	data_out=16'h8962;
17'h1585c:	data_out=16'h9e3;
17'h1585d:	data_out=16'h684;
17'h1585e:	data_out=16'h8878;
17'h1585f:	data_out=16'h9ff;
17'h15860:	data_out=16'h757;
17'h15861:	data_out=16'h9ec;
17'h15862:	data_out=16'h1f6;
17'h15863:	data_out=16'h9ff;
17'h15864:	data_out=16'h89cb;
17'h15865:	data_out=16'h89fb;
17'h15866:	data_out=16'h9e3;
17'h15867:	data_out=16'ha00;
17'h15868:	data_out=16'ha00;
17'h15869:	data_out=16'h3be;
17'h1586a:	data_out=16'ha00;
17'h1586b:	data_out=16'h8990;
17'h1586c:	data_out=16'h49a;
17'h1586d:	data_out=16'h9ff;
17'h1586e:	data_out=16'ha00;
17'h1586f:	data_out=16'h89fb;
17'h15870:	data_out=16'ha00;
17'h15871:	data_out=16'h9f2;
17'h15872:	data_out=16'h698;
17'h15873:	data_out=16'h9eb;
17'h15874:	data_out=16'h94c;
17'h15875:	data_out=16'h96f;
17'h15876:	data_out=16'h9d8;
17'h15877:	data_out=16'h89ff;
17'h15878:	data_out=16'h83a1;
17'h15879:	data_out=16'h9fa;
17'h1587a:	data_out=16'h9f2;
17'h1587b:	data_out=16'ha00;
17'h1587c:	data_out=16'ha00;
17'h1587d:	data_out=16'h85fe;
17'h1587e:	data_out=16'h89e0;
17'h1587f:	data_out=16'h197;
17'h15880:	data_out=16'h87f3;
17'h15881:	data_out=16'h48;
17'h15882:	data_out=16'h9ca;
17'h15883:	data_out=16'h8840;
17'h15884:	data_out=16'h878a;
17'h15885:	data_out=16'h8545;
17'h15886:	data_out=16'h8977;
17'h15887:	data_out=16'h8a00;
17'h15888:	data_out=16'h33a;
17'h15889:	data_out=16'h89fe;
17'h1588a:	data_out=16'h838e;
17'h1588b:	data_out=16'h6a2;
17'h1588c:	data_out=16'h8a00;
17'h1588d:	data_out=16'h86b6;
17'h1588e:	data_out=16'h9ff;
17'h1588f:	data_out=16'h837;
17'h15890:	data_out=16'h89e3;
17'h15891:	data_out=16'h89fa;
17'h15892:	data_out=16'h9fb;
17'h15893:	data_out=16'h89f5;
17'h15894:	data_out=16'h9f1;
17'h15895:	data_out=16'h88db;
17'h15896:	data_out=16'h89db;
17'h15897:	data_out=16'h9e7;
17'h15898:	data_out=16'h9fc;
17'h15899:	data_out=16'h549;
17'h1589a:	data_out=16'h869b;
17'h1589b:	data_out=16'h9f2;
17'h1589c:	data_out=16'h5e3;
17'h1589d:	data_out=16'h8852;
17'h1589e:	data_out=16'h9ff;
17'h1589f:	data_out=16'h3e6;
17'h158a0:	data_out=16'h83dc;
17'h158a1:	data_out=16'h9ff;
17'h158a2:	data_out=16'h9b4;
17'h158a3:	data_out=16'h8a00;
17'h158a4:	data_out=16'h8a00;
17'h158a5:	data_out=16'h89fe;
17'h158a6:	data_out=16'h915;
17'h158a7:	data_out=16'h887b;
17'h158a8:	data_out=16'h9ff;
17'h158a9:	data_out=16'ha00;
17'h158aa:	data_out=16'h87b3;
17'h158ab:	data_out=16'h150;
17'h158ac:	data_out=16'h89c3;
17'h158ad:	data_out=16'ha00;
17'h158ae:	data_out=16'h9dc;
17'h158af:	data_out=16'h86c5;
17'h158b0:	data_out=16'h20c;
17'h158b1:	data_out=16'h89b9;
17'h158b2:	data_out=16'h898d;
17'h158b3:	data_out=16'ha00;
17'h158b4:	data_out=16'h8569;
17'h158b5:	data_out=16'h8599;
17'h158b6:	data_out=16'h863d;
17'h158b7:	data_out=16'h9ea;
17'h158b8:	data_out=16'h869b;
17'h158b9:	data_out=16'ha00;
17'h158ba:	data_out=16'h89cb;
17'h158bb:	data_out=16'h89fe;
17'h158bc:	data_out=16'ha00;
17'h158bd:	data_out=16'h81fb;
17'h158be:	data_out=16'h9ff;
17'h158bf:	data_out=16'h8534;
17'h158c0:	data_out=16'h89f1;
17'h158c1:	data_out=16'h883;
17'h158c2:	data_out=16'h89ff;
17'h158c3:	data_out=16'h82f1;
17'h158c4:	data_out=16'h85be;
17'h158c5:	data_out=16'h88e8;
17'h158c6:	data_out=16'ha00;
17'h158c7:	data_out=16'h88c2;
17'h158c8:	data_out=16'h8426;
17'h158c9:	data_out=16'h89f9;
17'h158ca:	data_out=16'h88f8;
17'h158cb:	data_out=16'h89fe;
17'h158cc:	data_out=16'h89ff;
17'h158cd:	data_out=16'ha00;
17'h158ce:	data_out=16'h9ff;
17'h158cf:	data_out=16'h89ff;
17'h158d0:	data_out=16'h8714;
17'h158d1:	data_out=16'h9ef;
17'h158d2:	data_out=16'h8a00;
17'h158d3:	data_out=16'h58;
17'h158d4:	data_out=16'h83b3;
17'h158d5:	data_out=16'h98f;
17'h158d6:	data_out=16'h92c;
17'h158d7:	data_out=16'h9d8;
17'h158d8:	data_out=16'h9fb;
17'h158d9:	data_out=16'h85f0;
17'h158da:	data_out=16'ha00;
17'h158db:	data_out=16'h8597;
17'h158dc:	data_out=16'h75a;
17'h158dd:	data_out=16'h86d7;
17'h158de:	data_out=16'h87e5;
17'h158df:	data_out=16'h518;
17'h158e0:	data_out=16'hae;
17'h158e1:	data_out=16'h73d;
17'h158e2:	data_out=16'h60e;
17'h158e3:	data_out=16'ha00;
17'h158e4:	data_out=16'h89c9;
17'h158e5:	data_out=16'h89ef;
17'h158e6:	data_out=16'h9fa;
17'h158e7:	data_out=16'ha00;
17'h158e8:	data_out=16'h9ff;
17'h158e9:	data_out=16'h6b5;
17'h158ea:	data_out=16'ha00;
17'h158eb:	data_out=16'h874e;
17'h158ec:	data_out=16'h8500;
17'h158ed:	data_out=16'ha00;
17'h158ee:	data_out=16'ha00;
17'h158ef:	data_out=16'h89fa;
17'h158f0:	data_out=16'h9ff;
17'h158f1:	data_out=16'h7db;
17'h158f2:	data_out=16'h8625;
17'h158f3:	data_out=16'h765;
17'h158f4:	data_out=16'h192;
17'h158f5:	data_out=16'h986;
17'h158f6:	data_out=16'h9f3;
17'h158f7:	data_out=16'h89fd;
17'h158f8:	data_out=16'h89f8;
17'h158f9:	data_out=16'ha00;
17'h158fa:	data_out=16'h9ff;
17'h158fb:	data_out=16'h9ff;
17'h158fc:	data_out=16'h9fc;
17'h158fd:	data_out=16'hb8;
17'h158fe:	data_out=16'h89ee;
17'h158ff:	data_out=16'h9ba;
17'h15900:	data_out=16'h88c5;
17'h15901:	data_out=16'h87cf;
17'h15902:	data_out=16'h9e4;
17'h15903:	data_out=16'h8837;
17'h15904:	data_out=16'h8518;
17'h15905:	data_out=16'h873b;
17'h15906:	data_out=16'h89fd;
17'h15907:	data_out=16'h8a00;
17'h15908:	data_out=16'h8993;
17'h15909:	data_out=16'h89fd;
17'h1590a:	data_out=16'h8253;
17'h1590b:	data_out=16'h897b;
17'h1590c:	data_out=16'h89ff;
17'h1590d:	data_out=16'h84ae;
17'h1590e:	data_out=16'ha00;
17'h1590f:	data_out=16'h84a9;
17'h15910:	data_out=16'h89f3;
17'h15911:	data_out=16'h89f7;
17'h15912:	data_out=16'h597;
17'h15913:	data_out=16'h88e3;
17'h15914:	data_out=16'h9c8;
17'h15915:	data_out=16'h83fe;
17'h15916:	data_out=16'h89f1;
17'h15917:	data_out=16'h904;
17'h15918:	data_out=16'h9fd;
17'h15919:	data_out=16'h8363;
17'h1591a:	data_out=16'h86ea;
17'h1591b:	data_out=16'h8035;
17'h1591c:	data_out=16'hdb;
17'h1591d:	data_out=16'h8a00;
17'h1591e:	data_out=16'h9f2;
17'h1591f:	data_out=16'hbf;
17'h15920:	data_out=16'h888d;
17'h15921:	data_out=16'ha00;
17'h15922:	data_out=16'ha00;
17'h15923:	data_out=16'h87a9;
17'h15924:	data_out=16'h87af;
17'h15925:	data_out=16'h85fc;
17'h15926:	data_out=16'h9fb;
17'h15927:	data_out=16'h89df;
17'h15928:	data_out=16'ha00;
17'h15929:	data_out=16'h9fe;
17'h1592a:	data_out=16'h89c1;
17'h1592b:	data_out=16'h87ff;
17'h1592c:	data_out=16'h89ef;
17'h1592d:	data_out=16'h9f4;
17'h1592e:	data_out=16'h8113;
17'h1592f:	data_out=16'h89c1;
17'h15930:	data_out=16'hf7;
17'h15931:	data_out=16'h89f6;
17'h15932:	data_out=16'h88b3;
17'h15933:	data_out=16'h9e1;
17'h15934:	data_out=16'h89e0;
17'h15935:	data_out=16'h86d4;
17'h15936:	data_out=16'h8989;
17'h15937:	data_out=16'h9ef;
17'h15938:	data_out=16'h89ca;
17'h15939:	data_out=16'ha00;
17'h1593a:	data_out=16'h89d0;
17'h1593b:	data_out=16'h89ff;
17'h1593c:	data_out=16'ha00;
17'h1593d:	data_out=16'h835c;
17'h1593e:	data_out=16'ha00;
17'h1593f:	data_out=16'h870c;
17'h15940:	data_out=16'h8840;
17'h15941:	data_out=16'h86fc;
17'h15942:	data_out=16'h89fe;
17'h15943:	data_out=16'h860a;
17'h15944:	data_out=16'h8886;
17'h15945:	data_out=16'h84d5;
17'h15946:	data_out=16'ha00;
17'h15947:	data_out=16'h8987;
17'h15948:	data_out=16'h89b1;
17'h15949:	data_out=16'h83f3;
17'h1594a:	data_out=16'h89fd;
17'h1594b:	data_out=16'h89fd;
17'h1594c:	data_out=16'h8985;
17'h1594d:	data_out=16'h9fc;
17'h1594e:	data_out=16'h88ea;
17'h1594f:	data_out=16'h89f4;
17'h15950:	data_out=16'h861e;
17'h15951:	data_out=16'h9ea;
17'h15952:	data_out=16'h8184;
17'h15953:	data_out=16'h8977;
17'h15954:	data_out=16'h88c2;
17'h15955:	data_out=16'h848;
17'h15956:	data_out=16'h9e6;
17'h15957:	data_out=16'h9ff;
17'h15958:	data_out=16'h9f7;
17'h15959:	data_out=16'h8248;
17'h1595a:	data_out=16'ha00;
17'h1595b:	data_out=16'h869f;
17'h1595c:	data_out=16'h8738;
17'h1595d:	data_out=16'h8943;
17'h1595e:	data_out=16'h89dc;
17'h1595f:	data_out=16'h89b1;
17'h15960:	data_out=16'h977;
17'h15961:	data_out=16'h212;
17'h15962:	data_out=16'h81;
17'h15963:	data_out=16'h770;
17'h15964:	data_out=16'h89df;
17'h15965:	data_out=16'h8a00;
17'h15966:	data_out=16'h86e8;
17'h15967:	data_out=16'h9fb;
17'h15968:	data_out=16'ha00;
17'h15969:	data_out=16'h841a;
17'h1596a:	data_out=16'ha00;
17'h1596b:	data_out=16'h884d;
17'h1596c:	data_out=16'h8809;
17'h1596d:	data_out=16'h7b4;
17'h1596e:	data_out=16'ha00;
17'h1596f:	data_out=16'h89ff;
17'h15970:	data_out=16'ha00;
17'h15971:	data_out=16'h8746;
17'h15972:	data_out=16'h1f;
17'h15973:	data_out=16'h445;
17'h15974:	data_out=16'heb;
17'h15975:	data_out=16'h9a8;
17'h15976:	data_out=16'h8150;
17'h15977:	data_out=16'h89f9;
17'h15978:	data_out=16'h89fd;
17'h15979:	data_out=16'h8265;
17'h1597a:	data_out=16'h992;
17'h1597b:	data_out=16'ha00;
17'h1597c:	data_out=16'h6b8;
17'h1597d:	data_out=16'h858b;
17'h1597e:	data_out=16'h89eb;
17'h1597f:	data_out=16'ha00;
17'h15980:	data_out=16'h89c5;
17'h15981:	data_out=16'h8a00;
17'h15982:	data_out=16'h9f8;
17'h15983:	data_out=16'h86f8;
17'h15984:	data_out=16'h882d;
17'h15985:	data_out=16'h899f;
17'h15986:	data_out=16'h8a00;
17'h15987:	data_out=16'h89ff;
17'h15988:	data_out=16'h89d6;
17'h15989:	data_out=16'h89ff;
17'h1598a:	data_out=16'h87ca;
17'h1598b:	data_out=16'h89e0;
17'h1598c:	data_out=16'h89ff;
17'h1598d:	data_out=16'h14;
17'h1598e:	data_out=16'ha00;
17'h1598f:	data_out=16'h89fc;
17'h15990:	data_out=16'h89f2;
17'h15991:	data_out=16'h8a00;
17'h15992:	data_out=16'h100;
17'h15993:	data_out=16'h8442;
17'h15994:	data_out=16'h9dc;
17'h15995:	data_out=16'h8940;
17'h15996:	data_out=16'h89fc;
17'h15997:	data_out=16'h88a;
17'h15998:	data_out=16'h9b6;
17'h15999:	data_out=16'h8770;
17'h1599a:	data_out=16'h89c3;
17'h1599b:	data_out=16'h8178;
17'h1599c:	data_out=16'h80c3;
17'h1599d:	data_out=16'h8a00;
17'h1599e:	data_out=16'h47a;
17'h1599f:	data_out=16'h2f1;
17'h159a0:	data_out=16'h89f6;
17'h159a1:	data_out=16'ha00;
17'h159a2:	data_out=16'ha00;
17'h159a3:	data_out=16'h86a0;
17'h159a4:	data_out=16'h86a7;
17'h159a5:	data_out=16'h8006;
17'h159a6:	data_out=16'ha00;
17'h159a7:	data_out=16'h8a00;
17'h159a8:	data_out=16'ha00;
17'h159a9:	data_out=16'ha00;
17'h159aa:	data_out=16'h89fd;
17'h159ab:	data_out=16'h88a3;
17'h159ac:	data_out=16'h89fb;
17'h159ad:	data_out=16'h691;
17'h159ae:	data_out=16'h8a00;
17'h159af:	data_out=16'h89ff;
17'h159b0:	data_out=16'h82fb;
17'h159b1:	data_out=16'h8a00;
17'h159b2:	data_out=16'h8a00;
17'h159b3:	data_out=16'h904;
17'h159b4:	data_out=16'h8a00;
17'h159b5:	data_out=16'h89f3;
17'h159b6:	data_out=16'h89fd;
17'h159b7:	data_out=16'h9fc;
17'h159b8:	data_out=16'h8a00;
17'h159b9:	data_out=16'h996;
17'h159ba:	data_out=16'h89fb;
17'h159bb:	data_out=16'h89ff;
17'h159bc:	data_out=16'ha00;
17'h159bd:	data_out=16'h889e;
17'h159be:	data_out=16'ha00;
17'h159bf:	data_out=16'h8981;
17'h159c0:	data_out=16'h89fe;
17'h159c1:	data_out=16'h87ea;
17'h159c2:	data_out=16'h89ff;
17'h159c3:	data_out=16'h85;
17'h159c4:	data_out=16'h89f1;
17'h159c5:	data_out=16'h8953;
17'h159c6:	data_out=16'ha00;
17'h159c7:	data_out=16'h89f1;
17'h159c8:	data_out=16'h89fe;
17'h159c9:	data_out=16'h801a;
17'h159ca:	data_out=16'h89ff;
17'h159cb:	data_out=16'h89ff;
17'h159cc:	data_out=16'h8996;
17'h159cd:	data_out=16'h9fe;
17'h159ce:	data_out=16'h8945;
17'h159cf:	data_out=16'h89f7;
17'h159d0:	data_out=16'h861d;
17'h159d1:	data_out=16'ha00;
17'h159d2:	data_out=16'h836e;
17'h159d3:	data_out=16'h89ff;
17'h159d4:	data_out=16'h89f5;
17'h159d5:	data_out=16'h921;
17'h159d6:	data_out=16'ha00;
17'h159d7:	data_out=16'ha00;
17'h159d8:	data_out=16'ha00;
17'h159d9:	data_out=16'h87a8;
17'h159da:	data_out=16'ha00;
17'h159db:	data_out=16'h8970;
17'h159dc:	data_out=16'h88b2;
17'h159dd:	data_out=16'h89fe;
17'h159de:	data_out=16'h89ff;
17'h159df:	data_out=16'h89fb;
17'h159e0:	data_out=16'h188;
17'h159e1:	data_out=16'h863f;
17'h159e2:	data_out=16'h8f;
17'h159e3:	data_out=16'h637;
17'h159e4:	data_out=16'h89f8;
17'h159e5:	data_out=16'h8a00;
17'h159e6:	data_out=16'h89ee;
17'h159e7:	data_out=16'h493;
17'h159e8:	data_out=16'ha00;
17'h159e9:	data_out=16'h5a;
17'h159ea:	data_out=16'ha00;
17'h159eb:	data_out=16'h89fe;
17'h159ec:	data_out=16'h89d5;
17'h159ed:	data_out=16'h684;
17'h159ee:	data_out=16'ha00;
17'h159ef:	data_out=16'h8a00;
17'h159f0:	data_out=16'ha00;
17'h159f1:	data_out=16'h89fd;
17'h159f2:	data_out=16'h886e;
17'h159f3:	data_out=16'h870d;
17'h159f4:	data_out=16'h8304;
17'h159f5:	data_out=16'h9de;
17'h159f6:	data_out=16'h89fc;
17'h159f7:	data_out=16'h89fd;
17'h159f8:	data_out=16'h864f;
17'h159f9:	data_out=16'h85bf;
17'h159fa:	data_out=16'h865;
17'h159fb:	data_out=16'ha00;
17'h159fc:	data_out=16'h844f;
17'h159fd:	data_out=16'h8962;
17'h159fe:	data_out=16'h85f3;
17'h159ff:	data_out=16'h679;
17'h15a00:	data_out=16'h89f9;
17'h15a01:	data_out=16'h8a00;
17'h15a02:	data_out=16'h9e0;
17'h15a03:	data_out=16'h214;
17'h15a04:	data_out=16'h891c;
17'h15a05:	data_out=16'h8a00;
17'h15a06:	data_out=16'h57a;
17'h15a07:	data_out=16'h8a00;
17'h15a08:	data_out=16'h8361;
17'h15a09:	data_out=16'h4f2;
17'h15a0a:	data_out=16'h89fb;
17'h15a0b:	data_out=16'h7d5;
17'h15a0c:	data_out=16'h8a00;
17'h15a0d:	data_out=16'h4c8;
17'h15a0e:	data_out=16'ha00;
17'h15a0f:	data_out=16'h89ff;
17'h15a10:	data_out=16'h81da;
17'h15a11:	data_out=16'h8a00;
17'h15a12:	data_out=16'h89f8;
17'h15a13:	data_out=16'h1ba;
17'h15a14:	data_out=16'h9fd;
17'h15a15:	data_out=16'h8763;
17'h15a16:	data_out=16'h89fc;
17'h15a17:	data_out=16'h9ec;
17'h15a18:	data_out=16'h885;
17'h15a19:	data_out=16'h8862;
17'h15a1a:	data_out=16'h8a00;
17'h15a1b:	data_out=16'h45;
17'h15a1c:	data_out=16'h809a;
17'h15a1d:	data_out=16'h8a00;
17'h15a1e:	data_out=16'h6e9;
17'h15a1f:	data_out=16'h835;
17'h15a20:	data_out=16'h8a00;
17'h15a21:	data_out=16'ha00;
17'h15a22:	data_out=16'ha00;
17'h15a23:	data_out=16'h8816;
17'h15a24:	data_out=16'h8817;
17'h15a25:	data_out=16'h725;
17'h15a26:	data_out=16'ha00;
17'h15a27:	data_out=16'h8a00;
17'h15a28:	data_out=16'ha00;
17'h15a29:	data_out=16'h19c;
17'h15a2a:	data_out=16'h89ff;
17'h15a2b:	data_out=16'h2f3;
17'h15a2c:	data_out=16'h89fc;
17'h15a2d:	data_out=16'h801b;
17'h15a2e:	data_out=16'h8a00;
17'h15a2f:	data_out=16'h8a00;
17'h15a30:	data_out=16'h872a;
17'h15a31:	data_out=16'h8a00;
17'h15a32:	data_out=16'h8a00;
17'h15a33:	data_out=16'h9fe;
17'h15a34:	data_out=16'h8a00;
17'h15a35:	data_out=16'h89f5;
17'h15a36:	data_out=16'h89ff;
17'h15a37:	data_out=16'h9cc;
17'h15a38:	data_out=16'h8a00;
17'h15a39:	data_out=16'ha00;
17'h15a3a:	data_out=16'h89f1;
17'h15a3b:	data_out=16'h89fc;
17'h15a3c:	data_out=16'ha00;
17'h15a3d:	data_out=16'h89c3;
17'h15a3e:	data_out=16'ha00;
17'h15a3f:	data_out=16'h89ff;
17'h15a40:	data_out=16'h89fc;
17'h15a41:	data_out=16'h80c4;
17'h15a42:	data_out=16'h89fd;
17'h15a43:	data_out=16'h9f5;
17'h15a44:	data_out=16'h89f5;
17'h15a45:	data_out=16'h884a;
17'h15a46:	data_out=16'ha00;
17'h15a47:	data_out=16'h89fe;
17'h15a48:	data_out=16'h8a00;
17'h15a49:	data_out=16'h828;
17'h15a4a:	data_out=16'h8a00;
17'h15a4b:	data_out=16'h89ff;
17'h15a4c:	data_out=16'h89ee;
17'h15a4d:	data_out=16'h9fc;
17'h15a4e:	data_out=16'h89dc;
17'h15a4f:	data_out=16'h89f7;
17'h15a50:	data_out=16'h5f0;
17'h15a51:	data_out=16'ha00;
17'h15a52:	data_out=16'h868a;
17'h15a53:	data_out=16'h8a00;
17'h15a54:	data_out=16'h8a00;
17'h15a55:	data_out=16'ha00;
17'h15a56:	data_out=16'ha00;
17'h15a57:	data_out=16'ha00;
17'h15a58:	data_out=16'ha00;
17'h15a59:	data_out=16'h89f2;
17'h15a5a:	data_out=16'ha00;
17'h15a5b:	data_out=16'h89f2;
17'h15a5c:	data_out=16'h88ec;
17'h15a5d:	data_out=16'h8a00;
17'h15a5e:	data_out=16'h8a00;
17'h15a5f:	data_out=16'h8a00;
17'h15a60:	data_out=16'h897c;
17'h15a61:	data_out=16'h898e;
17'h15a62:	data_out=16'h534;
17'h15a63:	data_out=16'h97b;
17'h15a64:	data_out=16'h8a00;
17'h15a65:	data_out=16'h8a00;
17'h15a66:	data_out=16'h8499;
17'h15a67:	data_out=16'h81ed;
17'h15a68:	data_out=16'ha00;
17'h15a69:	data_out=16'h7d7;
17'h15a6a:	data_out=16'ha00;
17'h15a6b:	data_out=16'h8a00;
17'h15a6c:	data_out=16'h89ff;
17'h15a6d:	data_out=16'h9bb;
17'h15a6e:	data_out=16'ha00;
17'h15a6f:	data_out=16'h8a00;
17'h15a70:	data_out=16'ha00;
17'h15a71:	data_out=16'h89ff;
17'h15a72:	data_out=16'h89fe;
17'h15a73:	data_out=16'h8a00;
17'h15a74:	data_out=16'h8767;
17'h15a75:	data_out=16'h9fb;
17'h15a76:	data_out=16'h12c;
17'h15a77:	data_out=16'h7ce;
17'h15a78:	data_out=16'h9e4;
17'h15a79:	data_out=16'h87dd;
17'h15a7a:	data_out=16'h9f4;
17'h15a7b:	data_out=16'ha00;
17'h15a7c:	data_out=16'h89fb;
17'h15a7d:	data_out=16'h5f2;
17'h15a7e:	data_out=16'ha00;
17'h15a7f:	data_out=16'h8003;
17'h15a80:	data_out=16'h89e9;
17'h15a81:	data_out=16'h8a00;
17'h15a82:	data_out=16'h3aa;
17'h15a83:	data_out=16'h5eb;
17'h15a84:	data_out=16'h88da;
17'h15a85:	data_out=16'h89fd;
17'h15a86:	data_out=16'h917;
17'h15a87:	data_out=16'h8a00;
17'h15a88:	data_out=16'h86ad;
17'h15a89:	data_out=16'h8a4;
17'h15a8a:	data_out=16'h8a00;
17'h15a8b:	data_out=16'h9f1;
17'h15a8c:	data_out=16'h89ff;
17'h15a8d:	data_out=16'h2fc;
17'h15a8e:	data_out=16'h4fc;
17'h15a8f:	data_out=16'h89ff;
17'h15a90:	data_out=16'h9f1;
17'h15a91:	data_out=16'h89fa;
17'h15a92:	data_out=16'h89f4;
17'h15a93:	data_out=16'h4b7;
17'h15a94:	data_out=16'ha00;
17'h15a95:	data_out=16'h82ca;
17'h15a96:	data_out=16'h89f0;
17'h15a97:	data_out=16'h9f7;
17'h15a98:	data_out=16'h489;
17'h15a99:	data_out=16'h8a00;
17'h15a9a:	data_out=16'h89f9;
17'h15a9b:	data_out=16'h8301;
17'h15a9c:	data_out=16'h8291;
17'h15a9d:	data_out=16'h8a00;
17'h15a9e:	data_out=16'h9ff;
17'h15a9f:	data_out=16'h983;
17'h15aa0:	data_out=16'h89da;
17'h15aa1:	data_out=16'h501;
17'h15aa2:	data_out=16'ha00;
17'h15aa3:	data_out=16'h89c1;
17'h15aa4:	data_out=16'h89c2;
17'h15aa5:	data_out=16'h6e8;
17'h15aa6:	data_out=16'h9fe;
17'h15aa7:	data_out=16'h8a00;
17'h15aa8:	data_out=16'h540;
17'h15aa9:	data_out=16'h2c6;
17'h15aaa:	data_out=16'h89ff;
17'h15aab:	data_out=16'h3e9;
17'h15aac:	data_out=16'h89c9;
17'h15aad:	data_out=16'h84e5;
17'h15aae:	data_out=16'h8a00;
17'h15aaf:	data_out=16'h89ff;
17'h15ab0:	data_out=16'h8900;
17'h15ab1:	data_out=16'h8a00;
17'h15ab2:	data_out=16'h8a00;
17'h15ab3:	data_out=16'ha00;
17'h15ab4:	data_out=16'h8a00;
17'h15ab5:	data_out=16'h89da;
17'h15ab6:	data_out=16'h89ff;
17'h15ab7:	data_out=16'h4d0;
17'h15ab8:	data_out=16'h8a00;
17'h15ab9:	data_out=16'ha00;
17'h15aba:	data_out=16'h8866;
17'h15abb:	data_out=16'h89ff;
17'h15abc:	data_out=16'ha00;
17'h15abd:	data_out=16'h892a;
17'h15abe:	data_out=16'h541;
17'h15abf:	data_out=16'h89fd;
17'h15ac0:	data_out=16'h87f4;
17'h15ac1:	data_out=16'ha00;
17'h15ac2:	data_out=16'h89fd;
17'h15ac3:	data_out=16'h9f6;
17'h15ac4:	data_out=16'h89a9;
17'h15ac5:	data_out=16'h8354;
17'h15ac6:	data_out=16'ha00;
17'h15ac7:	data_out=16'h89ff;
17'h15ac8:	data_out=16'h8a00;
17'h15ac9:	data_out=16'h891;
17'h15aca:	data_out=16'h8a00;
17'h15acb:	data_out=16'h89fe;
17'h15acc:	data_out=16'h89fc;
17'h15acd:	data_out=16'h9fd;
17'h15ace:	data_out=16'h89f7;
17'h15acf:	data_out=16'h89fc;
17'h15ad0:	data_out=16'h9ef;
17'h15ad1:	data_out=16'ha00;
17'h15ad2:	data_out=16'h88a0;
17'h15ad3:	data_out=16'h8a00;
17'h15ad4:	data_out=16'h89ff;
17'h15ad5:	data_out=16'ha00;
17'h15ad6:	data_out=16'ha00;
17'h15ad7:	data_out=16'ha00;
17'h15ad8:	data_out=16'ha00;
17'h15ad9:	data_out=16'h89c4;
17'h15ada:	data_out=16'h704;
17'h15adb:	data_out=16'h89c1;
17'h15adc:	data_out=16'h8998;
17'h15add:	data_out=16'h8a00;
17'h15ade:	data_out=16'h89ff;
17'h15adf:	data_out=16'h8a00;
17'h15ae0:	data_out=16'h89e5;
17'h15ae1:	data_out=16'h89fc;
17'h15ae2:	data_out=16'h83d;
17'h15ae3:	data_out=16'h9fd;
17'h15ae4:	data_out=16'h89ef;
17'h15ae5:	data_out=16'h8a00;
17'h15ae6:	data_out=16'h8356;
17'h15ae7:	data_out=16'h8014;
17'h15ae8:	data_out=16'h51e;
17'h15ae9:	data_out=16'h84ce;
17'h15aea:	data_out=16'h50e;
17'h15aeb:	data_out=16'h896d;
17'h15aec:	data_out=16'h89ff;
17'h15aed:	data_out=16'h9fe;
17'h15aee:	data_out=16'h50d;
17'h15aef:	data_out=16'h8a00;
17'h15af0:	data_out=16'h502;
17'h15af1:	data_out=16'h89ff;
17'h15af2:	data_out=16'h89cf;
17'h15af3:	data_out=16'h8a00;
17'h15af4:	data_out=16'h892c;
17'h15af5:	data_out=16'h79b;
17'h15af6:	data_out=16'h44a;
17'h15af7:	data_out=16'h940;
17'h15af8:	data_out=16'h9f1;
17'h15af9:	data_out=16'h88c4;
17'h15afa:	data_out=16'h9fe;
17'h15afb:	data_out=16'h540;
17'h15afc:	data_out=16'h89a7;
17'h15afd:	data_out=16'h9eb;
17'h15afe:	data_out=16'h9ff;
17'h15aff:	data_out=16'h81ef;
17'h15b00:	data_out=16'h8994;
17'h15b01:	data_out=16'h8a00;
17'h15b02:	data_out=16'h8334;
17'h15b03:	data_out=16'h811b;
17'h15b04:	data_out=16'h881c;
17'h15b05:	data_out=16'h89ee;
17'h15b06:	data_out=16'h8dc;
17'h15b07:	data_out=16'h8a00;
17'h15b08:	data_out=16'h845a;
17'h15b09:	data_out=16'h9de;
17'h15b0a:	data_out=16'h89f3;
17'h15b0b:	data_out=16'h9fb;
17'h15b0c:	data_out=16'h8a00;
17'h15b0d:	data_out=16'h832d;
17'h15b0e:	data_out=16'h229;
17'h15b0f:	data_out=16'h8a00;
17'h15b10:	data_out=16'ha00;
17'h15b11:	data_out=16'h8986;
17'h15b12:	data_out=16'h8657;
17'h15b13:	data_out=16'h833b;
17'h15b14:	data_out=16'ha00;
17'h15b15:	data_out=16'hb9;
17'h15b16:	data_out=16'h89d6;
17'h15b17:	data_out=16'h9ee;
17'h15b18:	data_out=16'h472;
17'h15b19:	data_out=16'h8a00;
17'h15b1a:	data_out=16'h89ca;
17'h15b1b:	data_out=16'h8775;
17'h15b1c:	data_out=16'h8609;
17'h15b1d:	data_out=16'h8a00;
17'h15b1e:	data_out=16'h52e;
17'h15b1f:	data_out=16'h955;
17'h15b20:	data_out=16'h8963;
17'h15b21:	data_out=16'h234;
17'h15b22:	data_out=16'ha00;
17'h15b23:	data_out=16'h89e2;
17'h15b24:	data_out=16'h89e2;
17'h15b25:	data_out=16'h6db;
17'h15b26:	data_out=16'h9fa;
17'h15b27:	data_out=16'h89de;
17'h15b28:	data_out=16'h268;
17'h15b29:	data_out=16'h814c;
17'h15b2a:	data_out=16'h8a00;
17'h15b2b:	data_out=16'h374;
17'h15b2c:	data_out=16'h8736;
17'h15b2d:	data_out=16'h834f;
17'h15b2e:	data_out=16'h8455;
17'h15b2f:	data_out=16'h8a00;
17'h15b30:	data_out=16'h899b;
17'h15b31:	data_out=16'h89e8;
17'h15b32:	data_out=16'h8a00;
17'h15b33:	data_out=16'ha00;
17'h15b34:	data_out=16'h8a00;
17'h15b35:	data_out=16'h892e;
17'h15b36:	data_out=16'h89fe;
17'h15b37:	data_out=16'h82b6;
17'h15b38:	data_out=16'h89dd;
17'h15b39:	data_out=16'ha00;
17'h15b3a:	data_out=16'h817b;
17'h15b3b:	data_out=16'h89ea;
17'h15b3c:	data_out=16'h8306;
17'h15b3d:	data_out=16'h770;
17'h15b3e:	data_out=16'h268;
17'h15b3f:	data_out=16'h89ed;
17'h15b40:	data_out=16'h594;
17'h15b41:	data_out=16'h8f8;
17'h15b42:	data_out=16'h89fe;
17'h15b43:	data_out=16'ha00;
17'h15b44:	data_out=16'h887d;
17'h15b45:	data_out=16'h6c;
17'h15b46:	data_out=16'h487;
17'h15b47:	data_out=16'h8640;
17'h15b48:	data_out=16'h87d9;
17'h15b49:	data_out=16'h8e8;
17'h15b4a:	data_out=16'h8a00;
17'h15b4b:	data_out=16'h89ff;
17'h15b4c:	data_out=16'h89ff;
17'h15b4d:	data_out=16'h9ff;
17'h15b4e:	data_out=16'h89fd;
17'h15b4f:	data_out=16'h88e7;
17'h15b50:	data_out=16'h9fd;
17'h15b51:	data_out=16'ha00;
17'h15b52:	data_out=16'h8795;
17'h15b53:	data_out=16'h8a00;
17'h15b54:	data_out=16'h89f2;
17'h15b55:	data_out=16'ha00;
17'h15b56:	data_out=16'ha00;
17'h15b57:	data_out=16'ha00;
17'h15b58:	data_out=16'ha00;
17'h15b59:	data_out=16'h4d3;
17'h15b5a:	data_out=16'h89d7;
17'h15b5b:	data_out=16'h890a;
17'h15b5c:	data_out=16'h89f7;
17'h15b5d:	data_out=16'h89fb;
17'h15b5e:	data_out=16'h89ff;
17'h15b5f:	data_out=16'h8a00;
17'h15b60:	data_out=16'h88be;
17'h15b61:	data_out=16'h89e3;
17'h15b62:	data_out=16'h707;
17'h15b63:	data_out=16'h9fd;
17'h15b64:	data_out=16'h8663;
17'h15b65:	data_out=16'h89ea;
17'h15b66:	data_out=16'h863c;
17'h15b67:	data_out=16'h3ad;
17'h15b68:	data_out=16'h24c;
17'h15b69:	data_out=16'h8492;
17'h15b6a:	data_out=16'h22f;
17'h15b6b:	data_out=16'h8919;
17'h15b6c:	data_out=16'h8a00;
17'h15b6d:	data_out=16'h9ff;
17'h15b6e:	data_out=16'h22f;
17'h15b6f:	data_out=16'h8a00;
17'h15b70:	data_out=16'h22a;
17'h15b71:	data_out=16'h8a00;
17'h15b72:	data_out=16'h8971;
17'h15b73:	data_out=16'h89f0;
17'h15b74:	data_out=16'h89a9;
17'h15b75:	data_out=16'h89b8;
17'h15b76:	data_out=16'h615;
17'h15b77:	data_out=16'h9ce;
17'h15b78:	data_out=16'h9ff;
17'h15b79:	data_out=16'h89b2;
17'h15b7a:	data_out=16'h9fd;
17'h15b7b:	data_out=16'h268;
17'h15b7c:	data_out=16'h84e7;
17'h15b7d:	data_out=16'h9fb;
17'h15b7e:	data_out=16'ha00;
17'h15b7f:	data_out=16'h2d3;
17'h15b80:	data_out=16'h8444;
17'h15b81:	data_out=16'h8a00;
17'h15b82:	data_out=16'h82b2;
17'h15b83:	data_out=16'h8242;
17'h15b84:	data_out=16'h88b0;
17'h15b85:	data_out=16'h8931;
17'h15b86:	data_out=16'h65c;
17'h15b87:	data_out=16'h8a00;
17'h15b88:	data_out=16'h342;
17'h15b89:	data_out=16'h9d9;
17'h15b8a:	data_out=16'h89e8;
17'h15b8b:	data_out=16'h9fe;
17'h15b8c:	data_out=16'h8a00;
17'h15b8d:	data_out=16'h86ae;
17'h15b8e:	data_out=16'he4;
17'h15b8f:	data_out=16'h89af;
17'h15b90:	data_out=16'h87c;
17'h15b91:	data_out=16'h89d2;
17'h15b92:	data_out=16'h8a00;
17'h15b93:	data_out=16'h857c;
17'h15b94:	data_out=16'h7a6;
17'h15b95:	data_out=16'h122;
17'h15b96:	data_out=16'h8681;
17'h15b97:	data_out=16'h226;
17'h15b98:	data_out=16'h17c;
17'h15b99:	data_out=16'h85b7;
17'h15b9a:	data_out=16'h89e3;
17'h15b9b:	data_out=16'h883a;
17'h15b9c:	data_out=16'h849d;
17'h15b9d:	data_out=16'h8a00;
17'h15b9e:	data_out=16'h8322;
17'h15b9f:	data_out=16'h8ca;
17'h15ba0:	data_out=16'h89dd;
17'h15ba1:	data_out=16'hea;
17'h15ba2:	data_out=16'h9d0;
17'h15ba3:	data_out=16'h8666;
17'h15ba4:	data_out=16'h865f;
17'h15ba5:	data_out=16'h47c;
17'h15ba6:	data_out=16'h9fc;
17'h15ba7:	data_out=16'h89fa;
17'h15ba8:	data_out=16'h10a;
17'h15ba9:	data_out=16'h8362;
17'h15baa:	data_out=16'h8a00;
17'h15bab:	data_out=16'h1de;
17'h15bac:	data_out=16'h83c6;
17'h15bad:	data_out=16'h218;
17'h15bae:	data_out=16'h87fd;
17'h15baf:	data_out=16'h8a00;
17'h15bb0:	data_out=16'h89b0;
17'h15bb1:	data_out=16'h89f5;
17'h15bb2:	data_out=16'h89ff;
17'h15bb3:	data_out=16'h6ab;
17'h15bb4:	data_out=16'h8a00;
17'h15bb5:	data_out=16'h8922;
17'h15bb6:	data_out=16'h87ff;
17'h15bb7:	data_out=16'h8261;
17'h15bb8:	data_out=16'h89fa;
17'h15bb9:	data_out=16'h466;
17'h15bba:	data_out=16'h829e;
17'h15bbb:	data_out=16'h89ce;
17'h15bbc:	data_out=16'h8109;
17'h15bbd:	data_out=16'h660;
17'h15bbe:	data_out=16'h10b;
17'h15bbf:	data_out=16'h8913;
17'h15bc0:	data_out=16'h748;
17'h15bc1:	data_out=16'h683;
17'h15bc2:	data_out=16'h89f4;
17'h15bc3:	data_out=16'ha00;
17'h15bc4:	data_out=16'h8342;
17'h15bc5:	data_out=16'hf7;
17'h15bc6:	data_out=16'h62f;
17'h15bc7:	data_out=16'h8606;
17'h15bc8:	data_out=16'h8a00;
17'h15bc9:	data_out=16'h6c2;
17'h15bca:	data_out=16'h8a00;
17'h15bcb:	data_out=16'h8a00;
17'h15bcc:	data_out=16'h8a00;
17'h15bcd:	data_out=16'h9de;
17'h15bce:	data_out=16'h8a00;
17'h15bcf:	data_out=16'h8981;
17'h15bd0:	data_out=16'h9ff;
17'h15bd1:	data_out=16'h930;
17'h15bd2:	data_out=16'h84fc;
17'h15bd3:	data_out=16'h8a00;
17'h15bd4:	data_out=16'h8a00;
17'h15bd5:	data_out=16'h9fe;
17'h15bd6:	data_out=16'ha00;
17'h15bd7:	data_out=16'ha00;
17'h15bd8:	data_out=16'ha00;
17'h15bd9:	data_out=16'h3ab;
17'h15bda:	data_out=16'h89e4;
17'h15bdb:	data_out=16'h8949;
17'h15bdc:	data_out=16'h89ee;
17'h15bdd:	data_out=16'h8a00;
17'h15bde:	data_out=16'h8a00;
17'h15bdf:	data_out=16'h8a00;
17'h15be0:	data_out=16'h84b3;
17'h15be1:	data_out=16'h8906;
17'h15be2:	data_out=16'h9b;
17'h15be3:	data_out=16'h61d;
17'h15be4:	data_out=16'h8339;
17'h15be5:	data_out=16'h89f5;
17'h15be6:	data_out=16'h826a;
17'h15be7:	data_out=16'h80b0;
17'h15be8:	data_out=16'hf9;
17'h15be9:	data_out=16'h269;
17'h15bea:	data_out=16'he8;
17'h15beb:	data_out=16'h8875;
17'h15bec:	data_out=16'h89fb;
17'h15bed:	data_out=16'h5d6;
17'h15bee:	data_out=16'he8;
17'h15bef:	data_out=16'h89ff;
17'h15bf0:	data_out=16'he5;
17'h15bf1:	data_out=16'h8a00;
17'h15bf2:	data_out=16'h89cc;
17'h15bf3:	data_out=16'h89f9;
17'h15bf4:	data_out=16'h89b2;
17'h15bf5:	data_out=16'h8739;
17'h15bf6:	data_out=16'h386;
17'h15bf7:	data_out=16'h9f0;
17'h15bf8:	data_out=16'h4e5;
17'h15bf9:	data_out=16'h89aa;
17'h15bfa:	data_out=16'h67d;
17'h15bfb:	data_out=16'h10a;
17'h15bfc:	data_out=16'h8423;
17'h15bfd:	data_out=16'h53b;
17'h15bfe:	data_out=16'ha00;
17'h15bff:	data_out=16'hba;
17'h15c00:	data_out=16'ha00;
17'h15c01:	data_out=16'h84d6;
17'h15c02:	data_out=16'h85b6;
17'h15c03:	data_out=16'h8209;
17'h15c04:	data_out=16'h2b6;
17'h15c05:	data_out=16'h80f9;
17'h15c06:	data_out=16'h840e;
17'h15c07:	data_out=16'h8595;
17'h15c08:	data_out=16'h8086;
17'h15c09:	data_out=16'h94e;
17'h15c0a:	data_out=16'h8386;
17'h15c0b:	data_out=16'h8720;
17'h15c0c:	data_out=16'h8a00;
17'h15c0d:	data_out=16'h86aa;
17'h15c0e:	data_out=16'h8152;
17'h15c0f:	data_out=16'h893d;
17'h15c10:	data_out=16'h4b2;
17'h15c11:	data_out=16'h8105;
17'h15c12:	data_out=16'h8a00;
17'h15c13:	data_out=16'h8571;
17'h15c14:	data_out=16'h8259;
17'h15c15:	data_out=16'h422;
17'h15c16:	data_out=16'h80f0;
17'h15c17:	data_out=16'h86d5;
17'h15c18:	data_out=16'h800e;
17'h15c19:	data_out=16'ha7;
17'h15c1a:	data_out=16'h8038;
17'h15c1b:	data_out=16'h89fb;
17'h15c1c:	data_out=16'h2ad;
17'h15c1d:	data_out=16'h8367;
17'h15c1e:	data_out=16'h851c;
17'h15c1f:	data_out=16'h1ce;
17'h15c20:	data_out=16'h87b;
17'h15c21:	data_out=16'h8156;
17'h15c22:	data_out=16'h581;
17'h15c23:	data_out=16'h8245;
17'h15c24:	data_out=16'h823f;
17'h15c25:	data_out=16'h38;
17'h15c26:	data_out=16'h8059;
17'h15c27:	data_out=16'h824c;
17'h15c28:	data_out=16'h815e;
17'h15c29:	data_out=16'h828a;
17'h15c2a:	data_out=16'h8a00;
17'h15c2b:	data_out=16'h3aa;
17'h15c2c:	data_out=16'h3d;
17'h15c2d:	data_out=16'h8574;
17'h15c2e:	data_out=16'h89ec;
17'h15c2f:	data_out=16'h82ac;
17'h15c30:	data_out=16'h8a00;
17'h15c31:	data_out=16'h8599;
17'h15c32:	data_out=16'h8a00;
17'h15c33:	data_out=16'h8098;
17'h15c34:	data_out=16'h81b6;
17'h15c35:	data_out=16'h8374;
17'h15c36:	data_out=16'h83db;
17'h15c37:	data_out=16'h8615;
17'h15c38:	data_out=16'h8033;
17'h15c39:	data_out=16'h80c7;
17'h15c3a:	data_out=16'h80f0;
17'h15c3b:	data_out=16'h8003;
17'h15c3c:	data_out=16'h85f0;
17'h15c3d:	data_out=16'h9ff;
17'h15c3e:	data_out=16'h815f;
17'h15c3f:	data_out=16'h80df;
17'h15c40:	data_out=16'h1ea;
17'h15c41:	data_out=16'h819c;
17'h15c42:	data_out=16'h8a00;
17'h15c43:	data_out=16'h82e3;
17'h15c44:	data_out=16'h3df;
17'h15c45:	data_out=16'h404;
17'h15c46:	data_out=16'h8053;
17'h15c47:	data_out=16'h8453;
17'h15c48:	data_out=16'h88e3;
17'h15c49:	data_out=16'h158;
17'h15c4a:	data_out=16'h8898;
17'h15c4b:	data_out=16'h8a00;
17'h15c4c:	data_out=16'h88f1;
17'h15c4d:	data_out=16'h5da;
17'h15c4e:	data_out=16'h8a00;
17'h15c4f:	data_out=16'h8679;
17'h15c50:	data_out=16'h416;
17'h15c51:	data_out=16'h811f;
17'h15c52:	data_out=16'h8121;
17'h15c53:	data_out=16'h8a00;
17'h15c54:	data_out=16'h1e2;
17'h15c55:	data_out=16'h108;
17'h15c56:	data_out=16'h114;
17'h15c57:	data_out=16'h1ca;
17'h15c58:	data_out=16'h8065;
17'h15c59:	data_out=16'ha3;
17'h15c5a:	data_out=16'h89ff;
17'h15c5b:	data_out=16'h15d;
17'h15c5c:	data_out=16'h83af;
17'h15c5d:	data_out=16'h8687;
17'h15c5e:	data_out=16'h832f;
17'h15c5f:	data_out=16'h8219;
17'h15c60:	data_out=16'h86e0;
17'h15c61:	data_out=16'h2d8;
17'h15c62:	data_out=16'h8a00;
17'h15c63:	data_out=16'h8129;
17'h15c64:	data_out=16'h458;
17'h15c65:	data_out=16'h8363;
17'h15c66:	data_out=16'haf;
17'h15c67:	data_out=16'h851f;
17'h15c68:	data_out=16'h8157;
17'h15c69:	data_out=16'h82b1;
17'h15c6a:	data_out=16'h814e;
17'h15c6b:	data_out=16'h444;
17'h15c6c:	data_out=16'h89e8;
17'h15c6d:	data_out=16'h810f;
17'h15c6e:	data_out=16'h814f;
17'h15c6f:	data_out=16'h8842;
17'h15c70:	data_out=16'h8151;
17'h15c71:	data_out=16'h8a00;
17'h15c72:	data_out=16'h81e7;
17'h15c73:	data_out=16'h1a7;
17'h15c74:	data_out=16'h8a00;
17'h15c75:	data_out=16'h8a00;
17'h15c76:	data_out=16'h296;
17'h15c77:	data_out=16'h619;
17'h15c78:	data_out=16'h8506;
17'h15c79:	data_out=16'h89db;
17'h15c7a:	data_out=16'h8226;
17'h15c7b:	data_out=16'h8160;
17'h15c7c:	data_out=16'h80ec;
17'h15c7d:	data_out=16'h849f;
17'h15c7e:	data_out=16'h995;
17'h15c7f:	data_out=16'h45f;
17'h15c80:	data_out=16'h45c;
17'h15c81:	data_out=16'h8209;
17'h15c82:	data_out=16'h838d;
17'h15c83:	data_out=16'h80cb;
17'h15c84:	data_out=16'h22d;
17'h15c85:	data_out=16'h4;
17'h15c86:	data_out=16'h34;
17'h15c87:	data_out=16'h8;
17'h15c88:	data_out=16'h83a9;
17'h15c89:	data_out=16'h466;
17'h15c8a:	data_out=16'h81df;
17'h15c8b:	data_out=16'h84ab;
17'h15c8c:	data_out=16'h86d2;
17'h15c8d:	data_out=16'h813b;
17'h15c8e:	data_out=16'h8125;
17'h15c8f:	data_out=16'h8374;
17'h15c90:	data_out=16'h42;
17'h15c91:	data_out=16'h19c;
17'h15c92:	data_out=16'h83c6;
17'h15c93:	data_out=16'h807b;
17'h15c94:	data_out=16'h8169;
17'h15c95:	data_out=16'h15b;
17'h15c96:	data_out=16'h80d6;
17'h15c97:	data_out=16'h8273;
17'h15c98:	data_out=16'h809a;
17'h15c99:	data_out=16'h1e8;
17'h15c9a:	data_out=16'h195;
17'h15c9b:	data_out=16'h8255;
17'h15c9c:	data_out=16'h77;
17'h15c9d:	data_out=16'h816f;
17'h15c9e:	data_out=16'h8131;
17'h15c9f:	data_out=16'he6;
17'h15ca0:	data_out=16'h354;
17'h15ca1:	data_out=16'h811f;
17'h15ca2:	data_out=16'h299;
17'h15ca3:	data_out=16'h82d3;
17'h15ca4:	data_out=16'h82d2;
17'h15ca5:	data_out=16'h4c;
17'h15ca6:	data_out=16'h80d8;
17'h15ca7:	data_out=16'h811e;
17'h15ca8:	data_out=16'h8118;
17'h15ca9:	data_out=16'h71;
17'h15caa:	data_out=16'h85a9;
17'h15cab:	data_out=16'h25c;
17'h15cac:	data_out=16'h800d;
17'h15cad:	data_out=16'h823b;
17'h15cae:	data_out=16'h847c;
17'h15caf:	data_out=16'h80e1;
17'h15cb0:	data_out=16'h83f1;
17'h15cb1:	data_out=16'h257;
17'h15cb2:	data_out=16'h83ab;
17'h15cb3:	data_out=16'h80b7;
17'h15cb4:	data_out=16'h282;
17'h15cb5:	data_out=16'h83e5;
17'h15cb6:	data_out=16'h84bf;
17'h15cb7:	data_out=16'h834a;
17'h15cb8:	data_out=16'h2f5;
17'h15cb9:	data_out=16'h12;
17'h15cba:	data_out=16'hb5;
17'h15cbb:	data_out=16'h7a;
17'h15cbc:	data_out=16'h85cd;
17'h15cbd:	data_out=16'h65c;
17'h15cbe:	data_out=16'h8115;
17'h15cbf:	data_out=16'h1c;
17'h15cc0:	data_out=16'h111;
17'h15cc1:	data_out=16'h8545;
17'h15cc2:	data_out=16'h8583;
17'h15cc3:	data_out=16'h8045;
17'h15cc4:	data_out=16'h148;
17'h15cc5:	data_out=16'h14d;
17'h15cc6:	data_out=16'h827c;
17'h15cc7:	data_out=16'h8059;
17'h15cc8:	data_out=16'h81b8;
17'h15cc9:	data_out=16'h110;
17'h15cca:	data_out=16'h8274;
17'h15ccb:	data_out=16'h87cc;
17'h15ccc:	data_out=16'h82d8;
17'h15ccd:	data_out=16'h311;
17'h15cce:	data_out=16'h8519;
17'h15ccf:	data_out=16'h81c7;
17'h15cd0:	data_out=16'hc2;
17'h15cd1:	data_out=16'h832f;
17'h15cd2:	data_out=16'h827e;
17'h15cd3:	data_out=16'h8220;
17'h15cd4:	data_out=16'h801b;
17'h15cd5:	data_out=16'h85cc;
17'h15cd6:	data_out=16'h80d3;
17'h15cd7:	data_out=16'h801c;
17'h15cd8:	data_out=16'h8662;
17'h15cd9:	data_out=16'h4;
17'h15cda:	data_out=16'h8467;
17'h15cdb:	data_out=16'h821c;
17'h15cdc:	data_out=16'h80a3;
17'h15cdd:	data_out=16'h82e1;
17'h15cde:	data_out=16'h8109;
17'h15cdf:	data_out=16'h809b;
17'h15ce0:	data_out=16'h827b;
17'h15ce1:	data_out=16'he1;
17'h15ce2:	data_out=16'h844e;
17'h15ce3:	data_out=16'h80d6;
17'h15ce4:	data_out=16'h3fd;
17'h15ce5:	data_out=16'h256;
17'h15ce6:	data_out=16'h28d;
17'h15ce7:	data_out=16'h81cd;
17'h15ce8:	data_out=16'h8120;
17'h15ce9:	data_out=16'h8591;
17'h15cea:	data_out=16'h8133;
17'h15ceb:	data_out=16'h439;
17'h15cec:	data_out=16'h850a;
17'h15ced:	data_out=16'h80cd;
17'h15cee:	data_out=16'h8132;
17'h15cef:	data_out=16'h808c;
17'h15cf0:	data_out=16'h8134;
17'h15cf1:	data_out=16'h8445;
17'h15cf2:	data_out=16'h49;
17'h15cf3:	data_out=16'h2b3;
17'h15cf4:	data_out=16'h8412;
17'h15cf5:	data_out=16'h8589;
17'h15cf6:	data_out=16'h27e;
17'h15cf7:	data_out=16'ha8;
17'h15cf8:	data_out=16'heb;
17'h15cf9:	data_out=16'h86d6;
17'h15cfa:	data_out=16'h8148;
17'h15cfb:	data_out=16'h8112;
17'h15cfc:	data_out=16'h812c;
17'h15cfd:	data_out=16'h87;
17'h15cfe:	data_out=16'h3d8;
17'h15cff:	data_out=16'h8a;
17'h15d00:	data_out=16'hf5;
17'h15d01:	data_out=16'h1e;
17'h15d02:	data_out=16'h8085;
17'h15d03:	data_out=16'h8004;
17'h15d04:	data_out=16'h8004;
17'h15d05:	data_out=16'h8003;
17'h15d06:	data_out=16'h805c;
17'h15d07:	data_out=16'h1c;
17'h15d08:	data_out=16'h48;
17'h15d09:	data_out=16'h9b;
17'h15d0a:	data_out=16'h8024;
17'h15d0b:	data_out=16'h8045;
17'h15d0c:	data_out=16'h802d;
17'h15d0d:	data_out=16'h72;
17'h15d0e:	data_out=16'h801a;
17'h15d0f:	data_out=16'h28;
17'h15d10:	data_out=16'h802c;
17'h15d11:	data_out=16'h51;
17'h15d12:	data_out=16'h807f;
17'h15d13:	data_out=16'h8a;
17'h15d14:	data_out=16'h8058;
17'h15d15:	data_out=16'ha1;
17'h15d16:	data_out=16'h9c;
17'h15d17:	data_out=16'h8052;
17'h15d18:	data_out=16'h8004;
17'h15d19:	data_out=16'hac;
17'h15d1a:	data_out=16'h11;
17'h15d1b:	data_out=16'h42;
17'h15d1c:	data_out=16'h32;
17'h15d1d:	data_out=16'h803c;
17'h15d1e:	data_out=16'h11;
17'h15d1f:	data_out=16'h8049;
17'h15d20:	data_out=16'h2f;
17'h15d21:	data_out=16'h8020;
17'h15d22:	data_out=16'hc;
17'h15d23:	data_out=16'h809d;
17'h15d24:	data_out=16'h8099;
17'h15d25:	data_out=16'h8025;
17'h15d26:	data_out=16'h64;
17'h15d27:	data_out=16'h8039;
17'h15d28:	data_out=16'h8021;
17'h15d29:	data_out=16'h13;
17'h15d2a:	data_out=16'h8022;
17'h15d2b:	data_out=16'h85;
17'h15d2c:	data_out=16'h23;
17'h15d2d:	data_out=16'h8055;
17'h15d2e:	data_out=16'h8082;
17'h15d2f:	data_out=16'h1b;
17'h15d30:	data_out=16'h801a;
17'h15d31:	data_out=16'he0;
17'h15d32:	data_out=16'h801d;
17'h15d33:	data_out=16'h8020;
17'h15d34:	data_out=16'h7d;
17'h15d35:	data_out=16'h8063;
17'h15d36:	data_out=16'h8092;
17'h15d37:	data_out=16'h8082;
17'h15d38:	data_out=16'h8a;
17'h15d39:	data_out=16'h30;
17'h15d3a:	data_out=16'h8060;
17'h15d3b:	data_out=16'ha2;
17'h15d3c:	data_out=16'h80a6;
17'h15d3d:	data_out=16'hef;
17'h15d3e:	data_out=16'h8024;
17'h15d3f:	data_out=16'h13;
17'h15d40:	data_out=16'h8064;
17'h15d41:	data_out=16'h8062;
17'h15d42:	data_out=16'h804c;
17'h15d43:	data_out=16'h805b;
17'h15d44:	data_out=16'h34;
17'h15d45:	data_out=16'h93;
17'h15d46:	data_out=16'h8068;
17'h15d47:	data_out=16'h806c;
17'h15d48:	data_out=16'h8063;
17'h15d49:	data_out=16'h8018;
17'h15d4a:	data_out=16'h8046;
17'h15d4b:	data_out=16'h807b;
17'h15d4c:	data_out=16'h8074;
17'h15d4d:	data_out=16'h4b;
17'h15d4e:	data_out=16'h8002;
17'h15d4f:	data_out=16'h8063;
17'h15d50:	data_out=16'h8067;
17'h15d51:	data_out=16'h5d;
17'h15d52:	data_out=16'h806a;
17'h15d53:	data_out=16'h8003;
17'h15d54:	data_out=16'h8002;
17'h15d55:	data_out=16'h809f;
17'h15d56:	data_out=16'h8064;
17'h15d57:	data_out=16'h8077;
17'h15d58:	data_out=16'h80b8;
17'h15d59:	data_out=16'h8087;
17'h15d5a:	data_out=16'h808a;
17'h15d5b:	data_out=16'h8043;
17'h15d5c:	data_out=16'h8014;
17'h15d5d:	data_out=16'h8001;
17'h15d5e:	data_out=16'h8;
17'h15d5f:	data_out=16'h8017;
17'h15d60:	data_out=16'h1a;
17'h15d61:	data_out=16'h57;
17'h15d62:	data_out=16'h805b;
17'h15d63:	data_out=16'h8034;
17'h15d64:	data_out=16'h4d;
17'h15d65:	data_out=16'h18;
17'h15d66:	data_out=16'h63;
17'h15d67:	data_out=16'h808d;
17'h15d68:	data_out=16'h801d;
17'h15d69:	data_out=16'h809b;
17'h15d6a:	data_out=16'h8028;
17'h15d6b:	data_out=16'hbb;
17'h15d6c:	data_out=16'h8068;
17'h15d6d:	data_out=16'h8022;
17'h15d6e:	data_out=16'h8024;
17'h15d6f:	data_out=16'ha;
17'h15d70:	data_out=16'h801e;
17'h15d71:	data_out=16'h8057;
17'h15d72:	data_out=16'h3;
17'h15d73:	data_out=16'h66;
17'h15d74:	data_out=16'h801f;
17'h15d75:	data_out=16'h800e;
17'h15d76:	data_out=16'h9f;
17'h15d77:	data_out=16'h8043;
17'h15d78:	data_out=16'h84;
17'h15d79:	data_out=16'h808a;
17'h15d7a:	data_out=16'h804a;
17'h15d7b:	data_out=16'h8016;
17'h15d7c:	data_out=16'h804b;
17'h15d7d:	data_out=16'h805b;
17'h15d7e:	data_out=16'h98;
17'h15d7f:	data_out=16'h8045;
17'h15d80:	data_out=16'h8001;
17'h15d81:	data_out=16'h8007;
17'h15d82:	data_out=16'h8004;
17'h15d83:	data_out=16'h1;
17'h15d84:	data_out=16'h8003;
17'h15d85:	data_out=16'h9;
17'h15d86:	data_out=16'h4;
17'h15d87:	data_out=16'h7;
17'h15d88:	data_out=16'h8006;
17'h15d89:	data_out=16'h6;
17'h15d8a:	data_out=16'h1;
17'h15d8b:	data_out=16'h8;
17'h15d8c:	data_out=16'h8007;
17'h15d8d:	data_out=16'h7;
17'h15d8e:	data_out=16'h8007;
17'h15d8f:	data_out=16'h5;
17'h15d90:	data_out=16'h2;
17'h15d91:	data_out=16'h8005;
17'h15d92:	data_out=16'h8003;
17'h15d93:	data_out=16'h8008;
17'h15d94:	data_out=16'h4;
17'h15d95:	data_out=16'h7;
17'h15d96:	data_out=16'h1;
17'h15d97:	data_out=16'h8001;
17'h15d98:	data_out=16'h8002;
17'h15d99:	data_out=16'h8006;
17'h15d9a:	data_out=16'h8003;
17'h15d9b:	data_out=16'h8008;
17'h15d9c:	data_out=16'h8006;
17'h15d9d:	data_out=16'h4;
17'h15d9e:	data_out=16'h9;
17'h15d9f:	data_out=16'h3;
17'h15da0:	data_out=16'h6;
17'h15da1:	data_out=16'h8004;
17'h15da2:	data_out=16'h8006;
17'h15da3:	data_out=16'h8006;
17'h15da4:	data_out=16'h8005;
17'h15da5:	data_out=16'h7;
17'h15da6:	data_out=16'h8007;
17'h15da7:	data_out=16'h8002;
17'h15da8:	data_out=16'h5;
17'h15da9:	data_out=16'h3;
17'h15daa:	data_out=16'h8003;
17'h15dab:	data_out=16'h7;
17'h15dac:	data_out=16'h0;
17'h15dad:	data_out=16'h8000;
17'h15dae:	data_out=16'h2;
17'h15daf:	data_out=16'h8007;
17'h15db0:	data_out=16'h4;
17'h15db1:	data_out=16'h8;
17'h15db2:	data_out=16'h8006;
17'h15db3:	data_out=16'h8001;
17'h15db4:	data_out=16'h6;
17'h15db5:	data_out=16'h4;
17'h15db6:	data_out=16'h7;
17'h15db7:	data_out=16'h8005;
17'h15db8:	data_out=16'h8;
17'h15db9:	data_out=16'h8004;
17'h15dba:	data_out=16'h8005;
17'h15dbb:	data_out=16'h8007;
17'h15dbc:	data_out=16'h9;
17'h15dbd:	data_out=16'h8005;
17'h15dbe:	data_out=16'h4;
17'h15dbf:	data_out=16'h6;
17'h15dc0:	data_out=16'h0;
17'h15dc1:	data_out=16'h8;
17'h15dc2:	data_out=16'h8009;
17'h15dc3:	data_out=16'h4;
17'h15dc4:	data_out=16'h6;
17'h15dc5:	data_out=16'h8007;
17'h15dc6:	data_out=16'h8007;
17'h15dc7:	data_out=16'h1;
17'h15dc8:	data_out=16'h5;
17'h15dc9:	data_out=16'h0;
17'h15dca:	data_out=16'h8001;
17'h15dcb:	data_out=16'h8004;
17'h15dcc:	data_out=16'h9;
17'h15dcd:	data_out=16'h8008;
17'h15dce:	data_out=16'h8001;
17'h15dcf:	data_out=16'h4;
17'h15dd0:	data_out=16'h8009;
17'h15dd1:	data_out=16'h2;
17'h15dd2:	data_out=16'h8007;
17'h15dd3:	data_out=16'h6;
17'h15dd4:	data_out=16'h8003;
17'h15dd5:	data_out=16'h8009;
17'h15dd6:	data_out=16'h8008;
17'h15dd7:	data_out=16'h8004;
17'h15dd8:	data_out=16'h8004;
17'h15dd9:	data_out=16'h8004;
17'h15dda:	data_out=16'h8002;
17'h15ddb:	data_out=16'h8004;
17'h15ddc:	data_out=16'h1;
17'h15ddd:	data_out=16'h8007;
17'h15dde:	data_out=16'h8007;
17'h15ddf:	data_out=16'h8009;
17'h15de0:	data_out=16'h8009;
17'h15de1:	data_out=16'h8006;
17'h15de2:	data_out=16'h5;
17'h15de3:	data_out=16'h6;
17'h15de4:	data_out=16'h8004;
17'h15de5:	data_out=16'h8;
17'h15de6:	data_out=16'h8001;
17'h15de7:	data_out=16'h8008;
17'h15de8:	data_out=16'h8002;
17'h15de9:	data_out=16'h7;
17'h15dea:	data_out=16'h8002;
17'h15deb:	data_out=16'h8002;
17'h15dec:	data_out=16'h8;
17'h15ded:	data_out=16'h6;
17'h15dee:	data_out=16'h8007;
17'h15def:	data_out=16'h9;
17'h15df0:	data_out=16'h8001;
17'h15df1:	data_out=16'h8005;
17'h15df2:	data_out=16'h6;
17'h15df3:	data_out=16'h5;
17'h15df4:	data_out=16'h8004;
17'h15df5:	data_out=16'h7;
17'h15df6:	data_out=16'h8009;
17'h15df7:	data_out=16'h1;
17'h15df8:	data_out=16'h8006;
17'h15df9:	data_out=16'h8002;
17'h15dfa:	data_out=16'h6;
17'h15dfb:	data_out=16'h4;
17'h15dfc:	data_out=16'h0;
17'h15dfd:	data_out=16'h9;
17'h15dfe:	data_out=16'h4;
17'h15dff:	data_out=16'h1;
17'h15e00:	data_out=16'h8007;
17'h15e01:	data_out=16'h0;
17'h15e02:	data_out=16'h8002;
17'h15e03:	data_out=16'h8001;
17'h15e04:	data_out=16'h8002;
17'h15e05:	data_out=16'h5;
17'h15e06:	data_out=16'h0;
17'h15e07:	data_out=16'h6;
17'h15e08:	data_out=16'h3;
17'h15e09:	data_out=16'h7;
17'h15e0a:	data_out=16'h8005;
17'h15e0b:	data_out=16'h2;
17'h15e0c:	data_out=16'h4;
17'h15e0d:	data_out=16'h8003;
17'h15e0e:	data_out=16'h2;
17'h15e0f:	data_out=16'h8007;
17'h15e10:	data_out=16'h1;
17'h15e11:	data_out=16'h8001;
17'h15e12:	data_out=16'h7;
17'h15e13:	data_out=16'h6;
17'h15e14:	data_out=16'h8003;
17'h15e15:	data_out=16'h8;
17'h15e16:	data_out=16'h8002;
17'h15e17:	data_out=16'h8000;
17'h15e18:	data_out=16'h8003;
17'h15e19:	data_out=16'h8005;
17'h15e1a:	data_out=16'h8006;
17'h15e1b:	data_out=16'h6;
17'h15e1c:	data_out=16'h8006;
17'h15e1d:	data_out=16'h8;
17'h15e1e:	data_out=16'h8002;
17'h15e1f:	data_out=16'h8003;
17'h15e20:	data_out=16'h8001;
17'h15e21:	data_out=16'h5;
17'h15e22:	data_out=16'h5;
17'h15e23:	data_out=16'h6;
17'h15e24:	data_out=16'h1;
17'h15e25:	data_out=16'h8005;
17'h15e26:	data_out=16'h3;
17'h15e27:	data_out=16'h8005;
17'h15e28:	data_out=16'h8007;
17'h15e29:	data_out=16'h7;
17'h15e2a:	data_out=16'h6;
17'h15e2b:	data_out=16'h6;
17'h15e2c:	data_out=16'h8005;
17'h15e2d:	data_out=16'h8001;
17'h15e2e:	data_out=16'h9;
17'h15e2f:	data_out=16'h5;
17'h15e30:	data_out=16'h7;
17'h15e31:	data_out=16'h7;
17'h15e32:	data_out=16'h1;
17'h15e33:	data_out=16'h8006;
17'h15e34:	data_out=16'h6;
17'h15e35:	data_out=16'h8;
17'h15e36:	data_out=16'h3;
17'h15e37:	data_out=16'h8007;
17'h15e38:	data_out=16'h8006;
17'h15e39:	data_out=16'h6;
17'h15e3a:	data_out=16'h9;
17'h15e3b:	data_out=16'h8003;
17'h15e3c:	data_out=16'h5;
17'h15e3d:	data_out=16'h8003;
17'h15e3e:	data_out=16'h3;
17'h15e3f:	data_out=16'h8006;
17'h15e40:	data_out=16'h8007;
17'h15e41:	data_out=16'h8002;
17'h15e42:	data_out=16'h8009;
17'h15e43:	data_out=16'h3;
17'h15e44:	data_out=16'h3;
17'h15e45:	data_out=16'h3;
17'h15e46:	data_out=16'h7;
17'h15e47:	data_out=16'h5;
17'h15e48:	data_out=16'h1;
17'h15e49:	data_out=16'h4;
17'h15e4a:	data_out=16'h3;
17'h15e4b:	data_out=16'h5;
17'h15e4c:	data_out=16'h8007;
17'h15e4d:	data_out=16'h2;
17'h15e4e:	data_out=16'h1;
17'h15e4f:	data_out=16'h8009;
17'h15e50:	data_out=16'h8000;
17'h15e51:	data_out=16'h8007;
17'h15e52:	data_out=16'h8006;
17'h15e53:	data_out=16'h8004;
17'h15e54:	data_out=16'h8008;
17'h15e55:	data_out=16'h7;
17'h15e56:	data_out=16'h8001;
17'h15e57:	data_out=16'h8005;
17'h15e58:	data_out=16'h4;
17'h15e59:	data_out=16'h8002;
17'h15e5a:	data_out=16'h1;
17'h15e5b:	data_out=16'h8001;
17'h15e5c:	data_out=16'h5;
17'h15e5d:	data_out=16'h8005;
17'h15e5e:	data_out=16'h3;
17'h15e5f:	data_out=16'h6;
17'h15e60:	data_out=16'h3;
17'h15e61:	data_out=16'h3;
17'h15e62:	data_out=16'h8000;
17'h15e63:	data_out=16'h8003;
17'h15e64:	data_out=16'h8003;
17'h15e65:	data_out=16'h8003;
17'h15e66:	data_out=16'h8007;
17'h15e67:	data_out=16'h8;
17'h15e68:	data_out=16'h8008;
17'h15e69:	data_out=16'h5;
17'h15e6a:	data_out=16'h4;
17'h15e6b:	data_out=16'h8006;
17'h15e6c:	data_out=16'h8003;
17'h15e6d:	data_out=16'h8004;
17'h15e6e:	data_out=16'h8006;
17'h15e6f:	data_out=16'h6;
17'h15e70:	data_out=16'h8002;
17'h15e71:	data_out=16'h8002;
17'h15e72:	data_out=16'h8007;
17'h15e73:	data_out=16'h8000;
17'h15e74:	data_out=16'h8005;
17'h15e75:	data_out=16'h1;
17'h15e76:	data_out=16'h4;
17'h15e77:	data_out=16'h8;
17'h15e78:	data_out=16'h9;
17'h15e79:	data_out=16'h8004;
17'h15e7a:	data_out=16'h8002;
17'h15e7b:	data_out=16'h4;
17'h15e7c:	data_out=16'h1;
17'h15e7d:	data_out=16'h8008;
17'h15e7e:	data_out=16'h1;
17'h15e7f:	data_out=16'h8006;
17'h15e80:	data_out=16'h4;
17'h15e81:	data_out=16'h8008;
17'h15e82:	data_out=16'h8000;
17'h15e83:	data_out=16'h8008;
17'h15e84:	data_out=16'h8002;
17'h15e85:	data_out=16'h2;
17'h15e86:	data_out=16'h8009;
17'h15e87:	data_out=16'h8001;
17'h15e88:	data_out=16'h8003;
17'h15e89:	data_out=16'h4;
17'h15e8a:	data_out=16'h2;
17'h15e8b:	data_out=16'h4;
17'h15e8c:	data_out=16'h8009;
17'h15e8d:	data_out=16'h5;
17'h15e8e:	data_out=16'h1;
17'h15e8f:	data_out=16'h8001;
17'h15e90:	data_out=16'h8006;
17'h15e91:	data_out=16'h4;
17'h15e92:	data_out=16'h7;
17'h15e93:	data_out=16'h8001;
17'h15e94:	data_out=16'h8004;
17'h15e95:	data_out=16'h2;
17'h15e96:	data_out=16'h8002;
17'h15e97:	data_out=16'h8005;
17'h15e98:	data_out=16'h7;
17'h15e99:	data_out=16'h5;
17'h15e9a:	data_out=16'h8;
17'h15e9b:	data_out=16'h8001;
17'h15e9c:	data_out=16'h6;
17'h15e9d:	data_out=16'h1;
17'h15e9e:	data_out=16'h2;
17'h15e9f:	data_out=16'h1;
17'h15ea0:	data_out=16'h2;
17'h15ea1:	data_out=16'h8007;
17'h15ea2:	data_out=16'h3;
17'h15ea3:	data_out=16'h9;
17'h15ea4:	data_out=16'h4;
17'h15ea5:	data_out=16'h3;
17'h15ea6:	data_out=16'h8001;
17'h15ea7:	data_out=16'h8008;
17'h15ea8:	data_out=16'h8002;
17'h15ea9:	data_out=16'h8009;
17'h15eaa:	data_out=16'h5;
17'h15eab:	data_out=16'h8001;
17'h15eac:	data_out=16'h6;
17'h15ead:	data_out=16'h8003;
17'h15eae:	data_out=16'h7;
17'h15eaf:	data_out=16'h8009;
17'h15eb0:	data_out=16'h8008;
17'h15eb1:	data_out=16'h5;
17'h15eb2:	data_out=16'h8001;
17'h15eb3:	data_out=16'h8004;
17'h15eb4:	data_out=16'h8002;
17'h15eb5:	data_out=16'h5;
17'h15eb6:	data_out=16'h1;
17'h15eb7:	data_out=16'h8004;
17'h15eb8:	data_out=16'h1;
17'h15eb9:	data_out=16'h8000;
17'h15eba:	data_out=16'h4;
17'h15ebb:	data_out=16'h8002;
17'h15ebc:	data_out=16'h8009;
17'h15ebd:	data_out=16'h8003;
17'h15ebe:	data_out=16'h8;
17'h15ebf:	data_out=16'h2;
17'h15ec0:	data_out=16'h8001;
17'h15ec1:	data_out=16'h2;
17'h15ec2:	data_out=16'h2;
17'h15ec3:	data_out=16'h8006;
17'h15ec4:	data_out=16'h8004;
17'h15ec5:	data_out=16'h8009;
17'h15ec6:	data_out=16'h8005;
17'h15ec7:	data_out=16'h3;
17'h15ec8:	data_out=16'h8009;
17'h15ec9:	data_out=16'h8008;
17'h15eca:	data_out=16'h8007;
17'h15ecb:	data_out=16'h7;
17'h15ecc:	data_out=16'h8002;
17'h15ecd:	data_out=16'h8;
17'h15ece:	data_out=16'h7;
17'h15ecf:	data_out=16'h8001;
17'h15ed0:	data_out=16'h4;
17'h15ed1:	data_out=16'h8004;
17'h15ed2:	data_out=16'h4;
17'h15ed3:	data_out=16'h8007;
17'h15ed4:	data_out=16'h8008;
17'h15ed5:	data_out=16'h8004;
17'h15ed6:	data_out=16'h8002;
17'h15ed7:	data_out=16'h3;
17'h15ed8:	data_out=16'h5;
17'h15ed9:	data_out=16'h8007;
17'h15eda:	data_out=16'h8008;
17'h15edb:	data_out=16'h5;
17'h15edc:	data_out=16'h8001;
17'h15edd:	data_out=16'h8009;
17'h15ede:	data_out=16'h8002;
17'h15edf:	data_out=16'h8;
17'h15ee0:	data_out=16'h2;
17'h15ee1:	data_out=16'h8;
17'h15ee2:	data_out=16'h8007;
17'h15ee3:	data_out=16'h7;
17'h15ee4:	data_out=16'h8;
17'h15ee5:	data_out=16'h8003;
17'h15ee6:	data_out=16'h1;
17'h15ee7:	data_out=16'h9;
17'h15ee8:	data_out=16'h8002;
17'h15ee9:	data_out=16'h3;
17'h15eea:	data_out=16'h6;
17'h15eeb:	data_out=16'h5;
17'h15eec:	data_out=16'h2;
17'h15eed:	data_out=16'h4;
17'h15eee:	data_out=16'h8005;
17'h15eef:	data_out=16'h8003;
17'h15ef0:	data_out=16'h9;
17'h15ef1:	data_out=16'h8;
17'h15ef2:	data_out=16'h8001;
17'h15ef3:	data_out=16'h8008;
17'h15ef4:	data_out=16'h8005;
17'h15ef5:	data_out=16'h6;
17'h15ef6:	data_out=16'h4;
17'h15ef7:	data_out=16'h9;
17'h15ef8:	data_out=16'h9;
17'h15ef9:	data_out=16'h4;
17'h15efa:	data_out=16'h5;
17'h15efb:	data_out=16'h8001;
17'h15efc:	data_out=16'h4;
17'h15efd:	data_out=16'h8007;
17'h15efe:	data_out=16'h8002;
17'h15eff:	data_out=16'h8003;
17'h15f00:	data_out=16'h800f;
17'h15f01:	data_out=16'h8002;
17'h15f02:	data_out=16'h8009;
17'h15f03:	data_out=16'h8017;
17'h15f04:	data_out=16'h8003;
17'h15f05:	data_out=16'h1f;
17'h15f06:	data_out=16'h27;
17'h15f07:	data_out=16'h8005;
17'h15f08:	data_out=16'ha;
17'h15f09:	data_out=16'h1d;
17'h15f0a:	data_out=16'h4;
17'h15f0b:	data_out=16'h20;
17'h15f0c:	data_out=16'h800f;
17'h15f0d:	data_out=16'h801a;
17'h15f0e:	data_out=16'h1;
17'h15f0f:	data_out=16'h7;
17'h15f10:	data_out=16'h8010;
17'h15f11:	data_out=16'h3;
17'h15f12:	data_out=16'h800b;
17'h15f13:	data_out=16'h8007;
17'h15f14:	data_out=16'h8007;
17'h15f15:	data_out=16'h800b;
17'h15f16:	data_out=16'h800a;
17'h15f17:	data_out=16'h8008;
17'h15f18:	data_out=16'h8007;
17'h15f19:	data_out=16'h8007;
17'h15f1a:	data_out=16'h800c;
17'h15f1b:	data_out=16'h8005;
17'h15f1c:	data_out=16'h0;
17'h15f1d:	data_out=16'h8015;
17'h15f1e:	data_out=16'h800a;
17'h15f1f:	data_out=16'h10;
17'h15f20:	data_out=16'h8009;
17'h15f21:	data_out=16'h3;
17'h15f22:	data_out=16'h8010;
17'h15f23:	data_out=16'h8002;
17'h15f24:	data_out=16'h800b;
17'h15f25:	data_out=16'h8007;
17'h15f26:	data_out=16'h1a;
17'h15f27:	data_out=16'h800e;
17'h15f28:	data_out=16'h2;
17'h15f29:	data_out=16'h8005;
17'h15f2a:	data_out=16'h8006;
17'h15f2b:	data_out=16'hc;
17'h15f2c:	data_out=16'h8009;
17'h15f2d:	data_out=16'h8004;
17'h15f2e:	data_out=16'h8008;
17'h15f2f:	data_out=16'h8007;
17'h15f30:	data_out=16'h9;
17'h15f31:	data_out=16'h800f;
17'h15f32:	data_out=16'h7;
17'h15f33:	data_out=16'h800e;
17'h15f34:	data_out=16'h800d;
17'h15f35:	data_out=16'h10;
17'h15f36:	data_out=16'h1a;
17'h15f37:	data_out=16'h0;
17'h15f38:	data_out=16'h14;
17'h15f39:	data_out=16'he;
17'h15f3a:	data_out=16'h8019;
17'h15f3b:	data_out=16'hc;
17'h15f3c:	data_out=16'h3;
17'h15f3d:	data_out=16'h8;
17'h15f3e:	data_out=16'h7;
17'h15f3f:	data_out=16'hf;
17'h15f40:	data_out=16'h800b;
17'h15f41:	data_out=16'h12;
17'h15f42:	data_out=16'h800d;
17'h15f43:	data_out=16'h26;
17'h15f44:	data_out=16'h9;
17'h15f45:	data_out=16'h8002;
17'h15f46:	data_out=16'h6;
17'h15f47:	data_out=16'h8014;
17'h15f48:	data_out=16'h800f;
17'h15f49:	data_out=16'h8004;
17'h15f4a:	data_out=16'h800e;
17'h15f4b:	data_out=16'h8022;
17'h15f4c:	data_out=16'h801e;
17'h15f4d:	data_out=16'h8010;
17'h15f4e:	data_out=16'h8008;
17'h15f4f:	data_out=16'h800c;
17'h15f50:	data_out=16'h8016;
17'h15f51:	data_out=16'h3;
17'h15f52:	data_out=16'h8006;
17'h15f53:	data_out=16'h8024;
17'h15f54:	data_out=16'h8002;
17'h15f55:	data_out=16'h1e;
17'h15f56:	data_out=16'h4;
17'h15f57:	data_out=16'h8001;
17'h15f58:	data_out=16'h14;
17'h15f59:	data_out=16'hc;
17'h15f5a:	data_out=16'h800a;
17'h15f5b:	data_out=16'h1d;
17'h15f5c:	data_out=16'h3;
17'h15f5d:	data_out=16'h8008;
17'h15f5e:	data_out=16'h6;
17'h15f5f:	data_out=16'h8014;
17'h15f60:	data_out=16'ha;
17'h15f61:	data_out=16'h2;
17'h15f62:	data_out=16'h1a;
17'h15f63:	data_out=16'h800f;
17'h15f64:	data_out=16'h3;
17'h15f65:	data_out=16'h5;
17'h15f66:	data_out=16'h7;
17'h15f67:	data_out=16'h8011;
17'h15f68:	data_out=16'h5;
17'h15f69:	data_out=16'h10;
17'h15f6a:	data_out=16'h8;
17'h15f6b:	data_out=16'hc;
17'h15f6c:	data_out=16'h801b;
17'h15f6d:	data_out=16'h800e;
17'h15f6e:	data_out=16'h9;
17'h15f6f:	data_out=16'h7;
17'h15f70:	data_out=16'h4;
17'h15f71:	data_out=16'h8011;
17'h15f72:	data_out=16'h1;
17'h15f73:	data_out=16'hd;
17'h15f74:	data_out=16'h8001;
17'h15f75:	data_out=16'h24;
17'h15f76:	data_out=16'hc;
17'h15f77:	data_out=16'h8004;
17'h15f78:	data_out=16'h23;
17'h15f79:	data_out=16'h8002;
17'h15f7a:	data_out=16'h800c;
17'h15f7b:	data_out=16'h2;
17'h15f7c:	data_out=16'h11;
17'h15f7d:	data_out=16'h3f;
17'h15f7e:	data_out=16'h16;
17'h15f7f:	data_out=16'h800a;
17'h15f80:	data_out=16'h5d;
17'h15f81:	data_out=16'h8008;
17'h15f82:	data_out=16'h183;
17'h15f83:	data_out=16'h80df;
17'h15f84:	data_out=16'h81c8;
17'h15f85:	data_out=16'h810e;
17'h15f86:	data_out=16'h82e0;
17'h15f87:	data_out=16'h81ff;
17'h15f88:	data_out=16'h80;
17'h15f89:	data_out=16'h81d8;
17'h15f8a:	data_out=16'h9d;
17'h15f8b:	data_out=16'h81b9;
17'h15f8c:	data_out=16'h8094;
17'h15f8d:	data_out=16'h80b0;
17'h15f8e:	data_out=16'h8082;
17'h15f8f:	data_out=16'h8011;
17'h15f90:	data_out=16'h8080;
17'h15f91:	data_out=16'h81d3;
17'h15f92:	data_out=16'h12c;
17'h15f93:	data_out=16'h81f1;
17'h15f94:	data_out=16'h92;
17'h15f95:	data_out=16'h80dc;
17'h15f96:	data_out=16'h80f1;
17'h15f97:	data_out=16'h8003;
17'h15f98:	data_out=16'h8065;
17'h15f99:	data_out=16'h8277;
17'h15f9a:	data_out=16'h8295;
17'h15f9b:	data_out=16'h80f6;
17'h15f9c:	data_out=16'h8001;
17'h15f9d:	data_out=16'h17f;
17'h15f9e:	data_out=16'h10c;
17'h15f9f:	data_out=16'h8110;
17'h15fa0:	data_out=16'h283;
17'h15fa1:	data_out=16'h808c;
17'h15fa2:	data_out=16'h23;
17'h15fa3:	data_out=16'h5b;
17'h15fa4:	data_out=16'h5d;
17'h15fa5:	data_out=16'h80f1;
17'h15fa6:	data_out=16'h8189;
17'h15fa7:	data_out=16'h1ce;
17'h15fa8:	data_out=16'h8080;
17'h15fa9:	data_out=16'h8139;
17'h15faa:	data_out=16'h36;
17'h15fab:	data_out=16'h80b6;
17'h15fac:	data_out=16'h80c1;
17'h15fad:	data_out=16'h8226;
17'h15fae:	data_out=16'h101;
17'h15faf:	data_out=16'hc;
17'h15fb0:	data_out=16'h82aa;
17'h15fb1:	data_out=16'h8128;
17'h15fb2:	data_out=16'h82d8;
17'h15fb3:	data_out=16'hda;
17'h15fb4:	data_out=16'h8260;
17'h15fb5:	data_out=16'h815e;
17'h15fb6:	data_out=16'h226;
17'h15fb7:	data_out=16'h174;
17'h15fb8:	data_out=16'h8159;
17'h15fb9:	data_out=16'h8086;
17'h15fba:	data_out=16'h10d;
17'h15fbb:	data_out=16'h80ca;
17'h15fbc:	data_out=16'h216;
17'h15fbd:	data_out=16'h815d;
17'h15fbe:	data_out=16'h8081;
17'h15fbf:	data_out=16'h820f;
17'h15fc0:	data_out=16'h80e2;
17'h15fc1:	data_out=16'h223;
17'h15fc2:	data_out=16'h8109;
17'h15fc3:	data_out=16'h825c;
17'h15fc4:	data_out=16'h8113;
17'h15fc5:	data_out=16'h80df;
17'h15fc6:	data_out=16'h14d;
17'h15fc7:	data_out=16'h8028;
17'h15fc8:	data_out=16'hba;
17'h15fc9:	data_out=16'h80e0;
17'h15fca:	data_out=16'h8124;
17'h15fcb:	data_out=16'h8082;
17'h15fcc:	data_out=16'h8153;
17'h15fcd:	data_out=16'h6b;
17'h15fce:	data_out=16'h8007;
17'h15fcf:	data_out=16'h8134;
17'h15fd0:	data_out=16'h80dd;
17'h15fd1:	data_out=16'h819c;
17'h15fd2:	data_out=16'h11;
17'h15fd3:	data_out=16'h190;
17'h15fd4:	data_out=16'hb0;
17'h15fd5:	data_out=16'h34;
17'h15fd6:	data_out=16'h5c;
17'h15fd7:	data_out=16'h69;
17'h15fd8:	data_out=16'h125;
17'h15fd9:	data_out=16'h801e;
17'h15fda:	data_out=16'ha3;
17'h15fdb:	data_out=16'h816e;
17'h15fdc:	data_out=16'h8032;
17'h15fdd:	data_out=16'h5c;
17'h15fde:	data_out=16'h8046;
17'h15fdf:	data_out=16'hb4;
17'h15fe0:	data_out=16'h81fc;
17'h15fe1:	data_out=16'h8174;
17'h15fe2:	data_out=16'h806f;
17'h15fe3:	data_out=16'hd6;
17'h15fe4:	data_out=16'h8286;
17'h15fe5:	data_out=16'h82bf;
17'h15fe6:	data_out=16'h832b;
17'h15fe7:	data_out=16'h15e;
17'h15fe8:	data_out=16'h8084;
17'h15fe9:	data_out=16'h155;
17'h15fea:	data_out=16'h808d;
17'h15feb:	data_out=16'h8218;
17'h15fec:	data_out=16'h312;
17'h15fed:	data_out=16'hd8;
17'h15fee:	data_out=16'h8088;
17'h15fef:	data_out=16'h8164;
17'h15ff0:	data_out=16'h8085;
17'h15ff1:	data_out=16'h8026;
17'h15ff2:	data_out=16'h82c2;
17'h15ff3:	data_out=16'h82b3;
17'h15ff4:	data_out=16'h82a3;
17'h15ff5:	data_out=16'h8163;
17'h15ff6:	data_out=16'h816a;
17'h15ff7:	data_out=16'h826b;
17'h15ff8:	data_out=16'h836e;
17'h15ff9:	data_out=16'h75;
17'h15ffa:	data_out=16'hba;
17'h15ffb:	data_out=16'h8084;
17'h15ffc:	data_out=16'h8049;
17'h15ffd:	data_out=16'h8324;
17'h15ffe:	data_out=16'h8297;
17'h15fff:	data_out=16'h8149;
17'h16000:	data_out=16'h82f1;
17'h16001:	data_out=16'h816d;
17'h16002:	data_out=16'h144;
17'h16003:	data_out=16'h85d4;
17'h16004:	data_out=16'h8a00;
17'h16005:	data_out=16'h8a00;
17'h16006:	data_out=16'h8a00;
17'h16007:	data_out=16'h8a00;
17'h16008:	data_out=16'ha00;
17'h16009:	data_out=16'h8207;
17'h1600a:	data_out=16'h896d;
17'h1600b:	data_out=16'ha00;
17'h1600c:	data_out=16'h896a;
17'h1600d:	data_out=16'hf5;
17'h1600e:	data_out=16'h83d7;
17'h1600f:	data_out=16'h160;
17'h16010:	data_out=16'h9c7;
17'h16011:	data_out=16'h8a00;
17'h16012:	data_out=16'h838;
17'h16013:	data_out=16'h85f3;
17'h16014:	data_out=16'h61f;
17'h16015:	data_out=16'h880b;
17'h16016:	data_out=16'h8a00;
17'h16017:	data_out=16'h613;
17'h16018:	data_out=16'h80b2;
17'h16019:	data_out=16'h89a4;
17'h1601a:	data_out=16'h8a00;
17'h1601b:	data_out=16'ha00;
17'h1601c:	data_out=16'h89b6;
17'h1601d:	data_out=16'h838d;
17'h1601e:	data_out=16'h57a;
17'h1601f:	data_out=16'h8a00;
17'h16020:	data_out=16'h6f3;
17'h16021:	data_out=16'h83c3;
17'h16022:	data_out=16'h557;
17'h16023:	data_out=16'h85d9;
17'h16024:	data_out=16'h85e5;
17'h16025:	data_out=16'h824f;
17'h16026:	data_out=16'h820b;
17'h16027:	data_out=16'h3f;
17'h16028:	data_out=16'h83b5;
17'h16029:	data_out=16'h5ef;
17'h1602a:	data_out=16'h64e;
17'h1602b:	data_out=16'h84a;
17'h1602c:	data_out=16'h8a00;
17'h1602d:	data_out=16'h4aa;
17'h1602e:	data_out=16'h9d8;
17'h1602f:	data_out=16'h9fc;
17'h16030:	data_out=16'h8a00;
17'h16031:	data_out=16'h8644;
17'h16032:	data_out=16'h8a00;
17'h16033:	data_out=16'h68c;
17'h16034:	data_out=16'h89ff;
17'h16035:	data_out=16'h8a00;
17'h16036:	data_out=16'ha00;
17'h16037:	data_out=16'h178;
17'h16038:	data_out=16'h89ff;
17'h16039:	data_out=16'h71c;
17'h1603a:	data_out=16'h200;
17'h1603b:	data_out=16'h8a00;
17'h1603c:	data_out=16'h9e2;
17'h1603d:	data_out=16'h8a00;
17'h1603e:	data_out=16'h83b5;
17'h1603f:	data_out=16'h8a00;
17'h16040:	data_out=16'h8a00;
17'h16041:	data_out=16'ha00;
17'h16042:	data_out=16'h7e5;
17'h16043:	data_out=16'h8a00;
17'h16044:	data_out=16'h8a00;
17'h16045:	data_out=16'h8859;
17'h16046:	data_out=16'h9d2;
17'h16047:	data_out=16'h88d0;
17'h16048:	data_out=16'h9e7;
17'h16049:	data_out=16'h8404;
17'h1604a:	data_out=16'h85d9;
17'h1604b:	data_out=16'h893;
17'h1604c:	data_out=16'h8427;
17'h1604d:	data_out=16'h630;
17'h1604e:	data_out=16'h6a9;
17'h1604f:	data_out=16'h8765;
17'h16050:	data_out=16'h8a00;
17'h16051:	data_out=16'h8a00;
17'h16052:	data_out=16'h8a00;
17'h16053:	data_out=16'h909;
17'h16054:	data_out=16'h9ff;
17'h16055:	data_out=16'h808a;
17'h16056:	data_out=16'h8a00;
17'h16057:	data_out=16'h8a00;
17'h16058:	data_out=16'h8027;
17'h16059:	data_out=16'h8a00;
17'h1605a:	data_out=16'ha00;
17'h1605b:	data_out=16'h8a00;
17'h1605c:	data_out=16'h8026;
17'h1605d:	data_out=16'h27e;
17'h1605e:	data_out=16'h9da;
17'h1605f:	data_out=16'h52a;
17'h16060:	data_out=16'h8a00;
17'h16061:	data_out=16'h8a00;
17'h16062:	data_out=16'h730;
17'h16063:	data_out=16'h72b;
17'h16064:	data_out=16'h89fd;
17'h16065:	data_out=16'h8a00;
17'h16066:	data_out=16'h8a00;
17'h16067:	data_out=16'h8c6;
17'h16068:	data_out=16'h83bc;
17'h16069:	data_out=16'ha00;
17'h1606a:	data_out=16'h83e7;
17'h1606b:	data_out=16'h8a00;
17'h1606c:	data_out=16'h14;
17'h1606d:	data_out=16'h6ef;
17'h1606e:	data_out=16'h83e7;
17'h1606f:	data_out=16'h8a00;
17'h16070:	data_out=16'h83de;
17'h16071:	data_out=16'h872f;
17'h16072:	data_out=16'h8a00;
17'h16073:	data_out=16'h8a00;
17'h16074:	data_out=16'h8a00;
17'h16075:	data_out=16'h8835;
17'h16076:	data_out=16'h814b;
17'h16077:	data_out=16'h8a00;
17'h16078:	data_out=16'h8a00;
17'h16079:	data_out=16'h8f7;
17'h1607a:	data_out=16'h75e;
17'h1607b:	data_out=16'h83b5;
17'h1607c:	data_out=16'hd0;
17'h1607d:	data_out=16'h8a00;
17'h1607e:	data_out=16'h8199;
17'h1607f:	data_out=16'h8a00;
17'h16080:	data_out=16'h89f7;
17'h16081:	data_out=16'h8a00;
17'h16082:	data_out=16'h55a;
17'h16083:	data_out=16'h8402;
17'h16084:	data_out=16'h8a00;
17'h16085:	data_out=16'h8a00;
17'h16086:	data_out=16'h8a00;
17'h16087:	data_out=16'h8a00;
17'h16088:	data_out=16'ha00;
17'h16089:	data_out=16'h204;
17'h1608a:	data_out=16'h8a00;
17'h1608b:	data_out=16'ha00;
17'h1608c:	data_out=16'h8992;
17'h1608d:	data_out=16'h31a;
17'h1608e:	data_out=16'h861d;
17'h1608f:	data_out=16'h35d;
17'h16090:	data_out=16'h9f7;
17'h16091:	data_out=16'h8a00;
17'h16092:	data_out=16'h9ff;
17'h16093:	data_out=16'h8699;
17'h16094:	data_out=16'h9fd;
17'h16095:	data_out=16'h8a00;
17'h16096:	data_out=16'h8a00;
17'h16097:	data_out=16'h9fd;
17'h16098:	data_out=16'h82ff;
17'h16099:	data_out=16'h8945;
17'h1609a:	data_out=16'h8a00;
17'h1609b:	data_out=16'ha00;
17'h1609c:	data_out=16'h87de;
17'h1609d:	data_out=16'h8a00;
17'h1609e:	data_out=16'h984;
17'h1609f:	data_out=16'h8a00;
17'h160a0:	data_out=16'h8156;
17'h160a1:	data_out=16'h85e1;
17'h160a2:	data_out=16'h990;
17'h160a3:	data_out=16'h89ff;
17'h160a4:	data_out=16'h89ff;
17'h160a5:	data_out=16'h802b;
17'h160a6:	data_out=16'h91b;
17'h160a7:	data_out=16'h8916;
17'h160a8:	data_out=16'h8590;
17'h160a9:	data_out=16'ha00;
17'h160aa:	data_out=16'h8c2;
17'h160ab:	data_out=16'ha00;
17'h160ac:	data_out=16'h8a00;
17'h160ad:	data_out=16'h86e;
17'h160ae:	data_out=16'h984;
17'h160af:	data_out=16'h9a3;
17'h160b0:	data_out=16'h8a00;
17'h160b1:	data_out=16'h8a00;
17'h160b2:	data_out=16'h8a00;
17'h160b3:	data_out=16'ha00;
17'h160b4:	data_out=16'h8a00;
17'h160b5:	data_out=16'h8a00;
17'h160b6:	data_out=16'h9fe;
17'h160b7:	data_out=16'h65b;
17'h160b8:	data_out=16'h89f2;
17'h160b9:	data_out=16'ha00;
17'h160ba:	data_out=16'h841c;
17'h160bb:	data_out=16'h8a00;
17'h160bc:	data_out=16'ha00;
17'h160bd:	data_out=16'h8a00;
17'h160be:	data_out=16'h858f;
17'h160bf:	data_out=16'h8a00;
17'h160c0:	data_out=16'h8a00;
17'h160c1:	data_out=16'ha00;
17'h160c2:	data_out=16'h9a6;
17'h160c3:	data_out=16'h888e;
17'h160c4:	data_out=16'h8a00;
17'h160c5:	data_out=16'h8a00;
17'h160c6:	data_out=16'ha00;
17'h160c7:	data_out=16'h89fe;
17'h160c8:	data_out=16'h963;
17'h160c9:	data_out=16'h82aa;
17'h160ca:	data_out=16'h85a3;
17'h160cb:	data_out=16'h709;
17'h160cc:	data_out=16'h8a00;
17'h160cd:	data_out=16'h986;
17'h160ce:	data_out=16'ha00;
17'h160cf:	data_out=16'h8a00;
17'h160d0:	data_out=16'h8a00;
17'h160d1:	data_out=16'h89de;
17'h160d2:	data_out=16'h8a00;
17'h160d3:	data_out=16'h9a6;
17'h160d4:	data_out=16'h94c;
17'h160d5:	data_out=16'h961;
17'h160d6:	data_out=16'h89fc;
17'h160d7:	data_out=16'h8a00;
17'h160d8:	data_out=16'ha00;
17'h160d9:	data_out=16'h8a00;
17'h160da:	data_out=16'ha00;
17'h160db:	data_out=16'h8a00;
17'h160dc:	data_out=16'h8206;
17'h160dd:	data_out=16'h854d;
17'h160de:	data_out=16'h933;
17'h160df:	data_out=16'h36b;
17'h160e0:	data_out=16'h8a00;
17'h160e1:	data_out=16'h8a00;
17'h160e2:	data_out=16'h9fd;
17'h160e3:	data_out=16'ha00;
17'h160e4:	data_out=16'h8a00;
17'h160e5:	data_out=16'h8a00;
17'h160e6:	data_out=16'h89e8;
17'h160e7:	data_out=16'h8bb;
17'h160e8:	data_out=16'h85be;
17'h160e9:	data_out=16'ha00;
17'h160ea:	data_out=16'h8647;
17'h160eb:	data_out=16'h8a00;
17'h160ec:	data_out=16'h8a00;
17'h160ed:	data_out=16'ha00;
17'h160ee:	data_out=16'h8646;
17'h160ef:	data_out=16'h8a00;
17'h160f0:	data_out=16'h8630;
17'h160f1:	data_out=16'h8905;
17'h160f2:	data_out=16'h8a00;
17'h160f3:	data_out=16'h8a00;
17'h160f4:	data_out=16'h8a00;
17'h160f5:	data_out=16'h89ff;
17'h160f6:	data_out=16'h280;
17'h160f7:	data_out=16'h89d5;
17'h160f8:	data_out=16'h89fd;
17'h160f9:	data_out=16'ha00;
17'h160fa:	data_out=16'h9ff;
17'h160fb:	data_out=16'h858e;
17'h160fc:	data_out=16'h820d;
17'h160fd:	data_out=16'h8a00;
17'h160fe:	data_out=16'h9af;
17'h160ff:	data_out=16'h8a00;
17'h16100:	data_out=16'h89fa;
17'h16101:	data_out=16'h8a00;
17'h16102:	data_out=16'h9ef;
17'h16103:	data_out=16'h19b;
17'h16104:	data_out=16'h8a00;
17'h16105:	data_out=16'h89ff;
17'h16106:	data_out=16'h8a00;
17'h16107:	data_out=16'h8a00;
17'h16108:	data_out=16'ha00;
17'h16109:	data_out=16'h8058;
17'h1610a:	data_out=16'h8a00;
17'h1610b:	data_out=16'ha00;
17'h1610c:	data_out=16'h89f9;
17'h1610d:	data_out=16'h741;
17'h1610e:	data_out=16'h8731;
17'h1610f:	data_out=16'h881;
17'h16110:	data_out=16'h9d5;
17'h16111:	data_out=16'h89e2;
17'h16112:	data_out=16'h9f4;
17'h16113:	data_out=16'h870e;
17'h16114:	data_out=16'h9fa;
17'h16115:	data_out=16'h8a00;
17'h16116:	data_out=16'h8a00;
17'h16117:	data_out=16'h9f9;
17'h16118:	data_out=16'h840d;
17'h16119:	data_out=16'h876e;
17'h1611a:	data_out=16'h8a00;
17'h1611b:	data_out=16'ha00;
17'h1611c:	data_out=16'h84fd;
17'h1611d:	data_out=16'h8a00;
17'h1611e:	data_out=16'h94e;
17'h1611f:	data_out=16'h8a00;
17'h16120:	data_out=16'h6c0;
17'h16121:	data_out=16'h86cc;
17'h16122:	data_out=16'h542;
17'h16123:	data_out=16'h89f8;
17'h16124:	data_out=16'h89f8;
17'h16125:	data_out=16'h833b;
17'h16126:	data_out=16'h805;
17'h16127:	data_out=16'h82bb;
17'h16128:	data_out=16'h861d;
17'h16129:	data_out=16'ha00;
17'h1612a:	data_out=16'h796;
17'h1612b:	data_out=16'h9ff;
17'h1612c:	data_out=16'h8a00;
17'h1612d:	data_out=16'h506;
17'h1612e:	data_out=16'h8e9;
17'h1612f:	data_out=16'h97a;
17'h16130:	data_out=16'h8a00;
17'h16131:	data_out=16'h89ff;
17'h16132:	data_out=16'h8a00;
17'h16133:	data_out=16'h9ff;
17'h16134:	data_out=16'h8a00;
17'h16135:	data_out=16'h8a00;
17'h16136:	data_out=16'h9f4;
17'h16137:	data_out=16'h9f5;
17'h16138:	data_out=16'h8879;
17'h16139:	data_out=16'ha00;
17'h1613a:	data_out=16'h8a00;
17'h1613b:	data_out=16'h8a00;
17'h1613c:	data_out=16'ha00;
17'h1613d:	data_out=16'h8a00;
17'h1613e:	data_out=16'h8619;
17'h1613f:	data_out=16'h89ff;
17'h16140:	data_out=16'h8a00;
17'h16141:	data_out=16'ha00;
17'h16142:	data_out=16'h7db;
17'h16143:	data_out=16'h852f;
17'h16144:	data_out=16'h89fe;
17'h16145:	data_out=16'h8a00;
17'h16146:	data_out=16'ha00;
17'h16147:	data_out=16'h8a00;
17'h16148:	data_out=16'h8b5;
17'h16149:	data_out=16'h84cf;
17'h1614a:	data_out=16'h81f8;
17'h1614b:	data_out=16'h9ae;
17'h1614c:	data_out=16'h8a00;
17'h1614d:	data_out=16'h605;
17'h1614e:	data_out=16'ha00;
17'h1614f:	data_out=16'h8a00;
17'h16150:	data_out=16'h8a00;
17'h16151:	data_out=16'h86dc;
17'h16152:	data_out=16'h8a00;
17'h16153:	data_out=16'h9e7;
17'h16154:	data_out=16'h822;
17'h16155:	data_out=16'h9a9;
17'h16156:	data_out=16'h89ec;
17'h16157:	data_out=16'h8a00;
17'h16158:	data_out=16'ha00;
17'h16159:	data_out=16'h8a00;
17'h1615a:	data_out=16'ha00;
17'h1615b:	data_out=16'h89ff;
17'h1615c:	data_out=16'ha00;
17'h1615d:	data_out=16'h8568;
17'h1615e:	data_out=16'h8eb;
17'h1615f:	data_out=16'h352;
17'h16160:	data_out=16'h8a00;
17'h16161:	data_out=16'h89ff;
17'h16162:	data_out=16'h9f9;
17'h16163:	data_out=16'h9fe;
17'h16164:	data_out=16'h89fe;
17'h16165:	data_out=16'h8a00;
17'h16166:	data_out=16'h8663;
17'h16167:	data_out=16'h767;
17'h16168:	data_out=16'h8688;
17'h16169:	data_out=16'ha00;
17'h1616a:	data_out=16'h877a;
17'h1616b:	data_out=16'h8a00;
17'h1616c:	data_out=16'h89ff;
17'h1616d:	data_out=16'h9fe;
17'h1616e:	data_out=16'h8779;
17'h1616f:	data_out=16'h8a00;
17'h16170:	data_out=16'h8752;
17'h16171:	data_out=16'h87d6;
17'h16172:	data_out=16'h8a00;
17'h16173:	data_out=16'h8a00;
17'h16174:	data_out=16'h8a00;
17'h16175:	data_out=16'h30;
17'h16176:	data_out=16'h9cf;
17'h16177:	data_out=16'h88cf;
17'h16178:	data_out=16'h88ec;
17'h16179:	data_out=16'ha00;
17'h1617a:	data_out=16'h9fb;
17'h1617b:	data_out=16'h8617;
17'h1617c:	data_out=16'h82eb;
17'h1617d:	data_out=16'h8a00;
17'h1617e:	data_out=16'h8db;
17'h1617f:	data_out=16'h8a00;
17'h16180:	data_out=16'h89fb;
17'h16181:	data_out=16'h892c;
17'h16182:	data_out=16'ha00;
17'h16183:	data_out=16'h85e;
17'h16184:	data_out=16'h89ff;
17'h16185:	data_out=16'h89fc;
17'h16186:	data_out=16'h8a00;
17'h16187:	data_out=16'h8a00;
17'h16188:	data_out=16'ha00;
17'h16189:	data_out=16'h8a00;
17'h1618a:	data_out=16'h8a00;
17'h1618b:	data_out=16'ha00;
17'h1618c:	data_out=16'h85f4;
17'h1618d:	data_out=16'h9fe;
17'h1618e:	data_out=16'h8775;
17'h1618f:	data_out=16'h83d;
17'h16190:	data_out=16'h9bc;
17'h16191:	data_out=16'h88d7;
17'h16192:	data_out=16'h9e9;
17'h16193:	data_out=16'h8a00;
17'h16194:	data_out=16'h9f4;
17'h16195:	data_out=16'h8a00;
17'h16196:	data_out=16'h8a00;
17'h16197:	data_out=16'h9f5;
17'h16198:	data_out=16'h824b;
17'h16199:	data_out=16'h887d;
17'h1619a:	data_out=16'h89fc;
17'h1619b:	data_out=16'ha00;
17'h1619c:	data_out=16'h1aa;
17'h1619d:	data_out=16'h881a;
17'h1619e:	data_out=16'h921;
17'h1619f:	data_out=16'h8a00;
17'h161a0:	data_out=16'h571;
17'h161a1:	data_out=16'h86e2;
17'h161a2:	data_out=16'h82a5;
17'h161a3:	data_out=16'h89fe;
17'h161a4:	data_out=16'h89fe;
17'h161a5:	data_out=16'h8a00;
17'h161a6:	data_out=16'h8f6;
17'h161a7:	data_out=16'h648;
17'h161a8:	data_out=16'h85c4;
17'h161a9:	data_out=16'ha00;
17'h161aa:	data_out=16'h602;
17'h161ab:	data_out=16'h9fd;
17'h161ac:	data_out=16'h8a00;
17'h161ad:	data_out=16'h8054;
17'h161ae:	data_out=16'h7c5;
17'h161af:	data_out=16'h94d;
17'h161b0:	data_out=16'h89ff;
17'h161b1:	data_out=16'h89fc;
17'h161b2:	data_out=16'h89fe;
17'h161b3:	data_out=16'h9fd;
17'h161b4:	data_out=16'h8a00;
17'h161b5:	data_out=16'h870e;
17'h161b6:	data_out=16'h9f8;
17'h161b7:	data_out=16'h9ff;
17'h161b8:	data_out=16'h85f9;
17'h161b9:	data_out=16'ha00;
17'h161ba:	data_out=16'h8a00;
17'h161bb:	data_out=16'h89fd;
17'h161bc:	data_out=16'ha00;
17'h161bd:	data_out=16'h8a00;
17'h161be:	data_out=16'h85bc;
17'h161bf:	data_out=16'h89fc;
17'h161c0:	data_out=16'h8a00;
17'h161c1:	data_out=16'ha00;
17'h161c2:	data_out=16'h546;
17'h161c3:	data_out=16'h83a4;
17'h161c4:	data_out=16'h89fc;
17'h161c5:	data_out=16'h8a00;
17'h161c6:	data_out=16'ha00;
17'h161c7:	data_out=16'h8a00;
17'h161c8:	data_out=16'h679;
17'h161c9:	data_out=16'h8a00;
17'h161ca:	data_out=16'h667;
17'h161cb:	data_out=16'h800;
17'h161cc:	data_out=16'h8a00;
17'h161cd:	data_out=16'h8185;
17'h161ce:	data_out=16'ha00;
17'h161cf:	data_out=16'h8a00;
17'h161d0:	data_out=16'h8a00;
17'h161d1:	data_out=16'h81db;
17'h161d2:	data_out=16'h8a00;
17'h161d3:	data_out=16'h9e9;
17'h161d4:	data_out=16'h6d8;
17'h161d5:	data_out=16'h9a7;
17'h161d6:	data_out=16'h89b4;
17'h161d7:	data_out=16'h8a00;
17'h161d8:	data_out=16'ha00;
17'h161d9:	data_out=16'h8a00;
17'h161da:	data_out=16'ha00;
17'h161db:	data_out=16'h89fc;
17'h161dc:	data_out=16'ha00;
17'h161dd:	data_out=16'h13f;
17'h161de:	data_out=16'h871;
17'h161df:	data_out=16'h73c;
17'h161e0:	data_out=16'h8a00;
17'h161e1:	data_out=16'h89fc;
17'h161e2:	data_out=16'h9ec;
17'h161e3:	data_out=16'h9fd;
17'h161e4:	data_out=16'h89fc;
17'h161e5:	data_out=16'h8a00;
17'h161e6:	data_out=16'h89fe;
17'h161e7:	data_out=16'h500;
17'h161e8:	data_out=16'h867e;
17'h161e9:	data_out=16'ha00;
17'h161ea:	data_out=16'h87e2;
17'h161eb:	data_out=16'h89ff;
17'h161ec:	data_out=16'h8a00;
17'h161ed:	data_out=16'h9fc;
17'h161ee:	data_out=16'h87e1;
17'h161ef:	data_out=16'h89fe;
17'h161f0:	data_out=16'h87a3;
17'h161f1:	data_out=16'h82b0;
17'h161f2:	data_out=16'h8a00;
17'h161f3:	data_out=16'h8a00;
17'h161f4:	data_out=16'h89fd;
17'h161f5:	data_out=16'ha00;
17'h161f6:	data_out=16'h9ad;
17'h161f7:	data_out=16'h8922;
17'h161f8:	data_out=16'h86b8;
17'h161f9:	data_out=16'ha00;
17'h161fa:	data_out=16'h9f9;
17'h161fb:	data_out=16'h85b8;
17'h161fc:	data_out=16'h8054;
17'h161fd:	data_out=16'h89fe;
17'h161fe:	data_out=16'h487;
17'h161ff:	data_out=16'h8a00;
17'h16200:	data_out=16'h89f8;
17'h16201:	data_out=16'h89fc;
17'h16202:	data_out=16'h9fe;
17'h16203:	data_out=16'h9dc;
17'h16204:	data_out=16'h89fe;
17'h16205:	data_out=16'h8822;
17'h16206:	data_out=16'h89ff;
17'h16207:	data_out=16'h8a00;
17'h16208:	data_out=16'ha00;
17'h16209:	data_out=16'h8a00;
17'h1620a:	data_out=16'h89ff;
17'h1620b:	data_out=16'h9fe;
17'h1620c:	data_out=16'h8153;
17'h1620d:	data_out=16'h9fb;
17'h1620e:	data_out=16'h844b;
17'h1620f:	data_out=16'h8c8;
17'h16210:	data_out=16'h918;
17'h16211:	data_out=16'h85dd;
17'h16212:	data_out=16'h9c6;
17'h16213:	data_out=16'h885f;
17'h16214:	data_out=16'h9f4;
17'h16215:	data_out=16'h8a00;
17'h16216:	data_out=16'h8a00;
17'h16217:	data_out=16'h9f8;
17'h16218:	data_out=16'h82a8;
17'h16219:	data_out=16'h8928;
17'h1621a:	data_out=16'h895c;
17'h1621b:	data_out=16'ha00;
17'h1621c:	data_out=16'ha00;
17'h1621d:	data_out=16'h89f9;
17'h1621e:	data_out=16'h978;
17'h1621f:	data_out=16'h8099;
17'h16220:	data_out=16'h6a2;
17'h16221:	data_out=16'h8381;
17'h16222:	data_out=16'h89fc;
17'h16223:	data_out=16'h89fe;
17'h16224:	data_out=16'h89fe;
17'h16225:	data_out=16'h8a00;
17'h16226:	data_out=16'h82b;
17'h16227:	data_out=16'h7a6;
17'h16228:	data_out=16'h81bf;
17'h16229:	data_out=16'h9ff;
17'h1622a:	data_out=16'h38b;
17'h1622b:	data_out=16'h9fb;
17'h1622c:	data_out=16'h8a00;
17'h1622d:	data_out=16'h84d8;
17'h1622e:	data_out=16'h6d5;
17'h1622f:	data_out=16'h9e0;
17'h16230:	data_out=16'h89f7;
17'h16231:	data_out=16'h885a;
17'h16232:	data_out=16'h89f3;
17'h16233:	data_out=16'h9fe;
17'h16234:	data_out=16'h8a00;
17'h16235:	data_out=16'h803b;
17'h16236:	data_out=16'h9f9;
17'h16237:	data_out=16'h9ff;
17'h16238:	data_out=16'h261;
17'h16239:	data_out=16'h9fe;
17'h1623a:	data_out=16'h8a00;
17'h1623b:	data_out=16'h87d9;
17'h1623c:	data_out=16'ha00;
17'h1623d:	data_out=16'h8a00;
17'h1623e:	data_out=16'h81af;
17'h1623f:	data_out=16'h8834;
17'h16240:	data_out=16'h89ff;
17'h16241:	data_out=16'ha00;
17'h16242:	data_out=16'h89f6;
17'h16243:	data_out=16'h9f3;
17'h16244:	data_out=16'h889b;
17'h16245:	data_out=16'h8a00;
17'h16246:	data_out=16'ha00;
17'h16247:	data_out=16'h8a00;
17'h16248:	data_out=16'h2d8;
17'h16249:	data_out=16'h8a00;
17'h1624a:	data_out=16'h9d9;
17'h1624b:	data_out=16'h440;
17'h1624c:	data_out=16'h8a00;
17'h1624d:	data_out=16'h89fe;
17'h1624e:	data_out=16'ha00;
17'h1624f:	data_out=16'h8a00;
17'h16250:	data_out=16'h89b7;
17'h16251:	data_out=16'h9f2;
17'h16252:	data_out=16'h8a00;
17'h16253:	data_out=16'ha00;
17'h16254:	data_out=16'h6f1;
17'h16255:	data_out=16'h9e8;
17'h16256:	data_out=16'h88c2;
17'h16257:	data_out=16'h8a00;
17'h16258:	data_out=16'ha00;
17'h16259:	data_out=16'h8a00;
17'h1625a:	data_out=16'ha00;
17'h1625b:	data_out=16'h8966;
17'h1625c:	data_out=16'ha00;
17'h1625d:	data_out=16'h8285;
17'h1625e:	data_out=16'h9cb;
17'h1625f:	data_out=16'h6b2;
17'h16260:	data_out=16'h89ff;
17'h16261:	data_out=16'h898d;
17'h16262:	data_out=16'h9e5;
17'h16263:	data_out=16'h9ff;
17'h16264:	data_out=16'h8a00;
17'h16265:	data_out=16'h89fe;
17'h16266:	data_out=16'h89e5;
17'h16267:	data_out=16'h339;
17'h16268:	data_out=16'h82ed;
17'h16269:	data_out=16'h9fd;
17'h1626a:	data_out=16'h84da;
17'h1626b:	data_out=16'h89fe;
17'h1626c:	data_out=16'h8a00;
17'h1626d:	data_out=16'h9fe;
17'h1626e:	data_out=16'h84d8;
17'h1626f:	data_out=16'h89f4;
17'h16270:	data_out=16'h8486;
17'h16271:	data_out=16'h8188;
17'h16272:	data_out=16'h8a00;
17'h16273:	data_out=16'h89fc;
17'h16274:	data_out=16'h89f3;
17'h16275:	data_out=16'ha00;
17'h16276:	data_out=16'h961;
17'h16277:	data_out=16'h86aa;
17'h16278:	data_out=16'h63d;
17'h16279:	data_out=16'h9ff;
17'h1627a:	data_out=16'h9fb;
17'h1627b:	data_out=16'h81a8;
17'h1627c:	data_out=16'hb5;
17'h1627d:	data_out=16'h89fd;
17'h1627e:	data_out=16'h129;
17'h1627f:	data_out=16'h89ff;
17'h16280:	data_out=16'h89f0;
17'h16281:	data_out=16'h89b5;
17'h16282:	data_out=16'ha00;
17'h16283:	data_out=16'h9a6;
17'h16284:	data_out=16'h89f0;
17'h16285:	data_out=16'h83a7;
17'h16286:	data_out=16'h89ff;
17'h16287:	data_out=16'h8a00;
17'h16288:	data_out=16'ha00;
17'h16289:	data_out=16'h8a00;
17'h1628a:	data_out=16'h89e4;
17'h1628b:	data_out=16'h9af;
17'h1628c:	data_out=16'h6b4;
17'h1628d:	data_out=16'h9f0;
17'h1628e:	data_out=16'h994;
17'h1628f:	data_out=16'h97f;
17'h16290:	data_out=16'h600;
17'h16291:	data_out=16'h81fe;
17'h16292:	data_out=16'h9b9;
17'h16293:	data_out=16'h8a00;
17'h16294:	data_out=16'h9e9;
17'h16295:	data_out=16'h8a00;
17'h16296:	data_out=16'h8a00;
17'h16297:	data_out=16'h9eb;
17'h16298:	data_out=16'h742;
17'h16299:	data_out=16'h8965;
17'h1629a:	data_out=16'h8536;
17'h1629b:	data_out=16'ha00;
17'h1629c:	data_out=16'ha00;
17'h1629d:	data_out=16'h89e4;
17'h1629e:	data_out=16'h99a;
17'h1629f:	data_out=16'h992;
17'h162a0:	data_out=16'h6a5;
17'h162a1:	data_out=16'ha00;
17'h162a2:	data_out=16'h8a00;
17'h162a3:	data_out=16'h89e6;
17'h162a4:	data_out=16'h89e6;
17'h162a5:	data_out=16'h8a00;
17'h162a6:	data_out=16'h90a;
17'h162a7:	data_out=16'h9ea;
17'h162a8:	data_out=16'ha00;
17'h162a9:	data_out=16'ha00;
17'h162aa:	data_out=16'h5a6;
17'h162ab:	data_out=16'h9f1;
17'h162ac:	data_out=16'h8a00;
17'h162ad:	data_out=16'h8a00;
17'h162ae:	data_out=16'h88c;
17'h162af:	data_out=16'h9f2;
17'h162b0:	data_out=16'h87a9;
17'h162b1:	data_out=16'h8640;
17'h162b2:	data_out=16'h8721;
17'h162b3:	data_out=16'h9f1;
17'h162b4:	data_out=16'h89f2;
17'h162b5:	data_out=16'h41f;
17'h162b6:	data_out=16'h9f6;
17'h162b7:	data_out=16'ha00;
17'h162b8:	data_out=16'h7f2;
17'h162b9:	data_out=16'h9f2;
17'h162ba:	data_out=16'h8a00;
17'h162bb:	data_out=16'h8376;
17'h162bc:	data_out=16'ha00;
17'h162bd:	data_out=16'h8a00;
17'h162be:	data_out=16'ha00;
17'h162bf:	data_out=16'h83bd;
17'h162c0:	data_out=16'h89e8;
17'h162c1:	data_out=16'ha00;
17'h162c2:	data_out=16'h89fa;
17'h162c3:	data_out=16'h9f5;
17'h162c4:	data_out=16'h8528;
17'h162c5:	data_out=16'h8a00;
17'h162c6:	data_out=16'ha00;
17'h162c7:	data_out=16'h8a00;
17'h162c8:	data_out=16'h204;
17'h162c9:	data_out=16'h89ff;
17'h162ca:	data_out=16'h9f1;
17'h162cb:	data_out=16'h828b;
17'h162cc:	data_out=16'h8a00;
17'h162cd:	data_out=16'h89fb;
17'h162ce:	data_out=16'ha00;
17'h162cf:	data_out=16'h8a00;
17'h162d0:	data_out=16'h8a00;
17'h162d1:	data_out=16'h9f1;
17'h162d2:	data_out=16'h8a00;
17'h162d3:	data_out=16'ha00;
17'h162d4:	data_out=16'h75d;
17'h162d5:	data_out=16'h9eb;
17'h162d6:	data_out=16'h867c;
17'h162d7:	data_out=16'h89fb;
17'h162d8:	data_out=16'ha00;
17'h162d9:	data_out=16'h89fc;
17'h162da:	data_out=16'ha00;
17'h162db:	data_out=16'h8165;
17'h162dc:	data_out=16'ha00;
17'h162dd:	data_out=16'h89fd;
17'h162de:	data_out=16'h9e1;
17'h162df:	data_out=16'h4b0;
17'h162e0:	data_out=16'h8a00;
17'h162e1:	data_out=16'h84d0;
17'h162e2:	data_out=16'h85a;
17'h162e3:	data_out=16'h9f5;
17'h162e4:	data_out=16'h8a00;
17'h162e5:	data_out=16'h89ff;
17'h162e6:	data_out=16'h897a;
17'h162e7:	data_out=16'h523;
17'h162e8:	data_out=16'ha00;
17'h162e9:	data_out=16'h9fe;
17'h162ea:	data_out=16'h854;
17'h162eb:	data_out=16'h89fb;
17'h162ec:	data_out=16'h89ee;
17'h162ed:	data_out=16'h9f3;
17'h162ee:	data_out=16'h855;
17'h162ef:	data_out=16'h8728;
17'h162f0:	data_out=16'h8fa;
17'h162f1:	data_out=16'h917;
17'h162f2:	data_out=16'h8a00;
17'h162f3:	data_out=16'h89e8;
17'h162f4:	data_out=16'h870f;
17'h162f5:	data_out=16'ha00;
17'h162f6:	data_out=16'h854;
17'h162f7:	data_out=16'h495;
17'h162f8:	data_out=16'ha00;
17'h162f9:	data_out=16'h9ff;
17'h162fa:	data_out=16'h9f3;
17'h162fb:	data_out=16'ha00;
17'h162fc:	data_out=16'h687;
17'h162fd:	data_out=16'h853;
17'h162fe:	data_out=16'h815e;
17'h162ff:	data_out=16'h89f6;
17'h16300:	data_out=16'h8a00;
17'h16301:	data_out=16'h885c;
17'h16302:	data_out=16'ha00;
17'h16303:	data_out=16'h741;
17'h16304:	data_out=16'h89db;
17'h16305:	data_out=16'h8362;
17'h16306:	data_out=16'h8a00;
17'h16307:	data_out=16'h89ff;
17'h16308:	data_out=16'ha00;
17'h16309:	data_out=16'h8a00;
17'h1630a:	data_out=16'h89cd;
17'h1630b:	data_out=16'h7f5;
17'h1630c:	data_out=16'h1dc;
17'h1630d:	data_out=16'h8cf;
17'h1630e:	data_out=16'ha00;
17'h1630f:	data_out=16'h9b0;
17'h16310:	data_out=16'h31a;
17'h16311:	data_out=16'h57a;
17'h16312:	data_out=16'h8f6;
17'h16313:	data_out=16'h8a00;
17'h16314:	data_out=16'h9c4;
17'h16315:	data_out=16'h8a00;
17'h16316:	data_out=16'h8a00;
17'h16317:	data_out=16'h9bf;
17'h16318:	data_out=16'h7fd;
17'h16319:	data_out=16'h87d9;
17'h1631a:	data_out=16'h83da;
17'h1631b:	data_out=16'ha00;
17'h1631c:	data_out=16'ha00;
17'h1631d:	data_out=16'h89dc;
17'h1631e:	data_out=16'h82a;
17'h1631f:	data_out=16'h869;
17'h16320:	data_out=16'h898e;
17'h16321:	data_out=16'ha00;
17'h16322:	data_out=16'h892a;
17'h16323:	data_out=16'h8439;
17'h16324:	data_out=16'h8410;
17'h16325:	data_out=16'h89fe;
17'h16326:	data_out=16'h99a;
17'h16327:	data_out=16'h15;
17'h16328:	data_out=16'ha00;
17'h16329:	data_out=16'ha00;
17'h1632a:	data_out=16'hf8;
17'h1632b:	data_out=16'h999;
17'h1632c:	data_out=16'h8a00;
17'h1632d:	data_out=16'h8285;
17'h1632e:	data_out=16'h827;
17'h1632f:	data_out=16'h9db;
17'h16330:	data_out=16'h8527;
17'h16331:	data_out=16'h8792;
17'h16332:	data_out=16'h83f6;
17'h16333:	data_out=16'h9e4;
17'h16334:	data_out=16'h89f9;
17'h16335:	data_out=16'h8006;
17'h16336:	data_out=16'h9f8;
17'h16337:	data_out=16'ha00;
17'h16338:	data_out=16'h970;
17'h16339:	data_out=16'h9dc;
17'h1633a:	data_out=16'h8a00;
17'h1633b:	data_out=16'h8216;
17'h1633c:	data_out=16'ha00;
17'h1633d:	data_out=16'h8a00;
17'h1633e:	data_out=16'ha00;
17'h1633f:	data_out=16'h8375;
17'h16340:	data_out=16'h893b;
17'h16341:	data_out=16'ha00;
17'h16342:	data_out=16'h89fa;
17'h16343:	data_out=16'h9f1;
17'h16344:	data_out=16'h85e1;
17'h16345:	data_out=16'h8a00;
17'h16346:	data_out=16'ha00;
17'h16347:	data_out=16'h8a00;
17'h16348:	data_out=16'h8531;
17'h16349:	data_out=16'h89f3;
17'h1634a:	data_out=16'h9ea;
17'h1634b:	data_out=16'h8a00;
17'h1634c:	data_out=16'h89f9;
17'h1634d:	data_out=16'h8959;
17'h1634e:	data_out=16'ha00;
17'h1634f:	data_out=16'h8a00;
17'h16350:	data_out=16'h8a00;
17'h16351:	data_out=16'h9e8;
17'h16352:	data_out=16'h89f6;
17'h16353:	data_out=16'ha00;
17'h16354:	data_out=16'h2db;
17'h16355:	data_out=16'h9eb;
17'h16356:	data_out=16'h2d2;
17'h16357:	data_out=16'h89e0;
17'h16358:	data_out=16'ha00;
17'h16359:	data_out=16'h89ec;
17'h1635a:	data_out=16'ha00;
17'h1635b:	data_out=16'h9e7;
17'h1635c:	data_out=16'ha00;
17'h1635d:	data_out=16'h89fb;
17'h1635e:	data_out=16'h7a1;
17'h1635f:	data_out=16'h1bd;
17'h16360:	data_out=16'h89fa;
17'h16361:	data_out=16'h8169;
17'h16362:	data_out=16'h3c5;
17'h16363:	data_out=16'h9e8;
17'h16364:	data_out=16'h8a00;
17'h16365:	data_out=16'h89fc;
17'h16366:	data_out=16'h89dd;
17'h16367:	data_out=16'h6ff;
17'h16368:	data_out=16'ha00;
17'h16369:	data_out=16'h9fb;
17'h1636a:	data_out=16'ha00;
17'h1636b:	data_out=16'h89fd;
17'h1636c:	data_out=16'h89fa;
17'h1636d:	data_out=16'h9e7;
17'h1636e:	data_out=16'ha00;
17'h1636f:	data_out=16'h882e;
17'h16370:	data_out=16'ha00;
17'h16371:	data_out=16'h6d5;
17'h16372:	data_out=16'h89fe;
17'h16373:	data_out=16'h89b8;
17'h16374:	data_out=16'h8458;
17'h16375:	data_out=16'ha00;
17'h16376:	data_out=16'h7b2;
17'h16377:	data_out=16'h28b;
17'h16378:	data_out=16'ha00;
17'h16379:	data_out=16'ha00;
17'h1637a:	data_out=16'h9ea;
17'h1637b:	data_out=16'ha00;
17'h1637c:	data_out=16'h4b5;
17'h1637d:	data_out=16'h6c0;
17'h1637e:	data_out=16'h1bc;
17'h1637f:	data_out=16'h89fa;
17'h16380:	data_out=16'h89f2;
17'h16381:	data_out=16'h8707;
17'h16382:	data_out=16'ha00;
17'h16383:	data_out=16'h759;
17'h16384:	data_out=16'h89c1;
17'h16385:	data_out=16'h8249;
17'h16386:	data_out=16'h8a00;
17'h16387:	data_out=16'h89ff;
17'h16388:	data_out=16'ha00;
17'h16389:	data_out=16'h8a00;
17'h1638a:	data_out=16'h89b0;
17'h1638b:	data_out=16'h781;
17'h1638c:	data_out=16'h481;
17'h1638d:	data_out=16'h815;
17'h1638e:	data_out=16'ha00;
17'h1638f:	data_out=16'h968;
17'h16390:	data_out=16'h2b5;
17'h16391:	data_out=16'ha00;
17'h16392:	data_out=16'h8fc;
17'h16393:	data_out=16'h8a00;
17'h16394:	data_out=16'h947;
17'h16395:	data_out=16'h89fc;
17'h16396:	data_out=16'h8a00;
17'h16397:	data_out=16'h95e;
17'h16398:	data_out=16'h5a7;
17'h16399:	data_out=16'h932;
17'h1639a:	data_out=16'h844a;
17'h1639b:	data_out=16'ha00;
17'h1639c:	data_out=16'ha00;
17'h1639d:	data_out=16'h8993;
17'h1639e:	data_out=16'h80d;
17'h1639f:	data_out=16'h816c;
17'h163a0:	data_out=16'h2ed;
17'h163a1:	data_out=16'ha00;
17'h163a2:	data_out=16'h824e;
17'h163a3:	data_out=16'h3cb;
17'h163a4:	data_out=16'h3e8;
17'h163a5:	data_out=16'h8a00;
17'h163a6:	data_out=16'h957;
17'h163a7:	data_out=16'ha00;
17'h163a8:	data_out=16'ha00;
17'h163a9:	data_out=16'ha00;
17'h163aa:	data_out=16'h42f;
17'h163ab:	data_out=16'h9a1;
17'h163ac:	data_out=16'h8a00;
17'h163ad:	data_out=16'h922;
17'h163ae:	data_out=16'h844;
17'h163af:	data_out=16'h9bf;
17'h163b0:	data_out=16'h832e;
17'h163b1:	data_out=16'h88c1;
17'h163b2:	data_out=16'h8337;
17'h163b3:	data_out=16'h9a6;
17'h163b4:	data_out=16'h89ef;
17'h163b5:	data_out=16'h4f6;
17'h163b6:	data_out=16'h9ff;
17'h163b7:	data_out=16'ha00;
17'h163b8:	data_out=16'h9b6;
17'h163b9:	data_out=16'h985;
17'h163ba:	data_out=16'h8a00;
17'h163bb:	data_out=16'h810e;
17'h163bc:	data_out=16'ha00;
17'h163bd:	data_out=16'h89f5;
17'h163be:	data_out=16'ha00;
17'h163bf:	data_out=16'h82ce;
17'h163c0:	data_out=16'h8907;
17'h163c1:	data_out=16'ha00;
17'h163c2:	data_out=16'h8a00;
17'h163c3:	data_out=16'h4f8;
17'h163c4:	data_out=16'h8631;
17'h163c5:	data_out=16'h89fd;
17'h163c6:	data_out=16'ha00;
17'h163c7:	data_out=16'h8a00;
17'h163c8:	data_out=16'h8464;
17'h163c9:	data_out=16'h89fd;
17'h163ca:	data_out=16'h9f2;
17'h163cb:	data_out=16'h8a00;
17'h163cc:	data_out=16'h89ef;
17'h163cd:	data_out=16'h80c7;
17'h163ce:	data_out=16'ha00;
17'h163cf:	data_out=16'h8a00;
17'h163d0:	data_out=16'h8a00;
17'h163d1:	data_out=16'h9ec;
17'h163d2:	data_out=16'h89e9;
17'h163d3:	data_out=16'ha00;
17'h163d4:	data_out=16'h8f8;
17'h163d5:	data_out=16'h9c1;
17'h163d6:	data_out=16'h9fe;
17'h163d7:	data_out=16'h89d2;
17'h163d8:	data_out=16'ha00;
17'h163d9:	data_out=16'h89cf;
17'h163da:	data_out=16'ha00;
17'h163db:	data_out=16'ha00;
17'h163dc:	data_out=16'ha00;
17'h163dd:	data_out=16'h8279;
17'h163de:	data_out=16'h954;
17'h163df:	data_out=16'h362;
17'h163e0:	data_out=16'h89fb;
17'h163e1:	data_out=16'h6eb;
17'h163e2:	data_out=16'h449;
17'h163e3:	data_out=16'h9c9;
17'h163e4:	data_out=16'h8a00;
17'h163e5:	data_out=16'h89fb;
17'h163e6:	data_out=16'h83d8;
17'h163e7:	data_out=16'h9ed;
17'h163e8:	data_out=16'ha00;
17'h163e9:	data_out=16'h9e9;
17'h163ea:	data_out=16'ha00;
17'h163eb:	data_out=16'h89f8;
17'h163ec:	data_out=16'h89e9;
17'h163ed:	data_out=16'h9c2;
17'h163ee:	data_out=16'ha00;
17'h163ef:	data_out=16'h8909;
17'h163f0:	data_out=16'ha00;
17'h163f1:	data_out=16'h532;
17'h163f2:	data_out=16'h89e7;
17'h163f3:	data_out=16'h8997;
17'h163f4:	data_out=16'h813c;
17'h163f5:	data_out=16'ha00;
17'h163f6:	data_out=16'h962;
17'h163f7:	data_out=16'h480;
17'h163f8:	data_out=16'ha00;
17'h163f9:	data_out=16'ha00;
17'h163fa:	data_out=16'h9c1;
17'h163fb:	data_out=16'ha00;
17'h163fc:	data_out=16'h138;
17'h163fd:	data_out=16'h89f5;
17'h163fe:	data_out=16'h8934;
17'h163ff:	data_out=16'h89f5;
17'h16400:	data_out=16'h8a00;
17'h16401:	data_out=16'h873e;
17'h16402:	data_out=16'ha00;
17'h16403:	data_out=16'h758;
17'h16404:	data_out=16'h8645;
17'h16405:	data_out=16'h9af;
17'h16406:	data_out=16'h8a00;
17'h16407:	data_out=16'h8a00;
17'h16408:	data_out=16'ha00;
17'h16409:	data_out=16'h8a00;
17'h1640a:	data_out=16'h8a00;
17'h1640b:	data_out=16'h867;
17'h1640c:	data_out=16'h584;
17'h1640d:	data_out=16'h543;
17'h1640e:	data_out=16'ha00;
17'h1640f:	data_out=16'h8fd;
17'h16410:	data_out=16'h329;
17'h16411:	data_out=16'h9e9;
17'h16412:	data_out=16'h984;
17'h16413:	data_out=16'h8a00;
17'h16414:	data_out=16'h8fc;
17'h16415:	data_out=16'h8a00;
17'h16416:	data_out=16'h8a00;
17'h16417:	data_out=16'h916;
17'h16418:	data_out=16'h573;
17'h16419:	data_out=16'h9f8;
17'h1641a:	data_out=16'h4d2;
17'h1641b:	data_out=16'ha00;
17'h1641c:	data_out=16'ha00;
17'h1641d:	data_out=16'h89ff;
17'h1641e:	data_out=16'h80b;
17'h1641f:	data_out=16'h88de;
17'h16420:	data_out=16'h8a7;
17'h16421:	data_out=16'ha00;
17'h16422:	data_out=16'h496;
17'h16423:	data_out=16'h8391;
17'h16424:	data_out=16'h8366;
17'h16425:	data_out=16'h8a00;
17'h16426:	data_out=16'h7b1;
17'h16427:	data_out=16'h9b5;
17'h16428:	data_out=16'ha00;
17'h16429:	data_out=16'ha00;
17'h1642a:	data_out=16'h34a;
17'h1642b:	data_out=16'h991;
17'h1642c:	data_out=16'h8a00;
17'h1642d:	data_out=16'h9ac;
17'h1642e:	data_out=16'h7d7;
17'h1642f:	data_out=16'h953;
17'h16430:	data_out=16'h9fd;
17'h16431:	data_out=16'h89ff;
17'h16432:	data_out=16'haa;
17'h16433:	data_out=16'h9a7;
17'h16434:	data_out=16'h8a00;
17'h16435:	data_out=16'h654;
17'h16436:	data_out=16'h9e4;
17'h16437:	data_out=16'ha00;
17'h16438:	data_out=16'h9bc;
17'h16439:	data_out=16'h9b3;
17'h1643a:	data_out=16'h8a00;
17'h1643b:	data_out=16'h8416;
17'h1643c:	data_out=16'ha00;
17'h1643d:	data_out=16'h8a00;
17'h1643e:	data_out=16'ha00;
17'h1643f:	data_out=16'h940;
17'h16440:	data_out=16'h89ea;
17'h16441:	data_out=16'ha00;
17'h16442:	data_out=16'h8a00;
17'h16443:	data_out=16'h80b7;
17'h16444:	data_out=16'h850a;
17'h16445:	data_out=16'h8a00;
17'h16446:	data_out=16'ha00;
17'h16447:	data_out=16'h8a00;
17'h16448:	data_out=16'h86a5;
17'h16449:	data_out=16'h89fb;
17'h1644a:	data_out=16'h9bb;
17'h1644b:	data_out=16'h8a00;
17'h1644c:	data_out=16'h89f2;
17'h1644d:	data_out=16'h806;
17'h1644e:	data_out=16'h919;
17'h1644f:	data_out=16'h8a00;
17'h16450:	data_out=16'h89da;
17'h16451:	data_out=16'h9ed;
17'h16452:	data_out=16'h8a00;
17'h16453:	data_out=16'h9d8;
17'h16454:	data_out=16'h8e5;
17'h16455:	data_out=16'h918;
17'h16456:	data_out=16'h9fe;
17'h16457:	data_out=16'h89ea;
17'h16458:	data_out=16'ha00;
17'h16459:	data_out=16'h8a00;
17'h1645a:	data_out=16'ha00;
17'h1645b:	data_out=16'h9cf;
17'h1645c:	data_out=16'ha00;
17'h1645d:	data_out=16'h721;
17'h1645e:	data_out=16'h8e0;
17'h1645f:	data_out=16'h264;
17'h16460:	data_out=16'h89f5;
17'h16461:	data_out=16'h9f6;
17'h16462:	data_out=16'h636;
17'h16463:	data_out=16'h9b8;
17'h16464:	data_out=16'h8a00;
17'h16465:	data_out=16'h8a00;
17'h16466:	data_out=16'h3da;
17'h16467:	data_out=16'h9de;
17'h16468:	data_out=16'ha00;
17'h16469:	data_out=16'ha00;
17'h1646a:	data_out=16'ha00;
17'h1646b:	data_out=16'h8a00;
17'h1646c:	data_out=16'h8a00;
17'h1646d:	data_out=16'h9ab;
17'h1646e:	data_out=16'ha00;
17'h1646f:	data_out=16'h8a00;
17'h16470:	data_out=16'ha00;
17'h16471:	data_out=16'h83e5;
17'h16472:	data_out=16'h8a00;
17'h16473:	data_out=16'h8a00;
17'h16474:	data_out=16'ha00;
17'h16475:	data_out=16'ha00;
17'h16476:	data_out=16'h9b8;
17'h16477:	data_out=16'h439;
17'h16478:	data_out=16'ha00;
17'h16479:	data_out=16'ha00;
17'h1647a:	data_out=16'h978;
17'h1647b:	data_out=16'ha00;
17'h1647c:	data_out=16'h80f2;
17'h1647d:	data_out=16'h89ff;
17'h1647e:	data_out=16'h8964;
17'h1647f:	data_out=16'h8a00;
17'h16480:	data_out=16'h89fe;
17'h16481:	data_out=16'h80c0;
17'h16482:	data_out=16'ha00;
17'h16483:	data_out=16'h430;
17'h16484:	data_out=16'h89bf;
17'h16485:	data_out=16'h1bd;
17'h16486:	data_out=16'h8a00;
17'h16487:	data_out=16'h8a00;
17'h16488:	data_out=16'ha00;
17'h16489:	data_out=16'h8a00;
17'h1648a:	data_out=16'h8a00;
17'h1648b:	data_out=16'h8a3;
17'h1648c:	data_out=16'h80b8;
17'h1648d:	data_out=16'h84e3;
17'h1648e:	data_out=16'ha00;
17'h1648f:	data_out=16'h872;
17'h16490:	data_out=16'h8278;
17'h16491:	data_out=16'h6f2;
17'h16492:	data_out=16'h9ac;
17'h16493:	data_out=16'h8a00;
17'h16494:	data_out=16'h7c3;
17'h16495:	data_out=16'h8a00;
17'h16496:	data_out=16'h8a00;
17'h16497:	data_out=16'h7ba;
17'h16498:	data_out=16'h9a9;
17'h16499:	data_out=16'h9c2;
17'h1649a:	data_out=16'h8242;
17'h1649b:	data_out=16'ha00;
17'h1649c:	data_out=16'h9fb;
17'h1649d:	data_out=16'h8978;
17'h1649e:	data_out=16'h687;
17'h1649f:	data_out=16'h8848;
17'h164a0:	data_out=16'h1b2;
17'h164a1:	data_out=16'ha00;
17'h164a2:	data_out=16'h87b;
17'h164a3:	data_out=16'h899a;
17'h164a4:	data_out=16'h8988;
17'h164a5:	data_out=16'h8a00;
17'h164a6:	data_out=16'h6da;
17'h164a7:	data_out=16'h788;
17'h164a8:	data_out=16'ha00;
17'h164a9:	data_out=16'ha00;
17'h164aa:	data_out=16'h24a;
17'h164ab:	data_out=16'h41e;
17'h164ac:	data_out=16'h8a00;
17'h164ad:	data_out=16'h993;
17'h164ae:	data_out=16'h717;
17'h164af:	data_out=16'h834;
17'h164b0:	data_out=16'h9dd;
17'h164b1:	data_out=16'h8a00;
17'h164b2:	data_out=16'h82d2;
17'h164b3:	data_out=16'h976;
17'h164b4:	data_out=16'h8a00;
17'h164b5:	data_out=16'haa;
17'h164b6:	data_out=16'h9cb;
17'h164b7:	data_out=16'ha00;
17'h164b8:	data_out=16'h9b1;
17'h164b9:	data_out=16'h9a6;
17'h164ba:	data_out=16'h8a00;
17'h164bb:	data_out=16'h89ff;
17'h164bc:	data_out=16'ha00;
17'h164bd:	data_out=16'h8a00;
17'h164be:	data_out=16'ha00;
17'h164bf:	data_out=16'h175;
17'h164c0:	data_out=16'h8a00;
17'h164c1:	data_out=16'h9ff;
17'h164c2:	data_out=16'h8a00;
17'h164c3:	data_out=16'h8490;
17'h164c4:	data_out=16'h8a00;
17'h164c5:	data_out=16'h8a00;
17'h164c6:	data_out=16'ha00;
17'h164c7:	data_out=16'h8a00;
17'h164c8:	data_out=16'h8263;
17'h164c9:	data_out=16'h89ef;
17'h164ca:	data_out=16'h210;
17'h164cb:	data_out=16'h8a00;
17'h164cc:	data_out=16'h89da;
17'h164cd:	data_out=16'h8b3;
17'h164ce:	data_out=16'ha00;
17'h164cf:	data_out=16'h8a00;
17'h164d0:	data_out=16'h8a00;
17'h164d1:	data_out=16'h9d6;
17'h164d2:	data_out=16'h8a00;
17'h164d3:	data_out=16'h97d;
17'h164d4:	data_out=16'h7ca;
17'h164d5:	data_out=16'h7fa;
17'h164d6:	data_out=16'h9fa;
17'h164d7:	data_out=16'h423;
17'h164d8:	data_out=16'ha00;
17'h164d9:	data_out=16'h8a00;
17'h164da:	data_out=16'ha00;
17'h164db:	data_out=16'h51f;
17'h164dc:	data_out=16'h9f6;
17'h164dd:	data_out=16'h696;
17'h164de:	data_out=16'h6f8;
17'h164df:	data_out=16'h906;
17'h164e0:	data_out=16'h89f0;
17'h164e1:	data_out=16'h934;
17'h164e2:	data_out=16'h43a;
17'h164e3:	data_out=16'h963;
17'h164e4:	data_out=16'h8a00;
17'h164e5:	data_out=16'h8a00;
17'h164e6:	data_out=16'he9;
17'h164e7:	data_out=16'h9e2;
17'h164e8:	data_out=16'ha00;
17'h164e9:	data_out=16'ha00;
17'h164ea:	data_out=16'ha00;
17'h164eb:	data_out=16'h8a00;
17'h164ec:	data_out=16'h8a00;
17'h164ed:	data_out=16'h95d;
17'h164ee:	data_out=16'ha00;
17'h164ef:	data_out=16'h8a00;
17'h164f0:	data_out=16'ha00;
17'h164f1:	data_out=16'h144;
17'h164f2:	data_out=16'h8a00;
17'h164f3:	data_out=16'h88fb;
17'h164f4:	data_out=16'h9f8;
17'h164f5:	data_out=16'h9e4;
17'h164f6:	data_out=16'h9d4;
17'h164f7:	data_out=16'h14e;
17'h164f8:	data_out=16'h6b1;
17'h164f9:	data_out=16'ha00;
17'h164fa:	data_out=16'h8c9;
17'h164fb:	data_out=16'ha00;
17'h164fc:	data_out=16'h3ea;
17'h164fd:	data_out=16'h8a00;
17'h164fe:	data_out=16'h89f7;
17'h164ff:	data_out=16'h8618;
17'h16500:	data_out=16'h89f3;
17'h16501:	data_out=16'h889;
17'h16502:	data_out=16'ha00;
17'h16503:	data_out=16'h1af;
17'h16504:	data_out=16'h8a00;
17'h16505:	data_out=16'h8032;
17'h16506:	data_out=16'h8a00;
17'h16507:	data_out=16'h8a00;
17'h16508:	data_out=16'h9fc;
17'h16509:	data_out=16'h8a00;
17'h1650a:	data_out=16'h8a00;
17'h1650b:	data_out=16'h838;
17'h1650c:	data_out=16'h8a00;
17'h1650d:	data_out=16'h89f2;
17'h1650e:	data_out=16'ha00;
17'h1650f:	data_out=16'h8c3;
17'h16510:	data_out=16'h87de;
17'h16511:	data_out=16'h8204;
17'h16512:	data_out=16'h9d9;
17'h16513:	data_out=16'h8a00;
17'h16514:	data_out=16'h723;
17'h16515:	data_out=16'h8a00;
17'h16516:	data_out=16'h8a00;
17'h16517:	data_out=16'h747;
17'h16518:	data_out=16'h28e;
17'h16519:	data_out=16'h9d0;
17'h1651a:	data_out=16'h842d;
17'h1651b:	data_out=16'h9f3;
17'h1651c:	data_out=16'h9f0;
17'h1651d:	data_out=16'h23d;
17'h1651e:	data_out=16'h6f9;
17'h1651f:	data_out=16'h8a00;
17'h16520:	data_out=16'h588;
17'h16521:	data_out=16'ha00;
17'h16522:	data_out=16'h9da;
17'h16523:	data_out=16'h89e6;
17'h16524:	data_out=16'h89e6;
17'h16525:	data_out=16'h89fe;
17'h16526:	data_out=16'h8472;
17'h16527:	data_out=16'h696;
17'h16528:	data_out=16'ha00;
17'h16529:	data_out=16'ha00;
17'h1652a:	data_out=16'h491;
17'h1652b:	data_out=16'h8689;
17'h1652c:	data_out=16'h8a00;
17'h1652d:	data_out=16'h9e6;
17'h1652e:	data_out=16'h831;
17'h1652f:	data_out=16'h8e7;
17'h16530:	data_out=16'h9ea;
17'h16531:	data_out=16'h8a00;
17'h16532:	data_out=16'h162;
17'h16533:	data_out=16'h96a;
17'h16534:	data_out=16'h89fd;
17'h16535:	data_out=16'h80ab;
17'h16536:	data_out=16'h9db;
17'h16537:	data_out=16'ha00;
17'h16538:	data_out=16'h9ea;
17'h16539:	data_out=16'h99f;
17'h1653a:	data_out=16'h8a00;
17'h1653b:	data_out=16'h8a00;
17'h1653c:	data_out=16'h9f8;
17'h1653d:	data_out=16'h8a00;
17'h1653e:	data_out=16'ha00;
17'h1653f:	data_out=16'h806d;
17'h16540:	data_out=16'h8a00;
17'h16541:	data_out=16'h9f1;
17'h16542:	data_out=16'h8a00;
17'h16543:	data_out=16'h83a7;
17'h16544:	data_out=16'h8a00;
17'h16545:	data_out=16'h8a00;
17'h16546:	data_out=16'ha00;
17'h16547:	data_out=16'h89ff;
17'h16548:	data_out=16'h316;
17'h16549:	data_out=16'h89ef;
17'h1654a:	data_out=16'h830c;
17'h1654b:	data_out=16'h8a00;
17'h1654c:	data_out=16'h8669;
17'h1654d:	data_out=16'h9d7;
17'h1654e:	data_out=16'ha00;
17'h1654f:	data_out=16'h89fa;
17'h16550:	data_out=16'h8a00;
17'h16551:	data_out=16'h22a;
17'h16552:	data_out=16'h89f3;
17'h16553:	data_out=16'h9ad;
17'h16554:	data_out=16'h8b2;
17'h16555:	data_out=16'h714;
17'h16556:	data_out=16'h8cd;
17'h16557:	data_out=16'h46b;
17'h16558:	data_out=16'ha00;
17'h16559:	data_out=16'h8a00;
17'h1655a:	data_out=16'ha00;
17'h1655b:	data_out=16'h38f;
17'h1655c:	data_out=16'h9ef;
17'h1655d:	data_out=16'h805;
17'h1655e:	data_out=16'h7ce;
17'h1655f:	data_out=16'h982;
17'h16560:	data_out=16'h863d;
17'h16561:	data_out=16'h684;
17'h16562:	data_out=16'h508;
17'h16563:	data_out=16'h970;
17'h16564:	data_out=16'h89fe;
17'h16565:	data_out=16'h8a00;
17'h16566:	data_out=16'h842f;
17'h16567:	data_out=16'ha00;
17'h16568:	data_out=16'ha00;
17'h16569:	data_out=16'h9fd;
17'h1656a:	data_out=16'ha00;
17'h1656b:	data_out=16'h8a00;
17'h1656c:	data_out=16'h8704;
17'h1656d:	data_out=16'h96b;
17'h1656e:	data_out=16'ha00;
17'h1656f:	data_out=16'h8a00;
17'h16570:	data_out=16'ha00;
17'h16571:	data_out=16'h6f7;
17'h16572:	data_out=16'h88c2;
17'h16573:	data_out=16'h242;
17'h16574:	data_out=16'h9fe;
17'h16575:	data_out=16'h9d1;
17'h16576:	data_out=16'h9e2;
17'h16577:	data_out=16'h87a5;
17'h16578:	data_out=16'h8a7;
17'h16579:	data_out=16'ha00;
17'h1657a:	data_out=16'h8a2;
17'h1657b:	data_out=16'ha00;
17'h1657c:	data_out=16'h255;
17'h1657d:	data_out=16'h8a00;
17'h1657e:	data_out=16'h89ee;
17'h1657f:	data_out=16'h23c;
17'h16580:	data_out=16'h879b;
17'h16581:	data_out=16'h942;
17'h16582:	data_out=16'h9fc;
17'h16583:	data_out=16'h506;
17'h16584:	data_out=16'h8a00;
17'h16585:	data_out=16'h888b;
17'h16586:	data_out=16'h8a00;
17'h16587:	data_out=16'h8a00;
17'h16588:	data_out=16'h9f9;
17'h16589:	data_out=16'h8a00;
17'h1658a:	data_out=16'h8a00;
17'h1658b:	data_out=16'h943;
17'h1658c:	data_out=16'h8a00;
17'h1658d:	data_out=16'h8a00;
17'h1658e:	data_out=16'ha00;
17'h1658f:	data_out=16'h923;
17'h16590:	data_out=16'h70e;
17'h16591:	data_out=16'h8520;
17'h16592:	data_out=16'h9f5;
17'h16593:	data_out=16'h8a00;
17'h16594:	data_out=16'h6b3;
17'h16595:	data_out=16'h8a00;
17'h16596:	data_out=16'h8a00;
17'h16597:	data_out=16'h6d6;
17'h16598:	data_out=16'h4ed;
17'h16599:	data_out=16'h9df;
17'h1659a:	data_out=16'h8753;
17'h1659b:	data_out=16'h9dd;
17'h1659c:	data_out=16'h9d4;
17'h1659d:	data_out=16'h7db;
17'h1659e:	data_out=16'h7cd;
17'h1659f:	data_out=16'h8a00;
17'h165a0:	data_out=16'h6cb;
17'h165a1:	data_out=16'ha00;
17'h165a2:	data_out=16'ha00;
17'h165a3:	data_out=16'h89e5;
17'h165a4:	data_out=16'h89e5;
17'h165a5:	data_out=16'h89fd;
17'h165a6:	data_out=16'h8a5;
17'h165a7:	data_out=16'h70e;
17'h165a8:	data_out=16'ha00;
17'h165a9:	data_out=16'ha00;
17'h165aa:	data_out=16'h706;
17'h165ab:	data_out=16'h85a;
17'h165ac:	data_out=16'h8a00;
17'h165ad:	data_out=16'h9fb;
17'h165ae:	data_out=16'h8ed;
17'h165af:	data_out=16'h8ff;
17'h165b0:	data_out=16'h931;
17'h165b1:	data_out=16'h8a00;
17'h165b2:	data_out=16'h801f;
17'h165b3:	data_out=16'h96d;
17'h165b4:	data_out=16'h8378;
17'h165b5:	data_out=16'h85bb;
17'h165b6:	data_out=16'h9e4;
17'h165b7:	data_out=16'h9fe;
17'h165b8:	data_out=16'h9fa;
17'h165b9:	data_out=16'h9a8;
17'h165ba:	data_out=16'h8a00;
17'h165bb:	data_out=16'h8a00;
17'h165bc:	data_out=16'ha00;
17'h165bd:	data_out=16'h82a2;
17'h165be:	data_out=16'ha00;
17'h165bf:	data_out=16'h88be;
17'h165c0:	data_out=16'h8a00;
17'h165c1:	data_out=16'h9ea;
17'h165c2:	data_out=16'hcc;
17'h165c3:	data_out=16'h887f;
17'h165c4:	data_out=16'h8a00;
17'h165c5:	data_out=16'h8a00;
17'h165c6:	data_out=16'ha00;
17'h165c7:	data_out=16'h8a00;
17'h165c8:	data_out=16'h692;
17'h165c9:	data_out=16'h89f5;
17'h165ca:	data_out=16'h843b;
17'h165cb:	data_out=16'h8606;
17'h165cc:	data_out=16'h816a;
17'h165cd:	data_out=16'ha00;
17'h165ce:	data_out=16'ha00;
17'h165cf:	data_out=16'h89fe;
17'h165d0:	data_out=16'h8365;
17'h165d1:	data_out=16'h87ef;
17'h165d2:	data_out=16'h89ed;
17'h165d3:	data_out=16'h9b2;
17'h165d4:	data_out=16'h905;
17'h165d5:	data_out=16'h6b8;
17'h165d6:	data_out=16'h9a4;
17'h165d7:	data_out=16'h63d;
17'h165d8:	data_out=16'ha00;
17'h165d9:	data_out=16'h8560;
17'h165da:	data_out=16'ha00;
17'h165db:	data_out=16'h51d;
17'h165dc:	data_out=16'h9f9;
17'h165dd:	data_out=16'h953;
17'h165de:	data_out=16'h886;
17'h165df:	data_out=16'h9bc;
17'h165e0:	data_out=16'h74b;
17'h165e1:	data_out=16'h803d;
17'h165e2:	data_out=16'h624;
17'h165e3:	data_out=16'h97b;
17'h165e4:	data_out=16'h89ff;
17'h165e5:	data_out=16'h8a00;
17'h165e6:	data_out=16'h94;
17'h165e7:	data_out=16'h9fc;
17'h165e8:	data_out=16'ha00;
17'h165e9:	data_out=16'h9f0;
17'h165ea:	data_out=16'ha00;
17'h165eb:	data_out=16'h8a00;
17'h165ec:	data_out=16'h7a9;
17'h165ed:	data_out=16'h977;
17'h165ee:	data_out=16'ha00;
17'h165ef:	data_out=16'h8a00;
17'h165f0:	data_out=16'ha00;
17'h165f1:	data_out=16'h71e;
17'h165f2:	data_out=16'h84e4;
17'h165f3:	data_out=16'h581;
17'h165f4:	data_out=16'h9a9;
17'h165f5:	data_out=16'h9c8;
17'h165f6:	data_out=16'h9f4;
17'h165f7:	data_out=16'h81d0;
17'h165f8:	data_out=16'h16f;
17'h165f9:	data_out=16'ha00;
17'h165fa:	data_out=16'h899;
17'h165fb:	data_out=16'ha00;
17'h165fc:	data_out=16'h447;
17'h165fd:	data_out=16'h8a00;
17'h165fe:	data_out=16'h8927;
17'h165ff:	data_out=16'h58c;
17'h16600:	data_out=16'h8657;
17'h16601:	data_out=16'h9f4;
17'h16602:	data_out=16'ha00;
17'h16603:	data_out=16'h6a8;
17'h16604:	data_out=16'h7f5;
17'h16605:	data_out=16'h9a1;
17'h16606:	data_out=16'h880d;
17'h16607:	data_out=16'h8a00;
17'h16608:	data_out=16'ha00;
17'h16609:	data_out=16'h8a00;
17'h1660a:	data_out=16'h1a7;
17'h1660b:	data_out=16'h9a1;
17'h1660c:	data_out=16'h84ea;
17'h1660d:	data_out=16'h8a00;
17'h1660e:	data_out=16'ha00;
17'h1660f:	data_out=16'h9ca;
17'h16610:	data_out=16'h7a1;
17'h16611:	data_out=16'h9bb;
17'h16612:	data_out=16'h9ff;
17'h16613:	data_out=16'h8058;
17'h16614:	data_out=16'h7f6;
17'h16615:	data_out=16'h8a00;
17'h16616:	data_out=16'h8a00;
17'h16617:	data_out=16'h85e;
17'h16618:	data_out=16'h1cf;
17'h16619:	data_out=16'h9f4;
17'h1661a:	data_out=16'h9bb;
17'h1661b:	data_out=16'h9e3;
17'h1661c:	data_out=16'h9c2;
17'h1661d:	data_out=16'h9bd;
17'h1661e:	data_out=16'h986;
17'h1661f:	data_out=16'h88af;
17'h16620:	data_out=16'h9b6;
17'h16621:	data_out=16'ha00;
17'h16622:	data_out=16'ha00;
17'h16623:	data_out=16'h89f0;
17'h16624:	data_out=16'h89ef;
17'h16625:	data_out=16'h89f6;
17'h16626:	data_out=16'h8f6;
17'h16627:	data_out=16'h9dc;
17'h16628:	data_out=16'ha00;
17'h16629:	data_out=16'ha00;
17'h1662a:	data_out=16'h99c;
17'h1662b:	data_out=16'h9be;
17'h1662c:	data_out=16'h8a00;
17'h1662d:	data_out=16'ha00;
17'h1662e:	data_out=16'h9c4;
17'h1662f:	data_out=16'h9b8;
17'h16630:	data_out=16'h9fc;
17'h16631:	data_out=16'h8a00;
17'h16632:	data_out=16'h9eb;
17'h16633:	data_out=16'h9d0;
17'h16634:	data_out=16'h7df;
17'h16635:	data_out=16'h8d5;
17'h16636:	data_out=16'ha00;
17'h16637:	data_out=16'ha00;
17'h16638:	data_out=16'h9fe;
17'h16639:	data_out=16'h9df;
17'h1663a:	data_out=16'h8a00;
17'h1663b:	data_out=16'h88f4;
17'h1663c:	data_out=16'ha00;
17'h1663d:	data_out=16'h967;
17'h1663e:	data_out=16'ha00;
17'h1663f:	data_out=16'h9a3;
17'h16640:	data_out=16'h969;
17'h16641:	data_out=16'ha00;
17'h16642:	data_out=16'h763;
17'h16643:	data_out=16'h8a00;
17'h16644:	data_out=16'h80c4;
17'h16645:	data_out=16'h8a00;
17'h16646:	data_out=16'ha00;
17'h16647:	data_out=16'h8a00;
17'h16648:	data_out=16'h98a;
17'h16649:	data_out=16'h8946;
17'h1664a:	data_out=16'h3a7;
17'h1664b:	data_out=16'h1df;
17'h1664c:	data_out=16'h83e5;
17'h1664d:	data_out=16'ha00;
17'h1664e:	data_out=16'ha00;
17'h1664f:	data_out=16'h8a00;
17'h16650:	data_out=16'h604;
17'h16651:	data_out=16'h87c;
17'h16652:	data_out=16'h89f2;
17'h16653:	data_out=16'h9ff;
17'h16654:	data_out=16'h9e8;
17'h16655:	data_out=16'h852;
17'h16656:	data_out=16'h9f4;
17'h16657:	data_out=16'h88a;
17'h16658:	data_out=16'ha00;
17'h16659:	data_out=16'h8f3;
17'h1665a:	data_out=16'ha00;
17'h1665b:	data_out=16'h9e9;
17'h1665c:	data_out=16'ha00;
17'h1665d:	data_out=16'ha00;
17'h1665e:	data_out=16'h9c2;
17'h1665f:	data_out=16'h9f9;
17'h16660:	data_out=16'h886;
17'h16661:	data_out=16'h9f5;
17'h16662:	data_out=16'h7cd;
17'h16663:	data_out=16'h9e0;
17'h16664:	data_out=16'h14;
17'h16665:	data_out=16'h8a00;
17'h16666:	data_out=16'h9e0;
17'h16667:	data_out=16'h9f7;
17'h16668:	data_out=16'ha00;
17'h16669:	data_out=16'h9f9;
17'h1666a:	data_out=16'ha00;
17'h1666b:	data_out=16'h652;
17'h1666c:	data_out=16'h764;
17'h1666d:	data_out=16'h9de;
17'h1666e:	data_out=16'ha00;
17'h1666f:	data_out=16'h748;
17'h16670:	data_out=16'ha00;
17'h16671:	data_out=16'h8275;
17'h16672:	data_out=16'h767;
17'h16673:	data_out=16'h982;
17'h16674:	data_out=16'ha00;
17'h16675:	data_out=16'ha00;
17'h16676:	data_out=16'h9fb;
17'h16677:	data_out=16'h550;
17'h16678:	data_out=16'h8164;
17'h16679:	data_out=16'ha00;
17'h1667a:	data_out=16'h990;
17'h1667b:	data_out=16'ha00;
17'h1667c:	data_out=16'h81ef;
17'h1667d:	data_out=16'h89e8;
17'h1667e:	data_out=16'h8274;
17'h1667f:	data_out=16'h981;
17'h16680:	data_out=16'ha00;
17'h16681:	data_out=16'h9f3;
17'h16682:	data_out=16'ha00;
17'h16683:	data_out=16'h928;
17'h16684:	data_out=16'h92d;
17'h16685:	data_out=16'h9e2;
17'h16686:	data_out=16'h8113;
17'h16687:	data_out=16'h8a00;
17'h16688:	data_out=16'ha00;
17'h16689:	data_out=16'h8a00;
17'h1668a:	data_out=16'h84a;
17'h1668b:	data_out=16'ha00;
17'h1668c:	data_out=16'h821b;
17'h1668d:	data_out=16'h8756;
17'h1668e:	data_out=16'ha00;
17'h1668f:	data_out=16'h9f7;
17'h16690:	data_out=16'h95d;
17'h16691:	data_out=16'h9af;
17'h16692:	data_out=16'ha00;
17'h16693:	data_out=16'h747;
17'h16694:	data_out=16'h984;
17'h16695:	data_out=16'h8618;
17'h16696:	data_out=16'h8583;
17'h16697:	data_out=16'h99f;
17'h16698:	data_out=16'h8487;
17'h16699:	data_out=16'h9f4;
17'h1669a:	data_out=16'h9e1;
17'h1669b:	data_out=16'ha00;
17'h1669c:	data_out=16'ha00;
17'h1669d:	data_out=16'h9e5;
17'h1669e:	data_out=16'h9ff;
17'h1669f:	data_out=16'h80eb;
17'h166a0:	data_out=16'h9f7;
17'h166a1:	data_out=16'ha00;
17'h166a2:	data_out=16'ha00;
17'h166a3:	data_out=16'h89f6;
17'h166a4:	data_out=16'h89f6;
17'h166a5:	data_out=16'h88b2;
17'h166a6:	data_out=16'h9a3;
17'h166a7:	data_out=16'h9f3;
17'h166a8:	data_out=16'ha00;
17'h166a9:	data_out=16'ha00;
17'h166aa:	data_out=16'h9eb;
17'h166ab:	data_out=16'h9f7;
17'h166ac:	data_out=16'h87f2;
17'h166ad:	data_out=16'ha00;
17'h166ae:	data_out=16'h9eb;
17'h166af:	data_out=16'h9f8;
17'h166b0:	data_out=16'h9fd;
17'h166b1:	data_out=16'h8337;
17'h166b2:	data_out=16'h9e5;
17'h166b3:	data_out=16'h9ff;
17'h166b4:	data_out=16'h9e6;
17'h166b5:	data_out=16'h9bd;
17'h166b6:	data_out=16'ha00;
17'h166b7:	data_out=16'ha00;
17'h166b8:	data_out=16'h9f5;
17'h166b9:	data_out=16'ha00;
17'h166ba:	data_out=16'h8a00;
17'h166bb:	data_out=16'h22d;
17'h166bc:	data_out=16'ha00;
17'h166bd:	data_out=16'h9f5;
17'h166be:	data_out=16'ha00;
17'h166bf:	data_out=16'h9e2;
17'h166c0:	data_out=16'h9b4;
17'h166c1:	data_out=16'ha00;
17'h166c2:	data_out=16'h948;
17'h166c3:	data_out=16'h8a00;
17'h166c4:	data_out=16'h9d9;
17'h166c5:	data_out=16'h861b;
17'h166c6:	data_out=16'ha00;
17'h166c7:	data_out=16'h89f2;
17'h166c8:	data_out=16'h9ed;
17'h166c9:	data_out=16'h8708;
17'h166ca:	data_out=16'h83fe;
17'h166cb:	data_out=16'h5ef;
17'h166cc:	data_out=16'h862c;
17'h166cd:	data_out=16'ha00;
17'h166ce:	data_out=16'ha00;
17'h166cf:	data_out=16'h8a00;
17'h166d0:	data_out=16'h8e4;
17'h166d1:	data_out=16'h99f;
17'h166d2:	data_out=16'h89f0;
17'h166d3:	data_out=16'h9fb;
17'h166d4:	data_out=16'h9fe;
17'h166d5:	data_out=16'h949;
17'h166d6:	data_out=16'ha00;
17'h166d7:	data_out=16'h854;
17'h166d8:	data_out=16'ha00;
17'h166d9:	data_out=16'h95a;
17'h166da:	data_out=16'ha00;
17'h166db:	data_out=16'h9ea;
17'h166dc:	data_out=16'ha00;
17'h166dd:	data_out=16'ha00;
17'h166de:	data_out=16'h9fd;
17'h166df:	data_out=16'h419;
17'h166e0:	data_out=16'h984;
17'h166e1:	data_out=16'h9f3;
17'h166e2:	data_out=16'h9a7;
17'h166e3:	data_out=16'h9fb;
17'h166e4:	data_out=16'h70f;
17'h166e5:	data_out=16'h296;
17'h166e6:	data_out=16'h5e7;
17'h166e7:	data_out=16'h9fb;
17'h166e8:	data_out=16'ha00;
17'h166e9:	data_out=16'ha00;
17'h166ea:	data_out=16'ha00;
17'h166eb:	data_out=16'h90a;
17'h166ec:	data_out=16'h9fe;
17'h166ed:	data_out=16'h9fc;
17'h166ee:	data_out=16'ha00;
17'h166ef:	data_out=16'h92b;
17'h166f0:	data_out=16'ha00;
17'h166f1:	data_out=16'h88c2;
17'h166f2:	data_out=16'h8dd;
17'h166f3:	data_out=16'h9ad;
17'h166f4:	data_out=16'ha00;
17'h166f5:	data_out=16'h9f6;
17'h166f6:	data_out=16'h9fa;
17'h166f7:	data_out=16'h996;
17'h166f8:	data_out=16'h8204;
17'h166f9:	data_out=16'ha00;
17'h166fa:	data_out=16'h9fa;
17'h166fb:	data_out=16'ha00;
17'h166fc:	data_out=16'h8973;
17'h166fd:	data_out=16'h89fe;
17'h166fe:	data_out=16'h894;
17'h166ff:	data_out=16'h9f2;
17'h16700:	data_out=16'h854c;
17'h16701:	data_out=16'h955;
17'h16702:	data_out=16'ha00;
17'h16703:	data_out=16'ha00;
17'h16704:	data_out=16'h8569;
17'h16705:	data_out=16'h94e;
17'h16706:	data_out=16'h1ac;
17'h16707:	data_out=16'h8a00;
17'h16708:	data_out=16'ha00;
17'h16709:	data_out=16'h82ed;
17'h1670a:	data_out=16'h803d;
17'h1670b:	data_out=16'ha00;
17'h1670c:	data_out=16'h86d0;
17'h1670d:	data_out=16'h821;
17'h1670e:	data_out=16'ha00;
17'h1670f:	data_out=16'h9c9;
17'h16710:	data_out=16'h9e7;
17'h16711:	data_out=16'h8033;
17'h16712:	data_out=16'ha00;
17'h16713:	data_out=16'h9da;
17'h16714:	data_out=16'h9ff;
17'h16715:	data_out=16'h85d3;
17'h16716:	data_out=16'h8289;
17'h16717:	data_out=16'h9ff;
17'h16718:	data_out=16'h87a4;
17'h16719:	data_out=16'h9f1;
17'h1671a:	data_out=16'h445;
17'h1671b:	data_out=16'ha00;
17'h1671c:	data_out=16'ha00;
17'h1671d:	data_out=16'h69d;
17'h1671e:	data_out=16'ha00;
17'h1671f:	data_out=16'h359;
17'h16720:	data_out=16'hbd;
17'h16721:	data_out=16'ha00;
17'h16722:	data_out=16'ha00;
17'h16723:	data_out=16'h89f1;
17'h16724:	data_out=16'h89f1;
17'h16725:	data_out=16'h399;
17'h16726:	data_out=16'ha00;
17'h16727:	data_out=16'h9f2;
17'h16728:	data_out=16'ha00;
17'h16729:	data_out=16'ha00;
17'h1672a:	data_out=16'h8bd;
17'h1672b:	data_out=16'h9f9;
17'h1672c:	data_out=16'h8598;
17'h1672d:	data_out=16'ha00;
17'h1672e:	data_out=16'h987;
17'h1672f:	data_out=16'h9fc;
17'h16730:	data_out=16'ha00;
17'h16731:	data_out=16'h89ff;
17'h16732:	data_out=16'h54d;
17'h16733:	data_out=16'ha00;
17'h16734:	data_out=16'h86ba;
17'h16735:	data_out=16'h900;
17'h16736:	data_out=16'ha00;
17'h16737:	data_out=16'ha00;
17'h16738:	data_out=16'h9ec;
17'h16739:	data_out=16'ha00;
17'h1673a:	data_out=16'h8a00;
17'h1673b:	data_out=16'h88b1;
17'h1673c:	data_out=16'ha00;
17'h1673d:	data_out=16'h45c;
17'h1673e:	data_out=16'ha00;
17'h1673f:	data_out=16'h94d;
17'h16740:	data_out=16'h8d6;
17'h16741:	data_out=16'ha00;
17'h16742:	data_out=16'h9ed;
17'h16743:	data_out=16'h8557;
17'h16744:	data_out=16'h806c;
17'h16745:	data_out=16'h85a2;
17'h16746:	data_out=16'ha00;
17'h16747:	data_out=16'h89e5;
17'h16748:	data_out=16'h9ef;
17'h16749:	data_out=16'h541;
17'h1674a:	data_out=16'h8960;
17'h1674b:	data_out=16'h4c9;
17'h1674c:	data_out=16'h85d0;
17'h1674d:	data_out=16'ha00;
17'h1674e:	data_out=16'ha00;
17'h1674f:	data_out=16'h89fc;
17'h16750:	data_out=16'h9a6;
17'h16751:	data_out=16'h9c3;
17'h16752:	data_out=16'h89ea;
17'h16753:	data_out=16'h9f9;
17'h16754:	data_out=16'h9f9;
17'h16755:	data_out=16'h9bc;
17'h16756:	data_out=16'ha00;
17'h16757:	data_out=16'h887;
17'h16758:	data_out=16'ha00;
17'h16759:	data_out=16'h836;
17'h1675a:	data_out=16'ha00;
17'h1675b:	data_out=16'h3aa;
17'h1675c:	data_out=16'ha00;
17'h1675d:	data_out=16'h9fb;
17'h1675e:	data_out=16'h9fb;
17'h1675f:	data_out=16'h8983;
17'h16760:	data_out=16'ha00;
17'h16761:	data_out=16'h995;
17'h16762:	data_out=16'h9fa;
17'h16763:	data_out=16'h9ff;
17'h16764:	data_out=16'h820a;
17'h16765:	data_out=16'h88d6;
17'h16766:	data_out=16'h8385;
17'h16767:	data_out=16'h90e;
17'h16768:	data_out=16'ha00;
17'h16769:	data_out=16'ha00;
17'h1676a:	data_out=16'ha00;
17'h1676b:	data_out=16'h249;
17'h1676c:	data_out=16'h840e;
17'h1676d:	data_out=16'ha00;
17'h1676e:	data_out=16'ha00;
17'h1676f:	data_out=16'h8d2;
17'h16770:	data_out=16'ha00;
17'h16771:	data_out=16'h89b6;
17'h16772:	data_out=16'h815;
17'h16773:	data_out=16'h8c9;
17'h16774:	data_out=16'ha00;
17'h16775:	data_out=16'h9ec;
17'h16776:	data_out=16'h9f5;
17'h16777:	data_out=16'h9fa;
17'h16778:	data_out=16'h19d;
17'h16779:	data_out=16'ha00;
17'h1677a:	data_out=16'ha00;
17'h1677b:	data_out=16'ha00;
17'h1677c:	data_out=16'h89df;
17'h1677d:	data_out=16'h89fc;
17'h1677e:	data_out=16'h9a3;
17'h1677f:	data_out=16'h2fe;
17'h16780:	data_out=16'h8950;
17'h16781:	data_out=16'h82bb;
17'h16782:	data_out=16'h9fd;
17'h16783:	data_out=16'ha00;
17'h16784:	data_out=16'h894c;
17'h16785:	data_out=16'h55a;
17'h16786:	data_out=16'h981;
17'h16787:	data_out=16'h8a00;
17'h16788:	data_out=16'ha00;
17'h16789:	data_out=16'h84bd;
17'h1678a:	data_out=16'h89f5;
17'h1678b:	data_out=16'ha00;
17'h1678c:	data_out=16'h86e9;
17'h1678d:	data_out=16'h5db;
17'h1678e:	data_out=16'h6cc;
17'h1678f:	data_out=16'h35d;
17'h16790:	data_out=16'h9f3;
17'h16791:	data_out=16'h876b;
17'h16792:	data_out=16'h893;
17'h16793:	data_out=16'h9fd;
17'h16794:	data_out=16'ha00;
17'h16795:	data_out=16'h86e4;
17'h16796:	data_out=16'h82a3;
17'h16797:	data_out=16'ha00;
17'h16798:	data_out=16'h89fc;
17'h16799:	data_out=16'h9ff;
17'h1679a:	data_out=16'h823e;
17'h1679b:	data_out=16'ha00;
17'h1679c:	data_out=16'ha00;
17'h1679d:	data_out=16'h88b6;
17'h1679e:	data_out=16'ha00;
17'h1679f:	data_out=16'h5a3;
17'h167a0:	data_out=16'h881e;
17'h167a1:	data_out=16'h744;
17'h167a2:	data_out=16'ha00;
17'h167a3:	data_out=16'h89f5;
17'h167a4:	data_out=16'h89f5;
17'h167a5:	data_out=16'h81d7;
17'h167a6:	data_out=16'h9ff;
17'h167a7:	data_out=16'h8768;
17'h167a8:	data_out=16'h908;
17'h167a9:	data_out=16'h9fa;
17'h167aa:	data_out=16'h86f1;
17'h167ab:	data_out=16'ha00;
17'h167ac:	data_out=16'h8509;
17'h167ad:	data_out=16'h9f9;
17'h167ae:	data_out=16'h392;
17'h167af:	data_out=16'h9fa;
17'h167b0:	data_out=16'h294;
17'h167b1:	data_out=16'h8838;
17'h167b2:	data_out=16'h81b0;
17'h167b3:	data_out=16'ha00;
17'h167b4:	data_out=16'h899b;
17'h167b5:	data_out=16'h3a0;
17'h167b6:	data_out=16'h9fc;
17'h167b7:	data_out=16'h9ff;
17'h167b8:	data_out=16'h8287;
17'h167b9:	data_out=16'ha00;
17'h167ba:	data_out=16'h8a00;
17'h167bb:	data_out=16'h877d;
17'h167bc:	data_out=16'ha00;
17'h167bd:	data_out=16'h8848;
17'h167be:	data_out=16'h913;
17'h167bf:	data_out=16'h52f;
17'h167c0:	data_out=16'hc5;
17'h167c1:	data_out=16'ha00;
17'h167c2:	data_out=16'h9f3;
17'h167c3:	data_out=16'h9af;
17'h167c4:	data_out=16'h81c8;
17'h167c5:	data_out=16'h86ba;
17'h167c6:	data_out=16'ha00;
17'h167c7:	data_out=16'h8a00;
17'h167c8:	data_out=16'h82df;
17'h167c9:	data_out=16'h800b;
17'h167ca:	data_out=16'h899f;
17'h167cb:	data_out=16'h12f;
17'h167cc:	data_out=16'h89fd;
17'h167cd:	data_out=16'ha00;
17'h167ce:	data_out=16'h83db;
17'h167cf:	data_out=16'h8a00;
17'h167d0:	data_out=16'h9ff;
17'h167d1:	data_out=16'h9f4;
17'h167d2:	data_out=16'h89ef;
17'h167d3:	data_out=16'h9fa;
17'h167d4:	data_out=16'h5f1;
17'h167d5:	data_out=16'h9e3;
17'h167d6:	data_out=16'ha00;
17'h167d7:	data_out=16'h8c5;
17'h167d8:	data_out=16'ha00;
17'h167d9:	data_out=16'h831a;
17'h167da:	data_out=16'ha00;
17'h167db:	data_out=16'h4b9;
17'h167dc:	data_out=16'h78c;
17'h167dd:	data_out=16'h316;
17'h167de:	data_out=16'h9fa;
17'h167df:	data_out=16'h89f4;
17'h167e0:	data_out=16'h9fb;
17'h167e1:	data_out=16'h249;
17'h167e2:	data_out=16'h9f6;
17'h167e3:	data_out=16'ha00;
17'h167e4:	data_out=16'h888e;
17'h167e5:	data_out=16'h8903;
17'h167e6:	data_out=16'h20a;
17'h167e7:	data_out=16'h659;
17'h167e8:	data_out=16'h7c3;
17'h167e9:	data_out=16'ha00;
17'h167ea:	data_out=16'h679;
17'h167eb:	data_out=16'h8340;
17'h167ec:	data_out=16'h89be;
17'h167ed:	data_out=16'ha00;
17'h167ee:	data_out=16'h679;
17'h167ef:	data_out=16'h9da;
17'h167f0:	data_out=16'h6a7;
17'h167f1:	data_out=16'h89ff;
17'h167f2:	data_out=16'h8028;
17'h167f3:	data_out=16'h31;
17'h167f4:	data_out=16'h2e5;
17'h167f5:	data_out=16'ha00;
17'h167f6:	data_out=16'h45c;
17'h167f7:	data_out=16'h9f5;
17'h167f8:	data_out=16'h9ea;
17'h167f9:	data_out=16'h86d2;
17'h167fa:	data_out=16'ha00;
17'h167fb:	data_out=16'h917;
17'h167fc:	data_out=16'h89fd;
17'h167fd:	data_out=16'h8402;
17'h167fe:	data_out=16'h9d6;
17'h167ff:	data_out=16'h845f;
17'h16800:	data_out=16'h89f6;
17'h16801:	data_out=16'h8a00;
17'h16802:	data_out=16'h9f7;
17'h16803:	data_out=16'ha00;
17'h16804:	data_out=16'h88ff;
17'h16805:	data_out=16'h94;
17'h16806:	data_out=16'h9ee;
17'h16807:	data_out=16'h8a00;
17'h16808:	data_out=16'h9aa;
17'h16809:	data_out=16'h9e9;
17'h1680a:	data_out=16'h8a00;
17'h1680b:	data_out=16'ha00;
17'h1680c:	data_out=16'h886d;
17'h1680d:	data_out=16'h5e3;
17'h1680e:	data_out=16'h410;
17'h1680f:	data_out=16'h284;
17'h16810:	data_out=16'ha00;
17'h16811:	data_out=16'h88a1;
17'h16812:	data_out=16'h7c2;
17'h16813:	data_out=16'ha00;
17'h16814:	data_out=16'ha00;
17'h16815:	data_out=16'h83cd;
17'h16816:	data_out=16'ha;
17'h16817:	data_out=16'ha00;
17'h16818:	data_out=16'h884c;
17'h16819:	data_out=16'h22d;
17'h1681a:	data_out=16'h86ab;
17'h1681b:	data_out=16'ha00;
17'h1681c:	data_out=16'ha00;
17'h1681d:	data_out=16'h8a00;
17'h1681e:	data_out=16'ha00;
17'h1681f:	data_out=16'h9a2;
17'h16820:	data_out=16'h89d1;
17'h16821:	data_out=16'h440;
17'h16822:	data_out=16'ha00;
17'h16823:	data_out=16'h89fe;
17'h16824:	data_out=16'h89fe;
17'h16825:	data_out=16'ha00;
17'h16826:	data_out=16'ha00;
17'h16827:	data_out=16'h896b;
17'h16828:	data_out=16'h514;
17'h16829:	data_out=16'h9ff;
17'h1682a:	data_out=16'h8a00;
17'h1682b:	data_out=16'h938;
17'h1682c:	data_out=16'h80ba;
17'h1682d:	data_out=16'h9f3;
17'h1682e:	data_out=16'h197;
17'h1682f:	data_out=16'h38e;
17'h16830:	data_out=16'h8483;
17'h16831:	data_out=16'h8928;
17'h16832:	data_out=16'h86a6;
17'h16833:	data_out=16'ha00;
17'h16834:	data_out=16'h8a00;
17'h16835:	data_out=16'h386;
17'h16836:	data_out=16'h5b9;
17'h16837:	data_out=16'h9f8;
17'h16838:	data_out=16'h89b8;
17'h16839:	data_out=16'ha00;
17'h1683a:	data_out=16'h89ff;
17'h1683b:	data_out=16'h8922;
17'h1683c:	data_out=16'ha00;
17'h1683d:	data_out=16'h88f4;
17'h1683e:	data_out=16'h51d;
17'h1683f:	data_out=16'h73;
17'h16840:	data_out=16'h9eb;
17'h16841:	data_out=16'ha00;
17'h16842:	data_out=16'h845;
17'h16843:	data_out=16'ha00;
17'h16844:	data_out=16'h83f4;
17'h16845:	data_out=16'h8395;
17'h16846:	data_out=16'ha00;
17'h16847:	data_out=16'h8a00;
17'h16848:	data_out=16'h87b3;
17'h16849:	data_out=16'ha00;
17'h1684a:	data_out=16'h8a00;
17'h1684b:	data_out=16'h86ad;
17'h1684c:	data_out=16'h8a00;
17'h1684d:	data_out=16'ha00;
17'h1684e:	data_out=16'h8623;
17'h1684f:	data_out=16'h8a00;
17'h16850:	data_out=16'ha00;
17'h16851:	data_out=16'h9ff;
17'h16852:	data_out=16'h89f8;
17'h16853:	data_out=16'h88aa;
17'h16854:	data_out=16'h89f7;
17'h16855:	data_out=16'h9fc;
17'h16856:	data_out=16'ha00;
17'h16857:	data_out=16'h9ff;
17'h16858:	data_out=16'ha00;
17'h16859:	data_out=16'h2c4;
17'h1685a:	data_out=16'ha00;
17'h1685b:	data_out=16'h81da;
17'h1685c:	data_out=16'h8462;
17'h1685d:	data_out=16'h89a4;
17'h1685e:	data_out=16'h690;
17'h1685f:	data_out=16'h8a00;
17'h16860:	data_out=16'h9fd;
17'h16861:	data_out=16'h8463;
17'h16862:	data_out=16'h9f9;
17'h16863:	data_out=16'ha00;
17'h16864:	data_out=16'h89f4;
17'h16865:	data_out=16'h866f;
17'h16866:	data_out=16'h230;
17'h16867:	data_out=16'h61f;
17'h16868:	data_out=16'h484;
17'h16869:	data_out=16'ha00;
17'h1686a:	data_out=16'h3fb;
17'h1686b:	data_out=16'h845a;
17'h1686c:	data_out=16'h8a00;
17'h1686d:	data_out=16'ha00;
17'h1686e:	data_out=16'h3fc;
17'h1686f:	data_out=16'h9de;
17'h16870:	data_out=16'h409;
17'h16871:	data_out=16'h8a00;
17'h16872:	data_out=16'h838e;
17'h16873:	data_out=16'h831d;
17'h16874:	data_out=16'h84a9;
17'h16875:	data_out=16'ha00;
17'h16876:	data_out=16'h380;
17'h16877:	data_out=16'h9fe;
17'h16878:	data_out=16'h9ff;
17'h16879:	data_out=16'h880c;
17'h1687a:	data_out=16'ha00;
17'h1687b:	data_out=16'h520;
17'h1687c:	data_out=16'h8a00;
17'h1687d:	data_out=16'h88b;
17'h1687e:	data_out=16'h9ff;
17'h1687f:	data_out=16'h86d4;
17'h16880:	data_out=16'h89b7;
17'h16881:	data_out=16'h8a00;
17'h16882:	data_out=16'h9f8;
17'h16883:	data_out=16'ha00;
17'h16884:	data_out=16'h8951;
17'h16885:	data_out=16'h8950;
17'h16886:	data_out=16'h98b;
17'h16887:	data_out=16'h8a00;
17'h16888:	data_out=16'h9fe;
17'h16889:	data_out=16'h9ed;
17'h1688a:	data_out=16'h8a00;
17'h1688b:	data_out=16'ha00;
17'h1688c:	data_out=16'h8687;
17'h1688d:	data_out=16'h6ef;
17'h1688e:	data_out=16'h222;
17'h1688f:	data_out=16'h61f;
17'h16890:	data_out=16'ha00;
17'h16891:	data_out=16'h89be;
17'h16892:	data_out=16'h9fa;
17'h16893:	data_out=16'h9ff;
17'h16894:	data_out=16'ha00;
17'h16895:	data_out=16'h8298;
17'h16896:	data_out=16'h1c;
17'h16897:	data_out=16'ha00;
17'h16898:	data_out=16'h8124;
17'h16899:	data_out=16'h88df;
17'h1689a:	data_out=16'h898d;
17'h1689b:	data_out=16'ha00;
17'h1689c:	data_out=16'h81ea;
17'h1689d:	data_out=16'h8a00;
17'h1689e:	data_out=16'h9ff;
17'h1689f:	data_out=16'h3ae;
17'h168a0:	data_out=16'h89bb;
17'h168a1:	data_out=16'h239;
17'h168a2:	data_out=16'h7ed;
17'h168a3:	data_out=16'h89e9;
17'h168a4:	data_out=16'h89e7;
17'h168a5:	data_out=16'h734;
17'h168a6:	data_out=16'h9fa;
17'h168a7:	data_out=16'h899f;
17'h168a8:	data_out=16'h29c;
17'h168a9:	data_out=16'ha00;
17'h168aa:	data_out=16'h45;
17'h168ab:	data_out=16'h8155;
17'h168ac:	data_out=16'h80ce;
17'h168ad:	data_out=16'h9f6;
17'h168ae:	data_out=16'h85e;
17'h168af:	data_out=16'h7d;
17'h168b0:	data_out=16'h8894;
17'h168b1:	data_out=16'h89cc;
17'h168b2:	data_out=16'h89c2;
17'h168b3:	data_out=16'ha00;
17'h168b4:	data_out=16'h8a00;
17'h168b5:	data_out=16'h84ba;
17'h168b6:	data_out=16'h9f8;
17'h168b7:	data_out=16'h9f9;
17'h168b8:	data_out=16'h89f8;
17'h168b9:	data_out=16'ha00;
17'h168ba:	data_out=16'h89fd;
17'h168bb:	data_out=16'h8960;
17'h168bc:	data_out=16'ha00;
17'h168bd:	data_out=16'h8945;
17'h168be:	data_out=16'h2a1;
17'h168bf:	data_out=16'h8950;
17'h168c0:	data_out=16'h48c;
17'h168c1:	data_out=16'ha00;
17'h168c2:	data_out=16'h823d;
17'h168c3:	data_out=16'h9ee;
17'h168c4:	data_out=16'h892e;
17'h168c5:	data_out=16'h827d;
17'h168c6:	data_out=16'ha00;
17'h168c7:	data_out=16'h89ff;
17'h168c8:	data_out=16'h8079;
17'h168c9:	data_out=16'h7e2;
17'h168ca:	data_out=16'h8a00;
17'h168cb:	data_out=16'h89fb;
17'h168cc:	data_out=16'h8a00;
17'h168cd:	data_out=16'h709;
17'h168ce:	data_out=16'h343;
17'h168cf:	data_out=16'h8a00;
17'h168d0:	data_out=16'h99e;
17'h168d1:	data_out=16'h9fc;
17'h168d2:	data_out=16'h8912;
17'h168d3:	data_out=16'h8951;
17'h168d4:	data_out=16'h89b8;
17'h168d5:	data_out=16'h9f4;
17'h168d6:	data_out=16'ha00;
17'h168d7:	data_out=16'h9f9;
17'h168d8:	data_out=16'ha00;
17'h168d9:	data_out=16'h812a;
17'h168da:	data_out=16'ha00;
17'h168db:	data_out=16'h893e;
17'h168dc:	data_out=16'h8852;
17'h168dd:	data_out=16'h898b;
17'h168de:	data_out=16'h269;
17'h168df:	data_out=16'h8a00;
17'h168e0:	data_out=16'h9f9;
17'h168e1:	data_out=16'h8965;
17'h168e2:	data_out=16'h9fb;
17'h168e3:	data_out=16'ha00;
17'h168e4:	data_out=16'h89e9;
17'h168e5:	data_out=16'h8a00;
17'h168e6:	data_out=16'h864b;
17'h168e7:	data_out=16'h5b5;
17'h168e8:	data_out=16'h25a;
17'h168e9:	data_out=16'h9ff;
17'h168ea:	data_out=16'h219;
17'h168eb:	data_out=16'h893e;
17'h168ec:	data_out=16'h89fa;
17'h168ed:	data_out=16'ha00;
17'h168ee:	data_out=16'h219;
17'h168ef:	data_out=16'h8629;
17'h168f0:	data_out=16'h21f;
17'h168f1:	data_out=16'h8a00;
17'h168f2:	data_out=16'h89d6;
17'h168f3:	data_out=16'h89d4;
17'h168f4:	data_out=16'h889d;
17'h168f5:	data_out=16'h9f9;
17'h168f6:	data_out=16'h80e1;
17'h168f7:	data_out=16'h9fc;
17'h168f8:	data_out=16'h9f2;
17'h168f9:	data_out=16'h4d1;
17'h168fa:	data_out=16'ha00;
17'h168fb:	data_out=16'h2a2;
17'h168fc:	data_out=16'h89a2;
17'h168fd:	data_out=16'h508;
17'h168fe:	data_out=16'h9f3;
17'h168ff:	data_out=16'h889e;
17'h16900:	data_out=16'h8902;
17'h16901:	data_out=16'h8a00;
17'h16902:	data_out=16'h9f9;
17'h16903:	data_out=16'h28e;
17'h16904:	data_out=16'h8958;
17'h16905:	data_out=16'h8996;
17'h16906:	data_out=16'h81ba;
17'h16907:	data_out=16'h8a00;
17'h16908:	data_out=16'h9fc;
17'h16909:	data_out=16'h623;
17'h1690a:	data_out=16'h89fc;
17'h1690b:	data_out=16'h9f8;
17'h1690c:	data_out=16'h85d7;
17'h1690d:	data_out=16'h331;
17'h1690e:	data_out=16'h1b3;
17'h1690f:	data_out=16'h57f;
17'h16910:	data_out=16'h9de;
17'h16911:	data_out=16'h89f8;
17'h16912:	data_out=16'h73c;
17'h16913:	data_out=16'h277;
17'h16914:	data_out=16'h9fb;
17'h16915:	data_out=16'h804e;
17'h16916:	data_out=16'hd9;
17'h16917:	data_out=16'h9f6;
17'h16918:	data_out=16'h301;
17'h16919:	data_out=16'h89fe;
17'h1691a:	data_out=16'h89cc;
17'h1691b:	data_out=16'ha00;
17'h1691c:	data_out=16'h8758;
17'h1691d:	data_out=16'h8a00;
17'h1691e:	data_out=16'h62c;
17'h1691f:	data_out=16'h829e;
17'h16920:	data_out=16'h89b4;
17'h16921:	data_out=16'h1b3;
17'h16922:	data_out=16'h50;
17'h16923:	data_out=16'h843b;
17'h16924:	data_out=16'h8435;
17'h16925:	data_out=16'h811a;
17'h16926:	data_out=16'h9f8;
17'h16927:	data_out=16'h89c4;
17'h16928:	data_out=16'h1d5;
17'h16929:	data_out=16'h301;
17'h1692a:	data_out=16'h698;
17'h1692b:	data_out=16'h84e0;
17'h1692c:	data_out=16'h46;
17'h1692d:	data_out=16'h9f5;
17'h1692e:	data_out=16'h912;
17'h1692f:	data_out=16'h83aa;
17'h16930:	data_out=16'h8986;
17'h16931:	data_out=16'h89ee;
17'h16932:	data_out=16'h89ee;
17'h16933:	data_out=16'h8a0;
17'h16934:	data_out=16'h8a00;
17'h16935:	data_out=16'h84f0;
17'h16936:	data_out=16'h9f6;
17'h16937:	data_out=16'h9e1;
17'h16938:	data_out=16'h8a00;
17'h16939:	data_out=16'h7c0;
17'h1693a:	data_out=16'h89fd;
17'h1693b:	data_out=16'h8744;
17'h1693c:	data_out=16'ha00;
17'h1693d:	data_out=16'h896d;
17'h1693e:	data_out=16'h1d7;
17'h1693f:	data_out=16'h8992;
17'h16940:	data_out=16'h837b;
17'h16941:	data_out=16'ha00;
17'h16942:	data_out=16'h88eb;
17'h16943:	data_out=16'h287;
17'h16944:	data_out=16'h866a;
17'h16945:	data_out=16'h8046;
17'h16946:	data_out=16'ha00;
17'h16947:	data_out=16'h8a00;
17'h16948:	data_out=16'h8069;
17'h16949:	data_out=16'h8155;
17'h1694a:	data_out=16'h8a00;
17'h1694b:	data_out=16'h8a00;
17'h1694c:	data_out=16'h8a00;
17'h1694d:	data_out=16'ha;
17'h1694e:	data_out=16'h5c3;
17'h1694f:	data_out=16'h8a00;
17'h16950:	data_out=16'h161;
17'h16951:	data_out=16'h9ff;
17'h16952:	data_out=16'h841e;
17'h16953:	data_out=16'h89bf;
17'h16954:	data_out=16'h855a;
17'h16955:	data_out=16'h9fc;
17'h16956:	data_out=16'h61c;
17'h16957:	data_out=16'h5fb;
17'h16958:	data_out=16'ha00;
17'h16959:	data_out=16'h8545;
17'h1695a:	data_out=16'ha00;
17'h1695b:	data_out=16'h87cb;
17'h1695c:	data_out=16'h8975;
17'h1695d:	data_out=16'h84f1;
17'h1695e:	data_out=16'h8360;
17'h1695f:	data_out=16'h85f1;
17'h16960:	data_out=16'h433;
17'h16961:	data_out=16'h89aa;
17'h16962:	data_out=16'h9ee;
17'h16963:	data_out=16'h8f0;
17'h16964:	data_out=16'h89f2;
17'h16965:	data_out=16'h89fd;
17'h16966:	data_out=16'h89fd;
17'h16967:	data_out=16'h1f7;
17'h16968:	data_out=16'h1bb;
17'h16969:	data_out=16'h9fb;
17'h1696a:	data_out=16'h1b7;
17'h1696b:	data_out=16'h89d7;
17'h1696c:	data_out=16'h89a2;
17'h1696d:	data_out=16'h89c;
17'h1696e:	data_out=16'h1b7;
17'h1696f:	data_out=16'h89f6;
17'h16970:	data_out=16'h1b6;
17'h16971:	data_out=16'h84eb;
17'h16972:	data_out=16'h89fa;
17'h16973:	data_out=16'h89fb;
17'h16974:	data_out=16'h8980;
17'h16975:	data_out=16'ha00;
17'h16976:	data_out=16'h837d;
17'h16977:	data_out=16'h9f8;
17'h16978:	data_out=16'h808d;
17'h16979:	data_out=16'h9c9;
17'h1697a:	data_out=16'h9fb;
17'h1697b:	data_out=16'h1d8;
17'h1697c:	data_out=16'h81eb;
17'h1697d:	data_out=16'h817a;
17'h1697e:	data_out=16'h9d8;
17'h1697f:	data_out=16'h8765;
17'h16980:	data_out=16'h8462;
17'h16981:	data_out=16'h887f;
17'h16982:	data_out=16'h660;
17'h16983:	data_out=16'h8169;
17'h16984:	data_out=16'h878b;
17'h16985:	data_out=16'h8373;
17'h16986:	data_out=16'h81e1;
17'h16987:	data_out=16'h82bd;
17'h16988:	data_out=16'ha00;
17'h16989:	data_out=16'h34d;
17'h1698a:	data_out=16'h86b4;
17'h1698b:	data_out=16'h4da;
17'h1698c:	data_out=16'h803b;
17'h1698d:	data_out=16'h80dc;
17'h1698e:	data_out=16'h14f;
17'h1698f:	data_out=16'h3ed;
17'h16990:	data_out=16'hbc;
17'h16991:	data_out=16'h8984;
17'h16992:	data_out=16'h84;
17'h16993:	data_out=16'h822c;
17'h16994:	data_out=16'h19d;
17'h16995:	data_out=16'h1ac;
17'h16996:	data_out=16'h2b8;
17'h16997:	data_out=16'h809f;
17'h16998:	data_out=16'h3e3;
17'h16999:	data_out=16'h8838;
17'h1699a:	data_out=16'h8924;
17'h1699b:	data_out=16'h86a4;
17'h1699c:	data_out=16'h8365;
17'h1699d:	data_out=16'h8a00;
17'h1699e:	data_out=16'h809a;
17'h1699f:	data_out=16'h5c0;
17'h169a0:	data_out=16'h89f5;
17'h169a1:	data_out=16'h148;
17'h169a2:	data_out=16'h8228;
17'h169a3:	data_out=16'hd9;
17'h169a4:	data_out=16'hdb;
17'h169a5:	data_out=16'h81ae;
17'h169a6:	data_out=16'h78d;
17'h169a7:	data_out=16'h89ee;
17'h169a8:	data_out=16'h148;
17'h169a9:	data_out=16'h829c;
17'h169aa:	data_out=16'h3a9;
17'h169ab:	data_out=16'h8674;
17'h169ac:	data_out=16'h287;
17'h169ad:	data_out=16'h820f;
17'h169ae:	data_out=16'h581;
17'h169af:	data_out=16'h894d;
17'h169b0:	data_out=16'h87f5;
17'h169b1:	data_out=16'h89ef;
17'h169b2:	data_out=16'h8906;
17'h169b3:	data_out=16'h122;
17'h169b4:	data_out=16'h8a00;
17'h169b5:	data_out=16'he6;
17'h169b6:	data_out=16'h47d;
17'h169b7:	data_out=16'h5ad;
17'h169b8:	data_out=16'h8a00;
17'h169b9:	data_out=16'h99;
17'h169ba:	data_out=16'h8196;
17'h169bb:	data_out=16'ha5;
17'h169bc:	data_out=16'h72e;
17'h169bd:	data_out=16'h83a0;
17'h169be:	data_out=16'h148;
17'h169bf:	data_out=16'h8367;
17'h169c0:	data_out=16'hdb;
17'h169c1:	data_out=16'ha00;
17'h169c2:	data_out=16'h88a0;
17'h169c3:	data_out=16'h110;
17'h169c4:	data_out=16'h80b3;
17'h169c5:	data_out=16'h1bd;
17'h169c6:	data_out=16'h3a;
17'h169c7:	data_out=16'h826e;
17'h169c8:	data_out=16'h82e7;
17'h169c9:	data_out=16'h818c;
17'h169ca:	data_out=16'h8471;
17'h169cb:	data_out=16'h8a00;
17'h169cc:	data_out=16'h863d;
17'h169cd:	data_out=16'h828e;
17'h169ce:	data_out=16'h8098;
17'h169cf:	data_out=16'h8555;
17'h169d0:	data_out=16'h334;
17'h169d1:	data_out=16'ha00;
17'h169d2:	data_out=16'h1a5;
17'h169d3:	data_out=16'h8a00;
17'h169d4:	data_out=16'h8705;
17'h169d5:	data_out=16'ha00;
17'h169d6:	data_out=16'h563;
17'h169d7:	data_out=16'h517;
17'h169d8:	data_out=16'ha00;
17'h169d9:	data_out=16'h12d;
17'h169da:	data_out=16'h82ae;
17'h169db:	data_out=16'h12a;
17'h169dc:	data_out=16'h88e6;
17'h169dd:	data_out=16'h841f;
17'h169de:	data_out=16'h8925;
17'h169df:	data_out=16'h82c7;
17'h169e0:	data_out=16'h241;
17'h169e1:	data_out=16'h8126;
17'h169e2:	data_out=16'h122;
17'h169e3:	data_out=16'hf3;
17'h169e4:	data_out=16'h89ff;
17'h169e5:	data_out=16'h8a00;
17'h169e6:	data_out=16'h8617;
17'h169e7:	data_out=16'h104;
17'h169e8:	data_out=16'h146;
17'h169e9:	data_out=16'ha00;
17'h169ea:	data_out=16'h158;
17'h169eb:	data_out=16'h873a;
17'h169ec:	data_out=16'h898d;
17'h169ed:	data_out=16'hd3;
17'h169ee:	data_out=16'h157;
17'h169ef:	data_out=16'h8882;
17'h169f0:	data_out=16'h154;
17'h169f1:	data_out=16'h2b8;
17'h169f2:	data_out=16'h8747;
17'h169f3:	data_out=16'h8864;
17'h169f4:	data_out=16'h87ca;
17'h169f5:	data_out=16'h49c;
17'h169f6:	data_out=16'h832d;
17'h169f7:	data_out=16'h88d;
17'h169f8:	data_out=16'h8217;
17'h169f9:	data_out=16'h531;
17'h169fa:	data_out=16'h15f;
17'h169fb:	data_out=16'h148;
17'h169fc:	data_out=16'h9f;
17'h169fd:	data_out=16'h803f;
17'h169fe:	data_out=16'h2bf;
17'h169ff:	data_out=16'h2a1;
17'h16a00:	data_out=16'h1a9;
17'h16a01:	data_out=16'hc7;
17'h16a02:	data_out=16'h33b;
17'h16a03:	data_out=16'h8205;
17'h16a04:	data_out=16'h81db;
17'h16a05:	data_out=16'h810c;
17'h16a06:	data_out=16'h8474;
17'h16a07:	data_out=16'h8321;
17'h16a08:	data_out=16'h5f5;
17'h16a09:	data_out=16'h81a0;
17'h16a0a:	data_out=16'h41;
17'h16a0b:	data_out=16'h836e;
17'h16a0c:	data_out=16'h19e;
17'h16a0d:	data_out=16'h81e0;
17'h16a0e:	data_out=16'h10;
17'h16a0f:	data_out=16'haf;
17'h16a10:	data_out=16'h6d;
17'h16a11:	data_out=16'h82ce;
17'h16a12:	data_out=16'h8477;
17'h16a13:	data_out=16'h838e;
17'h16a14:	data_out=16'h81f9;
17'h16a15:	data_out=16'h116;
17'h16a16:	data_out=16'h19b;
17'h16a17:	data_out=16'h8369;
17'h16a18:	data_out=16'h156;
17'h16a19:	data_out=16'h83b8;
17'h16a1a:	data_out=16'h8302;
17'h16a1b:	data_out=16'h8500;
17'h16a1c:	data_out=16'h80cb;
17'h16a1d:	data_out=16'h8127;
17'h16a1e:	data_out=16'h81ed;
17'h16a1f:	data_out=16'h8012;
17'h16a20:	data_out=16'h80cb;
17'h16a21:	data_out=16'h8;
17'h16a22:	data_out=16'h8241;
17'h16a23:	data_out=16'h1c1;
17'h16a24:	data_out=16'h1c5;
17'h16a25:	data_out=16'h8324;
17'h16a26:	data_out=16'h64;
17'h16a27:	data_out=16'h80f1;
17'h16a28:	data_out=16'h1;
17'h16a29:	data_out=16'h82e5;
17'h16a2a:	data_out=16'h8120;
17'h16a2b:	data_out=16'h82cb;
17'h16a2c:	data_out=16'h176;
17'h16a2d:	data_out=16'h83fb;
17'h16a2e:	data_out=16'h15a;
17'h16a2f:	data_out=16'h8274;
17'h16a30:	data_out=16'h8256;
17'h16a31:	data_out=16'h8648;
17'h16a32:	data_out=16'h82f7;
17'h16a33:	data_out=16'h819a;
17'h16a34:	data_out=16'h8652;
17'h16a35:	data_out=16'h2be;
17'h16a36:	data_out=16'h478;
17'h16a37:	data_out=16'h179;
17'h16a38:	data_out=16'h8470;
17'h16a39:	data_out=16'h8169;
17'h16a3a:	data_out=16'h8211;
17'h16a3b:	data_out=16'h278;
17'h16a3c:	data_out=16'h359;
17'h16a3d:	data_out=16'h8072;
17'h16a3e:	data_out=16'h6;
17'h16a3f:	data_out=16'h8101;
17'h16a40:	data_out=16'h825e;
17'h16a41:	data_out=16'h552;
17'h16a42:	data_out=16'h8421;
17'h16a43:	data_out=16'h82bc;
17'h16a44:	data_out=16'h109;
17'h16a45:	data_out=16'h165;
17'h16a46:	data_out=16'h8034;
17'h16a47:	data_out=16'h836b;
17'h16a48:	data_out=16'h8296;
17'h16a49:	data_out=16'h831c;
17'h16a4a:	data_out=16'h8182;
17'h16a4b:	data_out=16'h84e2;
17'h16a4c:	data_out=16'h83e3;
17'h16a4d:	data_out=16'h8244;
17'h16a4e:	data_out=16'h81cc;
17'h16a4f:	data_out=16'h83cb;
17'h16a50:	data_out=16'h8192;
17'h16a51:	data_out=16'h490;
17'h16a52:	data_out=16'h13d;
17'h16a53:	data_out=16'h84f5;
17'h16a54:	data_out=16'h801f;
17'h16a55:	data_out=16'h7ca;
17'h16a56:	data_out=16'h808e;
17'h16a57:	data_out=16'h5e;
17'h16a58:	data_out=16'h7f9;
17'h16a59:	data_out=16'h8013;
17'h16a5a:	data_out=16'h820b;
17'h16a5b:	data_out=16'h406;
17'h16a5c:	data_out=16'h80e1;
17'h16a5d:	data_out=16'h35;
17'h16a5e:	data_out=16'h82b3;
17'h16a5f:	data_out=16'h15;
17'h16a60:	data_out=16'h8152;
17'h16a61:	data_out=16'h212;
17'h16a62:	data_out=16'h8344;
17'h16a63:	data_out=16'h81b1;
17'h16a64:	data_out=16'h85b1;
17'h16a65:	data_out=16'h871f;
17'h16a66:	data_out=16'h8396;
17'h16a67:	data_out=16'h81d0;
17'h16a68:	data_out=16'h2;
17'h16a69:	data_out=16'h5af;
17'h16a6a:	data_out=16'h8;
17'h16a6b:	data_out=16'h8225;
17'h16a6c:	data_out=16'ha0;
17'h16a6d:	data_out=16'h81af;
17'h16a6e:	data_out=16'h1d;
17'h16a6f:	data_out=16'h84ee;
17'h16a70:	data_out=16'h17;
17'h16a71:	data_out=16'h194;
17'h16a72:	data_out=16'h81b0;
17'h16a73:	data_out=16'h836b;
17'h16a74:	data_out=16'h823a;
17'h16a75:	data_out=16'h80be;
17'h16a76:	data_out=16'h829d;
17'h16a77:	data_out=16'h80a3;
17'h16a78:	data_out=16'h8569;
17'h16a79:	data_out=16'h30a;
17'h16a7a:	data_out=16'h81c1;
17'h16a7b:	data_out=16'h4;
17'h16a7c:	data_out=16'h176;
17'h16a7d:	data_out=16'h848d;
17'h16a7e:	data_out=16'h81f8;
17'h16a7f:	data_out=16'h15e;
17'h16a80:	data_out=16'h7c;
17'h16a81:	data_out=16'h8060;
17'h16a82:	data_out=16'h8039;
17'h16a83:	data_out=16'h8039;
17'h16a84:	data_out=16'h80a0;
17'h16a85:	data_out=16'h8090;
17'h16a86:	data_out=16'h8075;
17'h16a87:	data_out=16'h803a;
17'h16a88:	data_out=16'h3c;
17'h16a89:	data_out=16'hb9;
17'h16a8a:	data_out=16'h809b;
17'h16a8b:	data_out=16'h3c;
17'h16a8c:	data_out=16'h80bb;
17'h16a8d:	data_out=16'h11;
17'h16a8e:	data_out=16'h801d;
17'h16a8f:	data_out=16'h1;
17'h16a90:	data_out=16'h2e;
17'h16a91:	data_out=16'h8074;
17'h16a92:	data_out=16'h8085;
17'h16a93:	data_out=16'h4b;
17'h16a94:	data_out=16'h805b;
17'h16a95:	data_out=16'h2d;
17'h16a96:	data_out=16'h2a;
17'h16a97:	data_out=16'h8055;
17'h16a98:	data_out=16'h801d;
17'h16a99:	data_out=16'h5e;
17'h16a9a:	data_out=16'h8095;
17'h16a9b:	data_out=16'he;
17'h16a9c:	data_out=16'h8072;
17'h16a9d:	data_out=16'h809c;
17'h16a9e:	data_out=16'h8025;
17'h16a9f:	data_out=16'h807e;
17'h16aa0:	data_out=16'h808c;
17'h16aa1:	data_out=16'h8021;
17'h16aa2:	data_out=16'h22;
17'h16aa3:	data_out=16'h80d6;
17'h16aa4:	data_out=16'h80de;
17'h16aa5:	data_out=16'h802d;
17'h16aa6:	data_out=16'had;
17'h16aa7:	data_out=16'h808a;
17'h16aa8:	data_out=16'h8023;
17'h16aa9:	data_out=16'hd;
17'h16aaa:	data_out=16'h8003;
17'h16aab:	data_out=16'h42;
17'h16aac:	data_out=16'h802d;
17'h16aad:	data_out=16'h8014;
17'h16aae:	data_out=16'h8014;
17'h16aaf:	data_out=16'h8033;
17'h16ab0:	data_out=16'h80e8;
17'h16ab1:	data_out=16'h800a;
17'h16ab2:	data_out=16'h80eb;
17'h16ab3:	data_out=16'h8047;
17'h16ab4:	data_out=16'h804f;
17'h16ab5:	data_out=16'h8108;
17'h16ab6:	data_out=16'h8072;
17'h16ab7:	data_out=16'h8072;
17'h16ab8:	data_out=16'h805c;
17'h16ab9:	data_out=16'h25;
17'h16aba:	data_out=16'h8078;
17'h16abb:	data_out=16'h10;
17'h16abc:	data_out=16'h8036;
17'h16abd:	data_out=16'h66;
17'h16abe:	data_out=16'h8023;
17'h16abf:	data_out=16'h8082;
17'h16ac0:	data_out=16'h80a3;
17'h16ac1:	data_out=16'h8030;
17'h16ac2:	data_out=16'h806c;
17'h16ac3:	data_out=16'h801e;
17'h16ac4:	data_out=16'h800b;
17'h16ac5:	data_out=16'h42;
17'h16ac6:	data_out=16'h803c;
17'h16ac7:	data_out=16'h80a8;
17'h16ac8:	data_out=16'h8036;
17'h16ac9:	data_out=16'h8013;
17'h16aca:	data_out=16'h80e4;
17'h16acb:	data_out=16'h80fa;
17'h16acc:	data_out=16'h80c4;
17'h16acd:	data_out=16'h31;
17'h16ace:	data_out=16'h8052;
17'h16acf:	data_out=16'h80ca;
17'h16ad0:	data_out=16'h8097;
17'h16ad1:	data_out=16'h18;
17'h16ad2:	data_out=16'h80ac;
17'h16ad3:	data_out=16'h80a9;
17'h16ad4:	data_out=16'h806b;
17'h16ad5:	data_out=16'h8028;
17'h16ad6:	data_out=16'h8058;
17'h16ad7:	data_out=16'h8016;
17'h16ad8:	data_out=16'h801c;
17'h16ad9:	data_out=16'h805b;
17'h16ada:	data_out=16'h802c;
17'h16adb:	data_out=16'h810c;
17'h16adc:	data_out=16'h8098;
17'h16add:	data_out=16'h8032;
17'h16ade:	data_out=16'h8039;
17'h16adf:	data_out=16'h8038;
17'h16ae0:	data_out=16'h22;
17'h16ae1:	data_out=16'h807b;
17'h16ae2:	data_out=16'h8032;
17'h16ae3:	data_out=16'h8059;
17'h16ae4:	data_out=16'h8025;
17'h16ae5:	data_out=16'h8023;
17'h16ae6:	data_out=16'h1c;
17'h16ae7:	data_out=16'h8050;
17'h16ae8:	data_out=16'h8025;
17'h16ae9:	data_out=16'h805d;
17'h16aea:	data_out=16'h802b;
17'h16aeb:	data_out=16'h801f;
17'h16aec:	data_out=16'h80c8;
17'h16aed:	data_out=16'h8048;
17'h16aee:	data_out=16'h8021;
17'h16aef:	data_out=16'h8060;
17'h16af0:	data_out=16'h801c;
17'h16af1:	data_out=16'h8069;
17'h16af2:	data_out=16'h805b;
17'h16af3:	data_out=16'h803f;
17'h16af4:	data_out=16'h80e0;
17'h16af5:	data_out=16'h8050;
17'h16af6:	data_out=16'h5c;
17'h16af7:	data_out=16'h802e;
17'h16af8:	data_out=16'h4c;
17'h16af9:	data_out=16'h805a;
17'h16afa:	data_out=16'h805a;
17'h16afb:	data_out=16'h8023;
17'h16afc:	data_out=16'h8035;
17'h16afd:	data_out=16'h8094;
17'h16afe:	data_out=16'hd4;
17'h16aff:	data_out=16'h8090;
17'h16b00:	data_out=16'h105;
17'h16b01:	data_out=16'hd;
17'h16b02:	data_out=16'h8084;
17'h16b03:	data_out=16'h801f;
17'h16b04:	data_out=16'h2;
17'h16b05:	data_out=16'h8006;
17'h16b06:	data_out=16'h8070;
17'h16b07:	data_out=16'h11;
17'h16b08:	data_out=16'h59;
17'h16b09:	data_out=16'had;
17'h16b0a:	data_out=16'h802d;
17'h16b0b:	data_out=16'h805d;
17'h16b0c:	data_out=16'h8039;
17'h16b0d:	data_out=16'h60;
17'h16b0e:	data_out=16'h8023;
17'h16b0f:	data_out=16'h23;
17'h16b10:	data_out=16'h8035;
17'h16b11:	data_out=16'h4e;
17'h16b12:	data_out=16'h8096;
17'h16b13:	data_out=16'h6d;
17'h16b14:	data_out=16'h8072;
17'h16b15:	data_out=16'h9a;
17'h16b16:	data_out=16'h8c;
17'h16b17:	data_out=16'h807c;
17'h16b18:	data_out=16'h8007;
17'h16b19:	data_out=16'hcc;
17'h16b1a:	data_out=16'h1c;
17'h16b1b:	data_out=16'h31;
17'h16b1c:	data_out=16'h38;
17'h16b1d:	data_out=16'h803e;
17'h16b1e:	data_out=16'h0;
17'h16b1f:	data_out=16'h804f;
17'h16b20:	data_out=16'h2b;
17'h16b21:	data_out=16'h801f;
17'h16b22:	data_out=16'h17;
17'h16b23:	data_out=16'h8090;
17'h16b24:	data_out=16'h8096;
17'h16b25:	data_out=16'h8034;
17'h16b26:	data_out=16'h68;
17'h16b27:	data_out=16'h8036;
17'h16b28:	data_out=16'h8022;
17'h16b29:	data_out=16'h9;
17'h16b2a:	data_out=16'h802a;
17'h16b2b:	data_out=16'h93;
17'h16b2c:	data_out=16'h6;
17'h16b2d:	data_out=16'h8051;
17'h16b2e:	data_out=16'h8086;
17'h16b2f:	data_out=16'he;
17'h16b30:	data_out=16'h803a;
17'h16b31:	data_out=16'he9;
17'h16b32:	data_out=16'h8027;
17'h16b33:	data_out=16'h803b;
17'h16b34:	data_out=16'h94;
17'h16b35:	data_out=16'h8070;
17'h16b36:	data_out=16'h809f;
17'h16b37:	data_out=16'h808c;
17'h16b38:	data_out=16'hb6;
17'h16b39:	data_out=16'h29;
17'h16b3a:	data_out=16'h8070;
17'h16b3b:	data_out=16'hb3;
17'h16b3c:	data_out=16'h80bb;
17'h16b3d:	data_out=16'hee;
17'h16b3e:	data_out=16'h8022;
17'h16b3f:	data_out=16'h11;
17'h16b40:	data_out=16'h8064;
17'h16b41:	data_out=16'h8069;
17'h16b42:	data_out=16'h8045;
17'h16b43:	data_out=16'h805f;
17'h16b44:	data_out=16'h3e;
17'h16b45:	data_out=16'h93;
17'h16b46:	data_out=16'h8063;
17'h16b47:	data_out=16'h807c;
17'h16b48:	data_out=16'h806a;
17'h16b49:	data_out=16'h8016;
17'h16b4a:	data_out=16'h804d;
17'h16b4b:	data_out=16'h8094;
17'h16b4c:	data_out=16'h8073;
17'h16b4d:	data_out=16'h4f;
17'h16b4e:	data_out=16'h7;
17'h16b4f:	data_out=16'h806c;
17'h16b50:	data_out=16'h806d;
17'h16b51:	data_out=16'h57;
17'h16b52:	data_out=16'h805d;
17'h16b53:	data_out=16'h801e;
17'h16b54:	data_out=16'h801a;
17'h16b55:	data_out=16'h80b3;
17'h16b56:	data_out=16'h8071;
17'h16b57:	data_out=16'h807f;
17'h16b58:	data_out=16'h80b9;
17'h16b59:	data_out=16'h808d;
17'h16b5a:	data_out=16'h80a1;
17'h16b5b:	data_out=16'h803d;
17'h16b5c:	data_out=16'h8016;
17'h16b5d:	data_out=16'h8002;
17'h16b5e:	data_out=16'h8012;
17'h16b5f:	data_out=16'h801d;
17'h16b60:	data_out=16'h2e;
17'h16b61:	data_out=16'h55;
17'h16b62:	data_out=16'h8078;
17'h16b63:	data_out=16'h804b;
17'h16b64:	data_out=16'h5b;
17'h16b65:	data_out=16'h12;
17'h16b66:	data_out=16'h6d;
17'h16b67:	data_out=16'h808e;
17'h16b68:	data_out=16'h8014;
17'h16b69:	data_out=16'h809e;
17'h16b6a:	data_out=16'h8019;
17'h16b6b:	data_out=16'hc0;
17'h16b6c:	data_out=16'h807c;
17'h16b6d:	data_out=16'h803f;
17'h16b6e:	data_out=16'h8016;
17'h16b6f:	data_out=16'h8;
17'h16b70:	data_out=16'h801c;
17'h16b71:	data_out=16'h8065;
17'h16b72:	data_out=16'h9;
17'h16b73:	data_out=16'h5d;
17'h16b74:	data_out=16'h802b;
17'h16b75:	data_out=16'h8019;
17'h16b76:	data_out=16'hac;
17'h16b77:	data_out=16'h804c;
17'h16b78:	data_out=16'h80;
17'h16b79:	data_out=16'h808e;
17'h16b7a:	data_out=16'h8076;
17'h16b7b:	data_out=16'h8015;
17'h16b7c:	data_out=16'h804e;
17'h16b7d:	data_out=16'h806d;
17'h16b7e:	data_out=16'haa;
17'h16b7f:	data_out=16'h804b;
17'h16b80:	data_out=16'h8009;
17'h16b81:	data_out=16'h7;
17'h16b82:	data_out=16'h8001;
17'h16b83:	data_out=16'h8000;
17'h16b84:	data_out=16'h8008;
17'h16b85:	data_out=16'h8004;
17'h16b86:	data_out=16'h8007;
17'h16b87:	data_out=16'h8008;
17'h16b88:	data_out=16'h1;
17'h16b89:	data_out=16'h8;
17'h16b8a:	data_out=16'h8000;
17'h16b8b:	data_out=16'h3;
17'h16b8c:	data_out=16'h8005;
17'h16b8d:	data_out=16'h8000;
17'h16b8e:	data_out=16'h8007;
17'h16b8f:	data_out=16'h6;
17'h16b90:	data_out=16'h6;
17'h16b91:	data_out=16'h5;
17'h16b92:	data_out=16'h8009;
17'h16b93:	data_out=16'h6;
17'h16b94:	data_out=16'h8008;
17'h16b95:	data_out=16'h4;
17'h16b96:	data_out=16'h8004;
17'h16b97:	data_out=16'h0;
17'h16b98:	data_out=16'h8001;
17'h16b99:	data_out=16'h1;
17'h16b9a:	data_out=16'h8002;
17'h16b9b:	data_out=16'h8002;
17'h16b9c:	data_out=16'h7;
17'h16b9d:	data_out=16'h8003;
17'h16b9e:	data_out=16'h8007;
17'h16b9f:	data_out=16'h8;
17'h16ba0:	data_out=16'h8006;
17'h16ba1:	data_out=16'h1;
17'h16ba2:	data_out=16'h8001;
17'h16ba3:	data_out=16'h8004;
17'h16ba4:	data_out=16'h6;
17'h16ba5:	data_out=16'h1;
17'h16ba6:	data_out=16'h8003;
17'h16ba7:	data_out=16'h8002;
17'h16ba8:	data_out=16'h8000;
17'h16ba9:	data_out=16'h6;
17'h16baa:	data_out=16'h8008;
17'h16bab:	data_out=16'h4;
17'h16bac:	data_out=16'h8004;
17'h16bad:	data_out=16'h8007;
17'h16bae:	data_out=16'h1;
17'h16baf:	data_out=16'h8007;
17'h16bb0:	data_out=16'h8;
17'h16bb1:	data_out=16'h1;
17'h16bb2:	data_out=16'h9;
17'h16bb3:	data_out=16'h8009;
17'h16bb4:	data_out=16'h8004;
17'h16bb5:	data_out=16'h8005;
17'h16bb6:	data_out=16'h0;
17'h16bb7:	data_out=16'h4;
17'h16bb8:	data_out=16'h5;
17'h16bb9:	data_out=16'h7;
17'h16bba:	data_out=16'h8007;
17'h16bbb:	data_out=16'h4;
17'h16bbc:	data_out=16'h8005;
17'h16bbd:	data_out=16'h8004;
17'h16bbe:	data_out=16'h2;
17'h16bbf:	data_out=16'h8002;
17'h16bc0:	data_out=16'h6;
17'h16bc1:	data_out=16'h8008;
17'h16bc2:	data_out=16'h3;
17'h16bc3:	data_out=16'h3;
17'h16bc4:	data_out=16'h2;
17'h16bc5:	data_out=16'h9;
17'h16bc6:	data_out=16'h8008;
17'h16bc7:	data_out=16'h8008;
17'h16bc8:	data_out=16'h5;
17'h16bc9:	data_out=16'h8008;
17'h16bca:	data_out=16'h5;
17'h16bcb:	data_out=16'h8007;
17'h16bcc:	data_out=16'h8005;
17'h16bcd:	data_out=16'h8003;
17'h16bce:	data_out=16'h8005;
17'h16bcf:	data_out=16'h8006;
17'h16bd0:	data_out=16'h7;
17'h16bd1:	data_out=16'h8005;
17'h16bd2:	data_out=16'h8006;
17'h16bd3:	data_out=16'h8006;
17'h16bd4:	data_out=16'h8001;
17'h16bd5:	data_out=16'h3;
17'h16bd6:	data_out=16'h7;
17'h16bd7:	data_out=16'h8005;
17'h16bd8:	data_out=16'h1;
17'h16bd9:	data_out=16'h8009;
17'h16bda:	data_out=16'h8;
17'h16bdb:	data_out=16'h5;
17'h16bdc:	data_out=16'h8004;
17'h16bdd:	data_out=16'h1;
17'h16bde:	data_out=16'h8005;
17'h16bdf:	data_out=16'h8007;
17'h16be0:	data_out=16'h2;
17'h16be1:	data_out=16'h7;
17'h16be2:	data_out=16'h5;
17'h16be3:	data_out=16'h8005;
17'h16be4:	data_out=16'h7;
17'h16be5:	data_out=16'h6;
17'h16be6:	data_out=16'h8004;
17'h16be7:	data_out=16'h3;
17'h16be8:	data_out=16'h7;
17'h16be9:	data_out=16'h8008;
17'h16bea:	data_out=16'h5;
17'h16beb:	data_out=16'h8007;
17'h16bec:	data_out=16'h8003;
17'h16bed:	data_out=16'h8009;
17'h16bee:	data_out=16'h8004;
17'h16bef:	data_out=16'h8005;
17'h16bf0:	data_out=16'h8005;
17'h16bf1:	data_out=16'h8001;
17'h16bf2:	data_out=16'h8002;
17'h16bf3:	data_out=16'h3;
17'h16bf4:	data_out=16'h8007;
17'h16bf5:	data_out=16'h8004;
17'h16bf6:	data_out=16'h8;
17'h16bf7:	data_out=16'h4;
17'h16bf8:	data_out=16'h8003;
17'h16bf9:	data_out=16'h6;
17'h16bfa:	data_out=16'h0;
17'h16bfb:	data_out=16'h2;
17'h16bfc:	data_out=16'h8002;
17'h16bfd:	data_out=16'h4;
17'h16bfe:	data_out=16'h4;
17'h16bff:	data_out=16'h8009;
17'h16c00:	data_out=16'h2;
17'h16c01:	data_out=16'h0;
17'h16c02:	data_out=16'h8005;
17'h16c03:	data_out=16'h8000;
17'h16c04:	data_out=16'h8003;
17'h16c05:	data_out=16'h8000;
17'h16c06:	data_out=16'h8006;
17'h16c07:	data_out=16'h8004;
17'h16c08:	data_out=16'h1;
17'h16c09:	data_out=16'h8;
17'h16c0a:	data_out=16'h8002;
17'h16c0b:	data_out=16'h7;
17'h16c0c:	data_out=16'h8;
17'h16c0d:	data_out=16'h3;
17'h16c0e:	data_out=16'h8007;
17'h16c0f:	data_out=16'h8007;
17'h16c10:	data_out=16'h8007;
17'h16c11:	data_out=16'h0;
17'h16c12:	data_out=16'h6;
17'h16c13:	data_out=16'h8005;
17'h16c14:	data_out=16'h5;
17'h16c15:	data_out=16'h4;
17'h16c16:	data_out=16'h8;
17'h16c17:	data_out=16'h8007;
17'h16c18:	data_out=16'h1;
17'h16c19:	data_out=16'h8001;
17'h16c1a:	data_out=16'h4;
17'h16c1b:	data_out=16'h9;
17'h16c1c:	data_out=16'h8006;
17'h16c1d:	data_out=16'h8001;
17'h16c1e:	data_out=16'h8009;
17'h16c1f:	data_out=16'h5;
17'h16c20:	data_out=16'h8;
17'h16c21:	data_out=16'h8005;
17'h16c22:	data_out=16'h8005;
17'h16c23:	data_out=16'h8004;
17'h16c24:	data_out=16'h4;
17'h16c25:	data_out=16'h8002;
17'h16c26:	data_out=16'h1;
17'h16c27:	data_out=16'h8004;
17'h16c28:	data_out=16'h8003;
17'h16c29:	data_out=16'h8;
17'h16c2a:	data_out=16'h8006;
17'h16c2b:	data_out=16'h8005;
17'h16c2c:	data_out=16'h2;
17'h16c2d:	data_out=16'h8004;
17'h16c2e:	data_out=16'h8003;
17'h16c2f:	data_out=16'h4;
17'h16c30:	data_out=16'h6;
17'h16c31:	data_out=16'h8006;
17'h16c32:	data_out=16'h8;
17'h16c33:	data_out=16'h2;
17'h16c34:	data_out=16'h7;
17'h16c35:	data_out=16'h7;
17'h16c36:	data_out=16'h4;
17'h16c37:	data_out=16'h8001;
17'h16c38:	data_out=16'h8003;
17'h16c39:	data_out=16'h8002;
17'h16c3a:	data_out=16'h8001;
17'h16c3b:	data_out=16'h0;
17'h16c3c:	data_out=16'h6;
17'h16c3d:	data_out=16'h8001;
17'h16c3e:	data_out=16'h8004;
17'h16c3f:	data_out=16'h5;
17'h16c40:	data_out=16'h3;
17'h16c41:	data_out=16'h1;
17'h16c42:	data_out=16'h8007;
17'h16c43:	data_out=16'h8002;
17'h16c44:	data_out=16'h8;
17'h16c45:	data_out=16'h3;
17'h16c46:	data_out=16'h3;
17'h16c47:	data_out=16'h8005;
17'h16c48:	data_out=16'h2;
17'h16c49:	data_out=16'h6;
17'h16c4a:	data_out=16'h8000;
17'h16c4b:	data_out=16'h8005;
17'h16c4c:	data_out=16'h8007;
17'h16c4d:	data_out=16'h6;
17'h16c4e:	data_out=16'h8;
17'h16c4f:	data_out=16'h8;
17'h16c50:	data_out=16'h8009;
17'h16c51:	data_out=16'h7;
17'h16c52:	data_out=16'h1;
17'h16c53:	data_out=16'h7;
17'h16c54:	data_out=16'h6;
17'h16c55:	data_out=16'h8004;
17'h16c56:	data_out=16'h8002;
17'h16c57:	data_out=16'h8007;
17'h16c58:	data_out=16'h3;
17'h16c59:	data_out=16'h6;
17'h16c5a:	data_out=16'h3;
17'h16c5b:	data_out=16'h0;
17'h16c5c:	data_out=16'h8004;
17'h16c5d:	data_out=16'h8;
17'h16c5e:	data_out=16'h8004;
17'h16c5f:	data_out=16'h8;
17'h16c60:	data_out=16'h8000;
17'h16c61:	data_out=16'h8002;
17'h16c62:	data_out=16'h8002;
17'h16c63:	data_out=16'h8002;
17'h16c64:	data_out=16'h8008;
17'h16c65:	data_out=16'h8009;
17'h16c66:	data_out=16'h3;
17'h16c67:	data_out=16'h4;
17'h16c68:	data_out=16'h7;
17'h16c69:	data_out=16'h8007;
17'h16c6a:	data_out=16'h8;
17'h16c6b:	data_out=16'h8009;
17'h16c6c:	data_out=16'h9;
17'h16c6d:	data_out=16'h7;
17'h16c6e:	data_out=16'h8;
17'h16c6f:	data_out=16'h9;
17'h16c70:	data_out=16'h5;
17'h16c71:	data_out=16'h0;
17'h16c72:	data_out=16'h7;
17'h16c73:	data_out=16'h2;
17'h16c74:	data_out=16'h5;
17'h16c75:	data_out=16'h8005;
17'h16c76:	data_out=16'h4;
17'h16c77:	data_out=16'h8001;
17'h16c78:	data_out=16'h8008;
17'h16c79:	data_out=16'h8002;
17'h16c7a:	data_out=16'h8;
17'h16c7b:	data_out=16'h8003;
17'h16c7c:	data_out=16'h8003;
17'h16c7d:	data_out=16'h8004;
17'h16c7e:	data_out=16'h8003;
17'h16c7f:	data_out=16'h6;
17'h16c80:	data_out=16'h3;
17'h16c81:	data_out=16'h3;
17'h16c82:	data_out=16'h8005;
17'h16c83:	data_out=16'h4;
17'h16c84:	data_out=16'h4;
17'h16c85:	data_out=16'h7;
17'h16c86:	data_out=16'h8001;
17'h16c87:	data_out=16'h1;
17'h16c88:	data_out=16'h8009;
17'h16c89:	data_out=16'h8002;
17'h16c8a:	data_out=16'h2;
17'h16c8b:	data_out=16'h9;
17'h16c8c:	data_out=16'h8005;
17'h16c8d:	data_out=16'h1;
17'h16c8e:	data_out=16'h9;
17'h16c8f:	data_out=16'h8008;
17'h16c90:	data_out=16'h8008;
17'h16c91:	data_out=16'h6;
17'h16c92:	data_out=16'h3;
17'h16c93:	data_out=16'h6;
17'h16c94:	data_out=16'h8008;
17'h16c95:	data_out=16'h8002;
17'h16c96:	data_out=16'h8004;
17'h16c97:	data_out=16'h8006;
17'h16c98:	data_out=16'h5;
17'h16c99:	data_out=16'h8005;
17'h16c9a:	data_out=16'h0;
17'h16c9b:	data_out=16'h8007;
17'h16c9c:	data_out=16'h8000;
17'h16c9d:	data_out=16'h6;
17'h16c9e:	data_out=16'h8;
17'h16c9f:	data_out=16'h8007;
17'h16ca0:	data_out=16'h8000;
17'h16ca1:	data_out=16'h8006;
17'h16ca2:	data_out=16'h7;
17'h16ca3:	data_out=16'h8005;
17'h16ca4:	data_out=16'h8009;
17'h16ca5:	data_out=16'h8003;
17'h16ca6:	data_out=16'h5;
17'h16ca7:	data_out=16'h8008;
17'h16ca8:	data_out=16'h3;
17'h16ca9:	data_out=16'h8002;
17'h16caa:	data_out=16'h8008;
17'h16cab:	data_out=16'h8;
17'h16cac:	data_out=16'h8;
17'h16cad:	data_out=16'h8009;
17'h16cae:	data_out=16'h9;
17'h16caf:	data_out=16'h9;
17'h16cb0:	data_out=16'h7;
17'h16cb1:	data_out=16'h2;
17'h16cb2:	data_out=16'h5;
17'h16cb3:	data_out=16'h8;
17'h16cb4:	data_out=16'h8009;
17'h16cb5:	data_out=16'h8008;
17'h16cb6:	data_out=16'h8007;
17'h16cb7:	data_out=16'h5;
17'h16cb8:	data_out=16'h8004;
17'h16cb9:	data_out=16'h2;
17'h16cba:	data_out=16'h7;
17'h16cbb:	data_out=16'h5;
17'h16cbc:	data_out=16'h8001;
17'h16cbd:	data_out=16'h6;
17'h16cbe:	data_out=16'h7;
17'h16cbf:	data_out=16'h8;
17'h16cc0:	data_out=16'h9;
17'h16cc1:	data_out=16'h5;
17'h16cc2:	data_out=16'h8007;
17'h16cc3:	data_out=16'h8009;
17'h16cc4:	data_out=16'h8007;
17'h16cc5:	data_out=16'h8;
17'h16cc6:	data_out=16'h8008;
17'h16cc7:	data_out=16'h5;
17'h16cc8:	data_out=16'h8004;
17'h16cc9:	data_out=16'h8007;
17'h16cca:	data_out=16'h4;
17'h16ccb:	data_out=16'h8005;
17'h16ccc:	data_out=16'h8007;
17'h16ccd:	data_out=16'h4;
17'h16cce:	data_out=16'h8006;
17'h16ccf:	data_out=16'h8009;
17'h16cd0:	data_out=16'h8003;
17'h16cd1:	data_out=16'h9;
17'h16cd2:	data_out=16'h8;
17'h16cd3:	data_out=16'h8003;
17'h16cd4:	data_out=16'h8008;
17'h16cd5:	data_out=16'h8008;
17'h16cd6:	data_out=16'h8006;
17'h16cd7:	data_out=16'h8003;
17'h16cd8:	data_out=16'h3;
17'h16cd9:	data_out=16'h8008;
17'h16cda:	data_out=16'h8008;
17'h16cdb:	data_out=16'h8007;
17'h16cdc:	data_out=16'h7;
17'h16cdd:	data_out=16'h9;
17'h16cde:	data_out=16'h8008;
17'h16cdf:	data_out=16'h7;
17'h16ce0:	data_out=16'h5;
17'h16ce1:	data_out=16'h8006;
17'h16ce2:	data_out=16'h7;
17'h16ce3:	data_out=16'h7;
17'h16ce4:	data_out=16'h8007;
17'h16ce5:	data_out=16'h8;
17'h16ce6:	data_out=16'h3;
17'h16ce7:	data_out=16'h8002;
17'h16ce8:	data_out=16'h8008;
17'h16ce9:	data_out=16'h8002;
17'h16cea:	data_out=16'h2;
17'h16ceb:	data_out=16'h8005;
17'h16cec:	data_out=16'h8007;
17'h16ced:	data_out=16'h5;
17'h16cee:	data_out=16'h8005;
17'h16cef:	data_out=16'h8001;
17'h16cf0:	data_out=16'h5;
17'h16cf1:	data_out=16'h8006;
17'h16cf2:	data_out=16'h6;
17'h16cf3:	data_out=16'h6;
17'h16cf4:	data_out=16'h8005;
17'h16cf5:	data_out=16'h8;
17'h16cf6:	data_out=16'h8007;
17'h16cf7:	data_out=16'h7;
17'h16cf8:	data_out=16'h8009;
17'h16cf9:	data_out=16'h8006;
17'h16cfa:	data_out=16'h9;
17'h16cfb:	data_out=16'h7;
17'h16cfc:	data_out=16'h8006;
17'h16cfd:	data_out=16'h8009;
17'h16cfe:	data_out=16'h5;
17'h16cff:	data_out=16'h8;
17'h16d00:	data_out=16'h8006;
17'h16d01:	data_out=16'h3;
17'h16d02:	data_out=16'h5;
17'h16d03:	data_out=16'h8004;
17'h16d04:	data_out=16'h2;
17'h16d05:	data_out=16'h8001;
17'h16d06:	data_out=16'h3;
17'h16d07:	data_out=16'h3;
17'h16d08:	data_out=16'h6;
17'h16d09:	data_out=16'h8004;
17'h16d0a:	data_out=16'h7;
17'h16d0b:	data_out=16'h8;
17'h16d0c:	data_out=16'h8008;
17'h16d0d:	data_out=16'h8008;
17'h16d0e:	data_out=16'h8002;
17'h16d0f:	data_out=16'h5;
17'h16d10:	data_out=16'h8005;
17'h16d11:	data_out=16'h8006;
17'h16d12:	data_out=16'h2;
17'h16d13:	data_out=16'h8001;
17'h16d14:	data_out=16'h8006;
17'h16d15:	data_out=16'h4;
17'h16d16:	data_out=16'h8004;
17'h16d17:	data_out=16'h8006;
17'h16d18:	data_out=16'h8;
17'h16d19:	data_out=16'h8004;
17'h16d1a:	data_out=16'h8008;
17'h16d1b:	data_out=16'h8008;
17'h16d1c:	data_out=16'h8004;
17'h16d1d:	data_out=16'h6;
17'h16d1e:	data_out=16'h8009;
17'h16d1f:	data_out=16'h8000;
17'h16d20:	data_out=16'h8000;
17'h16d21:	data_out=16'h5;
17'h16d22:	data_out=16'h5;
17'h16d23:	data_out=16'h8008;
17'h16d24:	data_out=16'h8005;
17'h16d25:	data_out=16'h8001;
17'h16d26:	data_out=16'h4;
17'h16d27:	data_out=16'h8008;
17'h16d28:	data_out=16'h3;
17'h16d29:	data_out=16'h2;
17'h16d2a:	data_out=16'h9;
17'h16d2b:	data_out=16'h4;
17'h16d2c:	data_out=16'h3;
17'h16d2d:	data_out=16'h8003;
17'h16d2e:	data_out=16'h0;
17'h16d2f:	data_out=16'h7;
17'h16d30:	data_out=16'h1;
17'h16d31:	data_out=16'h8007;
17'h16d32:	data_out=16'h8004;
17'h16d33:	data_out=16'h4;
17'h16d34:	data_out=16'h6;
17'h16d35:	data_out=16'h2;
17'h16d36:	data_out=16'h7;
17'h16d37:	data_out=16'h4;
17'h16d38:	data_out=16'h7;
17'h16d39:	data_out=16'h8;
17'h16d3a:	data_out=16'h6;
17'h16d3b:	data_out=16'h8006;
17'h16d3c:	data_out=16'h6;
17'h16d3d:	data_out=16'h6;
17'h16d3e:	data_out=16'h3;
17'h16d3f:	data_out=16'h8004;
17'h16d40:	data_out=16'h2;
17'h16d41:	data_out=16'h8002;
17'h16d42:	data_out=16'h8002;
17'h16d43:	data_out=16'h7;
17'h16d44:	data_out=16'h6;
17'h16d45:	data_out=16'h8007;
17'h16d46:	data_out=16'h7;
17'h16d47:	data_out=16'h0;
17'h16d48:	data_out=16'h4;
17'h16d49:	data_out=16'h7;
17'h16d4a:	data_out=16'h8005;
17'h16d4b:	data_out=16'h8002;
17'h16d4c:	data_out=16'h8005;
17'h16d4d:	data_out=16'h4;
17'h16d4e:	data_out=16'h8005;
17'h16d4f:	data_out=16'h5;
17'h16d50:	data_out=16'h6;
17'h16d51:	data_out=16'h1;
17'h16d52:	data_out=16'h8000;
17'h16d53:	data_out=16'h3;
17'h16d54:	data_out=16'h8006;
17'h16d55:	data_out=16'h8002;
17'h16d56:	data_out=16'h8002;
17'h16d57:	data_out=16'h8009;
17'h16d58:	data_out=16'h8003;
17'h16d59:	data_out=16'h8005;
17'h16d5a:	data_out=16'h8005;
17'h16d5b:	data_out=16'h8007;
17'h16d5c:	data_out=16'h8008;
17'h16d5d:	data_out=16'h6;
17'h16d5e:	data_out=16'h8001;
17'h16d5f:	data_out=16'h4;
17'h16d60:	data_out=16'h8004;
17'h16d61:	data_out=16'h6;
17'h16d62:	data_out=16'h1;
17'h16d63:	data_out=16'h8007;
17'h16d64:	data_out=16'h8;
17'h16d65:	data_out=16'h8001;
17'h16d66:	data_out=16'h2;
17'h16d67:	data_out=16'h3;
17'h16d68:	data_out=16'h8003;
17'h16d69:	data_out=16'h6;
17'h16d6a:	data_out=16'h8008;
17'h16d6b:	data_out=16'h2;
17'h16d6c:	data_out=16'h1;
17'h16d6d:	data_out=16'h8004;
17'h16d6e:	data_out=16'h8002;
17'h16d6f:	data_out=16'h8002;
17'h16d70:	data_out=16'h6;
17'h16d71:	data_out=16'h7;
17'h16d72:	data_out=16'h8008;
17'h16d73:	data_out=16'h9;
17'h16d74:	data_out=16'h8004;
17'h16d75:	data_out=16'h8001;
17'h16d76:	data_out=16'h8009;
17'h16d77:	data_out=16'h2;
17'h16d78:	data_out=16'h3;
17'h16d79:	data_out=16'h8005;
17'h16d7a:	data_out=16'h4;
17'h16d7b:	data_out=16'h5;
17'h16d7c:	data_out=16'h8008;
17'h16d7d:	data_out=16'h8006;
17'h16d7e:	data_out=16'h8001;
17'h16d7f:	data_out=16'h8003;
17'h16d80:	data_out=16'h802d;
17'h16d81:	data_out=16'h8041;
17'h16d82:	data_out=16'h10;
17'h16d83:	data_out=16'h8021;
17'h16d84:	data_out=16'h8046;
17'h16d85:	data_out=16'h8045;
17'h16d86:	data_out=16'h800a;
17'h16d87:	data_out=16'h8017;
17'h16d88:	data_out=16'h800e;
17'h16d89:	data_out=16'h10;
17'h16d8a:	data_out=16'h802f;
17'h16d8b:	data_out=16'h6;
17'h16d8c:	data_out=16'h8040;
17'h16d8d:	data_out=16'h8027;
17'h16d8e:	data_out=16'h8001;
17'h16d8f:	data_out=16'h8004;
17'h16d90:	data_out=16'h18;
17'h16d91:	data_out=16'h8036;
17'h16d92:	data_out=16'h5;
17'h16d93:	data_out=16'h800d;
17'h16d94:	data_out=16'h8010;
17'h16d95:	data_out=16'h801a;
17'h16d96:	data_out=16'h802b;
17'h16d97:	data_out=16'h8009;
17'h16d98:	data_out=16'h800e;
17'h16d99:	data_out=16'h8034;
17'h16d9a:	data_out=16'h8048;
17'h16d9b:	data_out=16'h8025;
17'h16d9c:	data_out=16'h804c;
17'h16d9d:	data_out=16'h8030;
17'h16d9e:	data_out=16'h801a;
17'h16d9f:	data_out=16'h8018;
17'h16da0:	data_out=16'h805a;
17'h16da1:	data_out=16'h2;
17'h16da2:	data_out=16'ha;
17'h16da3:	data_out=16'h8030;
17'h16da4:	data_out=16'h8029;
17'h16da5:	data_out=16'h801a;
17'h16da6:	data_out=16'h1c;
17'h16da7:	data_out=16'h8029;
17'h16da8:	data_out=16'h8002;
17'h16da9:	data_out=16'h8007;
17'h16daa:	data_out=16'hd;
17'h16dab:	data_out=16'h8023;
17'h16dac:	data_out=16'h8020;
17'h16dad:	data_out=16'h8003;
17'h16dae:	data_out=16'h2c;
17'h16daf:	data_out=16'h8026;
17'h16db0:	data_out=16'h8050;
17'h16db1:	data_out=16'h804f;
17'h16db2:	data_out=16'h805b;
17'h16db3:	data_out=16'h801b;
17'h16db4:	data_out=16'h8038;
17'h16db5:	data_out=16'h8043;
17'h16db6:	data_out=16'h801a;
17'h16db7:	data_out=16'h8004;
17'h16db8:	data_out=16'h8063;
17'h16db9:	data_out=16'h0;
17'h16dba:	data_out=16'h1;
17'h16dbb:	data_out=16'h8037;
17'h16dbc:	data_out=16'h3;
17'h16dbd:	data_out=16'h8031;
17'h16dbe:	data_out=16'h800b;
17'h16dbf:	data_out=16'h8035;
17'h16dc0:	data_out=16'h800d;
17'h16dc1:	data_out=16'h3;
17'h16dc2:	data_out=16'h8024;
17'h16dc3:	data_out=16'h13;
17'h16dc4:	data_out=16'h8017;
17'h16dc5:	data_out=16'h8015;
17'h16dc6:	data_out=16'h8005;
17'h16dc7:	data_out=16'h8021;
17'h16dc8:	data_out=16'h2b;
17'h16dc9:	data_out=16'h800d;
17'h16dca:	data_out=16'h8033;
17'h16dcb:	data_out=16'h805a;
17'h16dcc:	data_out=16'h8033;
17'h16dcd:	data_out=16'h8009;
17'h16dce:	data_out=16'h802e;
17'h16dcf:	data_out=16'h803a;
17'h16dd0:	data_out=16'h801a;
17'h16dd1:	data_out=16'h8018;
17'h16dd2:	data_out=16'h802c;
17'h16dd3:	data_out=16'h804e;
17'h16dd4:	data_out=16'h802b;
17'h16dd5:	data_out=16'h2e;
17'h16dd6:	data_out=16'h4;
17'h16dd7:	data_out=16'h2e;
17'h16dd8:	data_out=16'h26;
17'h16dd9:	data_out=16'h32;
17'h16dda:	data_out=16'h2a;
17'h16ddb:	data_out=16'h8058;
17'h16ddc:	data_out=16'h8031;
17'h16ddd:	data_out=16'h801b;
17'h16dde:	data_out=16'h8020;
17'h16ddf:	data_out=16'h8010;
17'h16de0:	data_out=16'h1;
17'h16de1:	data_out=16'h804d;
17'h16de2:	data_out=16'h8017;
17'h16de3:	data_out=16'h8016;
17'h16de4:	data_out=16'h8028;
17'h16de5:	data_out=16'h800a;
17'h16de6:	data_out=16'h8021;
17'h16de7:	data_out=16'h20;
17'h16de8:	data_out=16'h8007;
17'h16de9:	data_out=16'h0;
17'h16dea:	data_out=16'h8006;
17'h16deb:	data_out=16'h8053;
17'h16dec:	data_out=16'h8023;
17'h16ded:	data_out=16'h801e;
17'h16dee:	data_out=16'h8005;
17'h16def:	data_out=16'h802d;
17'h16df0:	data_out=16'h800f;
17'h16df1:	data_out=16'hf;
17'h16df2:	data_out=16'h8010;
17'h16df3:	data_out=16'h802f;
17'h16df4:	data_out=16'h805f;
17'h16df5:	data_out=16'h8020;
17'h16df6:	data_out=16'h801f;
17'h16df7:	data_out=16'h4;
17'h16df8:	data_out=16'h8017;
17'h16df9:	data_out=16'h13;
17'h16dfa:	data_out=16'h8010;
17'h16dfb:	data_out=16'h8007;
17'h16dfc:	data_out=16'h800a;
17'h16dfd:	data_out=16'h801d;
17'h16dfe:	data_out=16'h14;
17'h16dff:	data_out=16'h8020;
17'h16e00:	data_out=16'h837d;
17'h16e01:	data_out=16'h84cb;
17'h16e02:	data_out=16'hf0;
17'h16e03:	data_out=16'h82dd;
17'h16e04:	data_out=16'h88c8;
17'h16e05:	data_out=16'h86f8;
17'h16e06:	data_out=16'h803f;
17'h16e07:	data_out=16'h83e1;
17'h16e08:	data_out=16'h51;
17'h16e09:	data_out=16'h424;
17'h16e0a:	data_out=16'h8546;
17'h16e0b:	data_out=16'h47b;
17'h16e0c:	data_out=16'h87bd;
17'h16e0d:	data_out=16'h81e0;
17'h16e0e:	data_out=16'h80d5;
17'h16e0f:	data_out=16'h8048;
17'h16e10:	data_out=16'h372;
17'h16e11:	data_out=16'h883a;
17'h16e12:	data_out=16'h214;
17'h16e13:	data_out=16'h8193;
17'h16e14:	data_out=16'h1cc;
17'h16e15:	data_out=16'h829f;
17'h16e16:	data_out=16'h83d4;
17'h16e17:	data_out=16'h17b;
17'h16e18:	data_out=16'h8097;
17'h16e19:	data_out=16'h8436;
17'h16e1a:	data_out=16'h88c9;
17'h16e1b:	data_out=16'h26;
17'h16e1c:	data_out=16'h8811;
17'h16e1d:	data_out=16'h851d;
17'h16e1e:	data_out=16'hba;
17'h16e1f:	data_out=16'h8266;
17'h16e20:	data_out=16'h8664;
17'h16e21:	data_out=16'h80bc;
17'h16e22:	data_out=16'h3e1;
17'h16e23:	data_out=16'h81af;
17'h16e24:	data_out=16'h81af;
17'h16e25:	data_out=16'hab;
17'h16e26:	data_out=16'h461;
17'h16e27:	data_out=16'h8525;
17'h16e28:	data_out=16'h80a8;
17'h16e29:	data_out=16'hff;
17'h16e2a:	data_out=16'h23f;
17'h16e2b:	data_out=16'h81a6;
17'h16e2c:	data_out=16'h83ab;
17'h16e2d:	data_out=16'h406;
17'h16e2e:	data_out=16'h265;
17'h16e2f:	data_out=16'h819a;
17'h16e30:	data_out=16'h8949;
17'h16e31:	data_out=16'h8684;
17'h16e32:	data_out=16'h8969;
17'h16e33:	data_out=16'h156;
17'h16e34:	data_out=16'h865d;
17'h16e35:	data_out=16'h8823;
17'h16e36:	data_out=16'hb6;
17'h16e37:	data_out=16'h116;
17'h16e38:	data_out=16'h88c4;
17'h16e39:	data_out=16'haf;
17'h16e3a:	data_out=16'h11;
17'h16e3b:	data_out=16'h85e6;
17'h16e3c:	data_out=16'h101;
17'h16e3d:	data_out=16'h8503;
17'h16e3e:	data_out=16'h80b1;
17'h16e3f:	data_out=16'h86fb;
17'h16e40:	data_out=16'h8026;
17'h16e41:	data_out=16'h217;
17'h16e42:	data_out=16'h27;
17'h16e43:	data_out=16'h225;
17'h16e44:	data_out=16'h84a3;
17'h16e45:	data_out=16'h82ad;
17'h16e46:	data_out=16'h423;
17'h16e47:	data_out=16'h8085;
17'h16e48:	data_out=16'h318;
17'h16e49:	data_out=16'hdd;
17'h16e4a:	data_out=16'h8675;
17'h16e4b:	data_out=16'h84f3;
17'h16e4c:	data_out=16'h82c1;
17'h16e4d:	data_out=16'h293;
17'h16e4e:	data_out=16'h817a;
17'h16e4f:	data_out=16'h82f2;
17'h16e50:	data_out=16'h80bc;
17'h16e51:	data_out=16'h835c;
17'h16e52:	data_out=16'h81cf;
17'h16e53:	data_out=16'h8544;
17'h16e54:	data_out=16'h82ee;
17'h16e55:	data_out=16'h4ae;
17'h16e56:	data_out=16'h1d3;
17'h16e57:	data_out=16'h29c;
17'h16e58:	data_out=16'h2a8;
17'h16e59:	data_out=16'h37;
17'h16e5a:	data_out=16'h1c0;
17'h16e5b:	data_out=16'h8a00;
17'h16e5c:	data_out=16'h8649;
17'h16e5d:	data_out=16'h82cf;
17'h16e5e:	data_out=16'h8107;
17'h16e5f:	data_out=16'h8124;
17'h16e60:	data_out=16'h8e;
17'h16e61:	data_out=16'h892c;
17'h16e62:	data_out=16'ha3;
17'h16e63:	data_out=16'h151;
17'h16e64:	data_out=16'h83c9;
17'h16e65:	data_out=16'h830d;
17'h16e66:	data_out=16'h825f;
17'h16e67:	data_out=16'h315;
17'h16e68:	data_out=16'h80be;
17'h16e69:	data_out=16'h13b;
17'h16e6a:	data_out=16'h80df;
17'h16e6b:	data_out=16'h889d;
17'h16e6c:	data_out=16'h848e;
17'h16e6d:	data_out=16'h137;
17'h16e6e:	data_out=16'h80dd;
17'h16e6f:	data_out=16'h83fb;
17'h16e70:	data_out=16'h80d0;
17'h16e71:	data_out=16'h81b1;
17'h16e72:	data_out=16'h8815;
17'h16e73:	data_out=16'h8801;
17'h16e74:	data_out=16'h894f;
17'h16e75:	data_out=16'h8338;
17'h16e76:	data_out=16'h8046;
17'h16e77:	data_out=16'h181;
17'h16e78:	data_out=16'h8021;
17'h16e79:	data_out=16'h71;
17'h16e7a:	data_out=16'h1e0;
17'h16e7b:	data_out=16'h80a3;
17'h16e7c:	data_out=16'h80df;
17'h16e7d:	data_out=16'h8032;
17'h16e7e:	data_out=16'h56c;
17'h16e7f:	data_out=16'h84b4;
17'h16e80:	data_out=16'h8752;
17'h16e81:	data_out=16'h8620;
17'h16e82:	data_out=16'h31d;
17'h16e83:	data_out=16'h816b;
17'h16e84:	data_out=16'h8a00;
17'h16e85:	data_out=16'h8a00;
17'h16e86:	data_out=16'h187;
17'h16e87:	data_out=16'h842e;
17'h16e88:	data_out=16'h215;
17'h16e89:	data_out=16'h7f1;
17'h16e8a:	data_out=16'h89ea;
17'h16e8b:	data_out=16'h889;
17'h16e8c:	data_out=16'h89fe;
17'h16e8d:	data_out=16'h804b;
17'h16e8e:	data_out=16'h80a2;
17'h16e8f:	data_out=16'h356;
17'h16e90:	data_out=16'h742;
17'h16e91:	data_out=16'h8a00;
17'h16e92:	data_out=16'h609;
17'h16e93:	data_out=16'h8063;
17'h16e94:	data_out=16'h517;
17'h16e95:	data_out=16'h8438;
17'h16e96:	data_out=16'h862a;
17'h16e97:	data_out=16'h51c;
17'h16e98:	data_out=16'h42;
17'h16e99:	data_out=16'h882c;
17'h16e9a:	data_out=16'h8a00;
17'h16e9b:	data_out=16'h4b0;
17'h16e9c:	data_out=16'h8971;
17'h16e9d:	data_out=16'h8785;
17'h16e9e:	data_out=16'h2eb;
17'h16e9f:	data_out=16'h81ba;
17'h16ea0:	data_out=16'h8810;
17'h16ea1:	data_out=16'h807a;
17'h16ea2:	data_out=16'h854;
17'h16ea3:	data_out=16'h825b;
17'h16ea4:	data_out=16'h825c;
17'h16ea5:	data_out=16'h375;
17'h16ea6:	data_out=16'h6a0;
17'h16ea7:	data_out=16'h8723;
17'h16ea8:	data_out=16'h803a;
17'h16ea9:	data_out=16'h406;
17'h16eaa:	data_out=16'h4ef;
17'h16eab:	data_out=16'h8076;
17'h16eac:	data_out=16'h8601;
17'h16ead:	data_out=16'h75f;
17'h16eae:	data_out=16'h53f;
17'h16eaf:	data_out=16'h9;
17'h16eb0:	data_out=16'h89ff;
17'h16eb1:	data_out=16'h8a00;
17'h16eb2:	data_out=16'h8a00;
17'h16eb3:	data_out=16'h4fa;
17'h16eb4:	data_out=16'h8a00;
17'h16eb5:	data_out=16'h89ff;
17'h16eb6:	data_out=16'h381;
17'h16eb7:	data_out=16'h373;
17'h16eb8:	data_out=16'h8a00;
17'h16eb9:	data_out=16'h44f;
17'h16eba:	data_out=16'h1ce;
17'h16ebb:	data_out=16'h8a00;
17'h16ebc:	data_out=16'h2a7;
17'h16ebd:	data_out=16'h8895;
17'h16ebe:	data_out=16'h8040;
17'h16ebf:	data_out=16'h8a00;
17'h16ec0:	data_out=16'h80fb;
17'h16ec1:	data_out=16'h443;
17'h16ec2:	data_out=16'h291;
17'h16ec3:	data_out=16'h3fb;
17'h16ec4:	data_out=16'h88d6;
17'h16ec5:	data_out=16'h8450;
17'h16ec6:	data_out=16'h84b;
17'h16ec7:	data_out=16'h267;
17'h16ec8:	data_out=16'h6c8;
17'h16ec9:	data_out=16'h35f;
17'h16eca:	data_out=16'h889a;
17'h16ecb:	data_out=16'h85f7;
17'h16ecc:	data_out=16'h8128;
17'h16ecd:	data_out=16'h7d3;
17'h16ece:	data_out=16'h82;
17'h16ecf:	data_out=16'h8263;
17'h16ed0:	data_out=16'h8002;
17'h16ed1:	data_out=16'h8369;
17'h16ed2:	data_out=16'h8301;
17'h16ed3:	data_out=16'h83f9;
17'h16ed4:	data_out=16'h8272;
17'h16ed5:	data_out=16'h892;
17'h16ed6:	data_out=16'h4bd;
17'h16ed7:	data_out=16'h5fe;
17'h16ed8:	data_out=16'h567;
17'h16ed9:	data_out=16'h80d9;
17'h16eda:	data_out=16'h62b;
17'h16edb:	data_out=16'h8a00;
17'h16edc:	data_out=16'h87ad;
17'h16edd:	data_out=16'h849e;
17'h16ede:	data_out=16'hf9;
17'h16edf:	data_out=16'h80a3;
17'h16ee0:	data_out=16'h125;
17'h16ee1:	data_out=16'h8a00;
17'h16ee2:	data_out=16'h300;
17'h16ee3:	data_out=16'h4ee;
17'h16ee4:	data_out=16'h852c;
17'h16ee5:	data_out=16'h8472;
17'h16ee6:	data_out=16'h846a;
17'h16ee7:	data_out=16'h7d7;
17'h16ee8:	data_out=16'h8066;
17'h16ee9:	data_out=16'h43a;
17'h16eea:	data_out=16'h80c7;
17'h16eeb:	data_out=16'h89ff;
17'h16eec:	data_out=16'h89e3;
17'h16eed:	data_out=16'h4cf;
17'h16eee:	data_out=16'h80c2;
17'h16eef:	data_out=16'h86fe;
17'h16ef0:	data_out=16'h8099;
17'h16ef1:	data_out=16'h81e5;
17'h16ef2:	data_out=16'h8a00;
17'h16ef3:	data_out=16'h8a00;
17'h16ef4:	data_out=16'h89ff;
17'h16ef5:	data_out=16'h841b;
17'h16ef6:	data_out=16'h29;
17'h16ef7:	data_out=16'h4a6;
17'h16ef8:	data_out=16'hd5;
17'h16ef9:	data_out=16'h299;
17'h16efa:	data_out=16'h4ff;
17'h16efb:	data_out=16'h802e;
17'h16efc:	data_out=16'h809b;
17'h16efd:	data_out=16'h176;
17'h16efe:	data_out=16'ha00;
17'h16eff:	data_out=16'h8727;
17'h16f00:	data_out=16'h876c;
17'h16f01:	data_out=16'h83e2;
17'h16f02:	data_out=16'ha00;
17'h16f03:	data_out=16'h81f;
17'h16f04:	data_out=16'h890a;
17'h16f05:	data_out=16'h81de;
17'h16f06:	data_out=16'h732;
17'h16f07:	data_out=16'he1;
17'h16f08:	data_out=16'h96d;
17'h16f09:	data_out=16'ha00;
17'h16f0a:	data_out=16'h86a5;
17'h16f0b:	data_out=16'ha00;
17'h16f0c:	data_out=16'h85aa;
17'h16f0d:	data_out=16'h5fa;
17'h16f0e:	data_out=16'h195;
17'h16f0f:	data_out=16'h969;
17'h16f10:	data_out=16'ha00;
17'h16f11:	data_out=16'h85e7;
17'h16f12:	data_out=16'h9e6;
17'h16f13:	data_out=16'h938;
17'h16f14:	data_out=16'ha00;
17'h16f15:	data_out=16'h813d;
17'h16f16:	data_out=16'h94;
17'h16f17:	data_out=16'ha00;
17'h16f18:	data_out=16'hc5;
17'h16f19:	data_out=16'h8747;
17'h16f1a:	data_out=16'h8822;
17'h16f1b:	data_out=16'ha00;
17'h16f1c:	data_out=16'h827b;
17'h16f1d:	data_out=16'h80df;
17'h16f1e:	data_out=16'h972;
17'h16f1f:	data_out=16'h2d9;
17'h16f20:	data_out=16'h8294;
17'h16f21:	data_out=16'h1ac;
17'h16f22:	data_out=16'ha00;
17'h16f23:	data_out=16'h81d4;
17'h16f24:	data_out=16'h81d3;
17'h16f25:	data_out=16'ha00;
17'h16f26:	data_out=16'ha00;
17'h16f27:	data_out=16'h802f;
17'h16f28:	data_out=16'h1e4;
17'h16f29:	data_out=16'ha00;
17'h16f2a:	data_out=16'h884;
17'h16f2b:	data_out=16'h4f3;
17'h16f2c:	data_out=16'h800f;
17'h16f2d:	data_out=16'h9b9;
17'h16f2e:	data_out=16'h9cc;
17'h16f2f:	data_out=16'h8f6;
17'h16f30:	data_out=16'h88f7;
17'h16f31:	data_out=16'h8796;
17'h16f32:	data_out=16'h8907;
17'h16f33:	data_out=16'ha00;
17'h16f34:	data_out=16'h8941;
17'h16f35:	data_out=16'h82ae;
17'h16f36:	data_out=16'h948;
17'h16f37:	data_out=16'ha00;
17'h16f38:	data_out=16'h887c;
17'h16f39:	data_out=16'ha00;
17'h16f3a:	data_out=16'h49e;
17'h16f3b:	data_out=16'h86d1;
17'h16f3c:	data_out=16'ha00;
17'h16f3d:	data_out=16'h8226;
17'h16f3e:	data_out=16'h1e7;
17'h16f3f:	data_out=16'h81f7;
17'h16f40:	data_out=16'h832;
17'h16f41:	data_out=16'ha00;
17'h16f42:	data_out=16'h692;
17'h16f43:	data_out=16'ha00;
17'h16f44:	data_out=16'h82d3;
17'h16f45:	data_out=16'h81ee;
17'h16f46:	data_out=16'ha00;
17'h16f47:	data_out=16'h786;
17'h16f48:	data_out=16'h9cc;
17'h16f49:	data_out=16'ha00;
17'h16f4a:	data_out=16'h82f6;
17'h16f4b:	data_out=16'h816f;
17'h16f4c:	data_out=16'h3a7;
17'h16f4d:	data_out=16'ha00;
17'h16f4e:	data_out=16'h99e;
17'h16f4f:	data_out=16'h2f5;
17'h16f50:	data_out=16'h851;
17'h16f51:	data_out=16'h407;
17'h16f52:	data_out=16'h8277;
17'h16f53:	data_out=16'h361;
17'h16f54:	data_out=16'h413;
17'h16f55:	data_out=16'ha00;
17'h16f56:	data_out=16'ha00;
17'h16f57:	data_out=16'h9ff;
17'h16f58:	data_out=16'ha00;
17'h16f59:	data_out=16'h6db;
17'h16f5a:	data_out=16'ha00;
17'h16f5b:	data_out=16'h89ff;
17'h16f5c:	data_out=16'h8008;
17'h16f5d:	data_out=16'h134;
17'h16f5e:	data_out=16'h92f;
17'h16f5f:	data_out=16'h8028;
17'h16f60:	data_out=16'h714;
17'h16f61:	data_out=16'h893e;
17'h16f62:	data_out=16'h9dd;
17'h16f63:	data_out=16'ha00;
17'h16f64:	data_out=16'ha0;
17'h16f65:	data_out=16'h61b;
17'h16f66:	data_out=16'h22;
17'h16f67:	data_out=16'h98c;
17'h16f68:	data_out=16'h1c1;
17'h16f69:	data_out=16'ha00;
17'h16f6a:	data_out=16'h189;
17'h16f6b:	data_out=16'h868c;
17'h16f6c:	data_out=16'h8a00;
17'h16f6d:	data_out=16'ha00;
17'h16f6e:	data_out=16'h189;
17'h16f6f:	data_out=16'h46a;
17'h16f70:	data_out=16'h18f;
17'h16f71:	data_out=16'h80f0;
17'h16f72:	data_out=16'h885f;
17'h16f73:	data_out=16'h8354;
17'h16f74:	data_out=16'h8913;
17'h16f75:	data_out=16'h797;
17'h16f76:	data_out=16'h64f;
17'h16f77:	data_out=16'ha00;
17'h16f78:	data_out=16'h834;
17'h16f79:	data_out=16'h9f3;
17'h16f7a:	data_out=16'ha00;
17'h16f7b:	data_out=16'h1e7;
17'h16f7c:	data_out=16'h8114;
17'h16f7d:	data_out=16'h67a;
17'h16f7e:	data_out=16'ha00;
17'h16f7f:	data_out=16'h828b;
17'h16f80:	data_out=16'h293;
17'h16f81:	data_out=16'h742;
17'h16f82:	data_out=16'ha00;
17'h16f83:	data_out=16'ha00;
17'h16f84:	data_out=16'h875;
17'h16f85:	data_out=16'h9e9;
17'h16f86:	data_out=16'ha00;
17'h16f87:	data_out=16'h8fc;
17'h16f88:	data_out=16'h9ff;
17'h16f89:	data_out=16'ha00;
17'h16f8a:	data_out=16'h885;
17'h16f8b:	data_out=16'ha00;
17'h16f8c:	data_out=16'ha00;
17'h16f8d:	data_out=16'ha00;
17'h16f8e:	data_out=16'h293;
17'h16f8f:	data_out=16'h9d7;
17'h16f90:	data_out=16'ha00;
17'h16f91:	data_out=16'ha00;
17'h16f92:	data_out=16'h9aa;
17'h16f93:	data_out=16'h9fb;
17'h16f94:	data_out=16'ha00;
17'h16f95:	data_out=16'h47e;
17'h16f96:	data_out=16'h9ff;
17'h16f97:	data_out=16'ha00;
17'h16f98:	data_out=16'h112;
17'h16f99:	data_out=16'h43c;
17'h16f9a:	data_out=16'h9c2;
17'h16f9b:	data_out=16'ha00;
17'h16f9c:	data_out=16'ha00;
17'h16f9d:	data_out=16'h816;
17'h16f9e:	data_out=16'ha00;
17'h16f9f:	data_out=16'h7fd;
17'h16fa0:	data_out=16'h85d;
17'h16fa1:	data_out=16'h2af;
17'h16fa2:	data_out=16'ha00;
17'h16fa3:	data_out=16'h80d7;
17'h16fa4:	data_out=16'h80d5;
17'h16fa5:	data_out=16'ha00;
17'h16fa6:	data_out=16'ha00;
17'h16fa7:	data_out=16'h8e0;
17'h16fa8:	data_out=16'h30d;
17'h16fa9:	data_out=16'ha00;
17'h16faa:	data_out=16'h8c0;
17'h16fab:	data_out=16'h9fe;
17'h16fac:	data_out=16'h9f2;
17'h16fad:	data_out=16'h9b9;
17'h16fae:	data_out=16'ha00;
17'h16faf:	data_out=16'h989;
17'h16fb0:	data_out=16'h9ff;
17'h16fb1:	data_out=16'h92b;
17'h16fb2:	data_out=16'h9ff;
17'h16fb3:	data_out=16'ha00;
17'h16fb4:	data_out=16'h81b0;
17'h16fb5:	data_out=16'h9b1;
17'h16fb6:	data_out=16'h9ab;
17'h16fb7:	data_out=16'ha00;
17'h16fb8:	data_out=16'h9f1;
17'h16fb9:	data_out=16'ha00;
17'h16fba:	data_out=16'h9fc;
17'h16fbb:	data_out=16'h930;
17'h16fbc:	data_out=16'ha00;
17'h16fbd:	data_out=16'h8da;
17'h16fbe:	data_out=16'h311;
17'h16fbf:	data_out=16'h9e1;
17'h16fc0:	data_out=16'h9ef;
17'h16fc1:	data_out=16'ha00;
17'h16fc2:	data_out=16'ha00;
17'h16fc3:	data_out=16'ha00;
17'h16fc4:	data_out=16'h996;
17'h16fc5:	data_out=16'h4ec;
17'h16fc6:	data_out=16'ha00;
17'h16fc7:	data_out=16'h8b7;
17'h16fc8:	data_out=16'h9f8;
17'h16fc9:	data_out=16'ha00;
17'h16fca:	data_out=16'h849;
17'h16fcb:	data_out=16'h9bc;
17'h16fcc:	data_out=16'h9fb;
17'h16fcd:	data_out=16'ha00;
17'h16fce:	data_out=16'h9db;
17'h16fcf:	data_out=16'h9e0;
17'h16fd0:	data_out=16'ha00;
17'h16fd1:	data_out=16'ha00;
17'h16fd2:	data_out=16'h811c;
17'h16fd3:	data_out=16'h927;
17'h16fd4:	data_out=16'h7d6;
17'h16fd5:	data_out=16'ha00;
17'h16fd6:	data_out=16'ha00;
17'h16fd7:	data_out=16'h9fe;
17'h16fd8:	data_out=16'ha00;
17'h16fd9:	data_out=16'h943;
17'h16fda:	data_out=16'ha00;
17'h16fdb:	data_out=16'h914;
17'h16fdc:	data_out=16'ha00;
17'h16fdd:	data_out=16'h8c6;
17'h16fde:	data_out=16'h9f6;
17'h16fdf:	data_out=16'h49f;
17'h16fe0:	data_out=16'ha00;
17'h16fe1:	data_out=16'h9e2;
17'h16fe2:	data_out=16'ha00;
17'h16fe3:	data_out=16'ha00;
17'h16fe4:	data_out=16'h92a;
17'h16fe5:	data_out=16'h9f9;
17'h16fe6:	data_out=16'h8bd;
17'h16fe7:	data_out=16'h9e4;
17'h16fe8:	data_out=16'h2cb;
17'h16fe9:	data_out=16'ha00;
17'h16fea:	data_out=16'h280;
17'h16feb:	data_out=16'h9fe;
17'h16fec:	data_out=16'h8235;
17'h16fed:	data_out=16'ha00;
17'h16fee:	data_out=16'h280;
17'h16fef:	data_out=16'ha00;
17'h16ff0:	data_out=16'h28b;
17'h16ff1:	data_out=16'h4a8;
17'h16ff2:	data_out=16'h962;
17'h16ff3:	data_out=16'h9ba;
17'h16ff4:	data_out=16'h9ff;
17'h16ff5:	data_out=16'ha00;
17'h16ff6:	data_out=16'ha00;
17'h16ff7:	data_out=16'ha00;
17'h16ff8:	data_out=16'ha00;
17'h16ff9:	data_out=16'h9d7;
17'h16ffa:	data_out=16'ha00;
17'h16ffb:	data_out=16'h313;
17'h16ffc:	data_out=16'hc5;
17'h16ffd:	data_out=16'h9b0;
17'h16ffe:	data_out=16'ha00;
17'h16fff:	data_out=16'h92d;
17'h17000:	data_out=16'h6eb;
17'h17001:	data_out=16'h757;
17'h17002:	data_out=16'ha00;
17'h17003:	data_out=16'ha00;
17'h17004:	data_out=16'h971;
17'h17005:	data_out=16'ha00;
17'h17006:	data_out=16'ha00;
17'h17007:	data_out=16'h90a;
17'h17008:	data_out=16'ha00;
17'h17009:	data_out=16'ha00;
17'h1700a:	data_out=16'h9f9;
17'h1700b:	data_out=16'ha00;
17'h1700c:	data_out=16'ha00;
17'h1700d:	data_out=16'ha00;
17'h1700e:	data_out=16'h513;
17'h1700f:	data_out=16'h9ff;
17'h17010:	data_out=16'ha00;
17'h17011:	data_out=16'ha00;
17'h17012:	data_out=16'h928;
17'h17013:	data_out=16'ha00;
17'h17014:	data_out=16'ha00;
17'h17015:	data_out=16'h9f5;
17'h17016:	data_out=16'ha00;
17'h17017:	data_out=16'ha00;
17'h17018:	data_out=16'h173;
17'h17019:	data_out=16'ha00;
17'h1701a:	data_out=16'ha00;
17'h1701b:	data_out=16'ha00;
17'h1701c:	data_out=16'ha00;
17'h1701d:	data_out=16'h834;
17'h1701e:	data_out=16'ha00;
17'h1701f:	data_out=16'ha00;
17'h17020:	data_out=16'h91d;
17'h17021:	data_out=16'h536;
17'h17022:	data_out=16'ha00;
17'h17023:	data_out=16'h195;
17'h17024:	data_out=16'h196;
17'h17025:	data_out=16'ha00;
17'h17026:	data_out=16'ha00;
17'h17027:	data_out=16'h9d7;
17'h17028:	data_out=16'h5c8;
17'h17029:	data_out=16'ha00;
17'h1702a:	data_out=16'h97c;
17'h1702b:	data_out=16'ha00;
17'h1702c:	data_out=16'ha00;
17'h1702d:	data_out=16'h9ff;
17'h1702e:	data_out=16'ha00;
17'h1702f:	data_out=16'ha00;
17'h17030:	data_out=16'ha00;
17'h17031:	data_out=16'h9fc;
17'h17032:	data_out=16'ha00;
17'h17033:	data_out=16'ha00;
17'h17034:	data_out=16'h52a;
17'h17035:	data_out=16'ha00;
17'h17036:	data_out=16'h9fc;
17'h17037:	data_out=16'ha00;
17'h17038:	data_out=16'h9ff;
17'h17039:	data_out=16'ha00;
17'h1703a:	data_out=16'ha00;
17'h1703b:	data_out=16'h9fc;
17'h1703c:	data_out=16'ha00;
17'h1703d:	data_out=16'h9fe;
17'h1703e:	data_out=16'h5cf;
17'h1703f:	data_out=16'ha00;
17'h17040:	data_out=16'ha00;
17'h17041:	data_out=16'ha00;
17'h17042:	data_out=16'ha00;
17'h17043:	data_out=16'ha00;
17'h17044:	data_out=16'h9f9;
17'h17045:	data_out=16'h9f9;
17'h17046:	data_out=16'ha00;
17'h17047:	data_out=16'h8ce;
17'h17048:	data_out=16'h9fb;
17'h17049:	data_out=16'ha00;
17'h1704a:	data_out=16'h84a;
17'h1704b:	data_out=16'ha00;
17'h1704c:	data_out=16'ha00;
17'h1704d:	data_out=16'ha00;
17'h1704e:	data_out=16'h9ee;
17'h1704f:	data_out=16'ha00;
17'h17050:	data_out=16'ha00;
17'h17051:	data_out=16'h9ff;
17'h17052:	data_out=16'h27b;
17'h17053:	data_out=16'h9e6;
17'h17054:	data_out=16'h878;
17'h17055:	data_out=16'ha00;
17'h17056:	data_out=16'ha00;
17'h17057:	data_out=16'h9ff;
17'h17058:	data_out=16'ha00;
17'h17059:	data_out=16'ha00;
17'h1705a:	data_out=16'ha00;
17'h1705b:	data_out=16'h9ff;
17'h1705c:	data_out=16'ha00;
17'h1705d:	data_out=16'h9fa;
17'h1705e:	data_out=16'ha00;
17'h1705f:	data_out=16'h7ca;
17'h17060:	data_out=16'ha00;
17'h17061:	data_out=16'ha00;
17'h17062:	data_out=16'ha00;
17'h17063:	data_out=16'ha00;
17'h17064:	data_out=16'h8bd;
17'h17065:	data_out=16'ha00;
17'h17066:	data_out=16'ha00;
17'h17067:	data_out=16'ha00;
17'h17068:	data_out=16'h55f;
17'h17069:	data_out=16'ha00;
17'h1706a:	data_out=16'h4fb;
17'h1706b:	data_out=16'ha00;
17'h1706c:	data_out=16'h31f;
17'h1706d:	data_out=16'ha00;
17'h1706e:	data_out=16'h4fb;
17'h1706f:	data_out=16'ha00;
17'h17070:	data_out=16'h508;
17'h17071:	data_out=16'h8bd;
17'h17072:	data_out=16'ha00;
17'h17073:	data_out=16'ha00;
17'h17074:	data_out=16'ha00;
17'h17075:	data_out=16'ha00;
17'h17076:	data_out=16'ha00;
17'h17077:	data_out=16'ha00;
17'h17078:	data_out=16'ha00;
17'h17079:	data_out=16'h9d5;
17'h1707a:	data_out=16'ha00;
17'h1707b:	data_out=16'h5d2;
17'h1707c:	data_out=16'hb4;
17'h1707d:	data_out=16'h9af;
17'h1707e:	data_out=16'ha00;
17'h1707f:	data_out=16'h954;
17'h17080:	data_out=16'h787;
17'h17081:	data_out=16'h6d2;
17'h17082:	data_out=16'ha00;
17'h17083:	data_out=16'ha00;
17'h17084:	data_out=16'h9df;
17'h17085:	data_out=16'ha00;
17'h17086:	data_out=16'ha00;
17'h17087:	data_out=16'h831;
17'h17088:	data_out=16'ha00;
17'h17089:	data_out=16'ha00;
17'h1708a:	data_out=16'h9ef;
17'h1708b:	data_out=16'ha00;
17'h1708c:	data_out=16'ha00;
17'h1708d:	data_out=16'h9fd;
17'h1708e:	data_out=16'h7f5;
17'h1708f:	data_out=16'ha00;
17'h17090:	data_out=16'ha00;
17'h17091:	data_out=16'ha00;
17'h17092:	data_out=16'h94f;
17'h17093:	data_out=16'ha00;
17'h17094:	data_out=16'ha00;
17'h17095:	data_out=16'h9fe;
17'h17096:	data_out=16'ha00;
17'h17097:	data_out=16'ha00;
17'h17098:	data_out=16'ha6;
17'h17099:	data_out=16'ha00;
17'h1709a:	data_out=16'ha00;
17'h1709b:	data_out=16'ha00;
17'h1709c:	data_out=16'ha00;
17'h1709d:	data_out=16'h856;
17'h1709e:	data_out=16'ha00;
17'h1709f:	data_out=16'h9fe;
17'h170a0:	data_out=16'h9ef;
17'h170a1:	data_out=16'h826;
17'h170a2:	data_out=16'ha00;
17'h170a3:	data_out=16'h79e;
17'h170a4:	data_out=16'h7a4;
17'h170a5:	data_out=16'ha00;
17'h170a6:	data_out=16'ha00;
17'h170a7:	data_out=16'ha00;
17'h170a8:	data_out=16'h8f3;
17'h170a9:	data_out=16'ha00;
17'h170aa:	data_out=16'h9fa;
17'h170ab:	data_out=16'ha00;
17'h170ac:	data_out=16'ha00;
17'h170ad:	data_out=16'ha00;
17'h170ae:	data_out=16'ha00;
17'h170af:	data_out=16'ha00;
17'h170b0:	data_out=16'ha00;
17'h170b1:	data_out=16'h99e;
17'h170b2:	data_out=16'ha00;
17'h170b3:	data_out=16'ha00;
17'h170b4:	data_out=16'h400;
17'h170b5:	data_out=16'ha00;
17'h170b6:	data_out=16'ha00;
17'h170b7:	data_out=16'ha00;
17'h170b8:	data_out=16'ha00;
17'h170b9:	data_out=16'ha00;
17'h170ba:	data_out=16'h283;
17'h170bb:	data_out=16'h9ff;
17'h170bc:	data_out=16'ha00;
17'h170bd:	data_out=16'ha00;
17'h170be:	data_out=16'h8fe;
17'h170bf:	data_out=16'ha00;
17'h170c0:	data_out=16'ha00;
17'h170c1:	data_out=16'ha00;
17'h170c2:	data_out=16'ha00;
17'h170c3:	data_out=16'ha00;
17'h170c4:	data_out=16'h9ff;
17'h170c5:	data_out=16'h9fe;
17'h170c6:	data_out=16'ha00;
17'h170c7:	data_out=16'h853;
17'h170c8:	data_out=16'h9fe;
17'h170c9:	data_out=16'ha00;
17'h170ca:	data_out=16'h7b7;
17'h170cb:	data_out=16'ha00;
17'h170cc:	data_out=16'ha00;
17'h170cd:	data_out=16'ha00;
17'h170ce:	data_out=16'ha00;
17'h170cf:	data_out=16'ha00;
17'h170d0:	data_out=16'ha00;
17'h170d1:	data_out=16'h9f4;
17'h170d2:	data_out=16'h942;
17'h170d3:	data_out=16'ha00;
17'h170d4:	data_out=16'h9af;
17'h170d5:	data_out=16'ha00;
17'h170d6:	data_out=16'ha00;
17'h170d7:	data_out=16'h9f7;
17'h170d8:	data_out=16'ha00;
17'h170d9:	data_out=16'ha00;
17'h170da:	data_out=16'ha00;
17'h170db:	data_out=16'ha00;
17'h170dc:	data_out=16'ha00;
17'h170dd:	data_out=16'ha00;
17'h170de:	data_out=16'ha00;
17'h170df:	data_out=16'h5d2;
17'h170e0:	data_out=16'ha00;
17'h170e1:	data_out=16'ha00;
17'h170e2:	data_out=16'ha00;
17'h170e3:	data_out=16'ha00;
17'h170e4:	data_out=16'h8eb;
17'h170e5:	data_out=16'ha00;
17'h170e6:	data_out=16'ha00;
17'h170e7:	data_out=16'ha00;
17'h170e8:	data_out=16'h860;
17'h170e9:	data_out=16'ha00;
17'h170ea:	data_out=16'h7d7;
17'h170eb:	data_out=16'ha00;
17'h170ec:	data_out=16'h83e9;
17'h170ed:	data_out=16'ha00;
17'h170ee:	data_out=16'h7d7;
17'h170ef:	data_out=16'ha00;
17'h170f0:	data_out=16'h7e8;
17'h170f1:	data_out=16'h80ba;
17'h170f2:	data_out=16'ha00;
17'h170f3:	data_out=16'ha00;
17'h170f4:	data_out=16'ha00;
17'h170f5:	data_out=16'ha00;
17'h170f6:	data_out=16'ha00;
17'h170f7:	data_out=16'ha00;
17'h170f8:	data_out=16'ha00;
17'h170f9:	data_out=16'h9fe;
17'h170fa:	data_out=16'ha00;
17'h170fb:	data_out=16'h901;
17'h170fc:	data_out=16'h82fd;
17'h170fd:	data_out=16'h8d2;
17'h170fe:	data_out=16'ha00;
17'h170ff:	data_out=16'h9a6;
17'h17100:	data_out=16'h815;
17'h17101:	data_out=16'h745;
17'h17102:	data_out=16'ha00;
17'h17103:	data_out=16'ha00;
17'h17104:	data_out=16'h9fc;
17'h17105:	data_out=16'ha00;
17'h17106:	data_out=16'ha00;
17'h17107:	data_out=16'h814;
17'h17108:	data_out=16'ha00;
17'h17109:	data_out=16'ha00;
17'h1710a:	data_out=16'h9f7;
17'h1710b:	data_out=16'ha00;
17'h1710c:	data_out=16'ha00;
17'h1710d:	data_out=16'h9f7;
17'h1710e:	data_out=16'ha00;
17'h1710f:	data_out=16'ha00;
17'h17110:	data_out=16'ha00;
17'h17111:	data_out=16'ha00;
17'h17112:	data_out=16'h8da;
17'h17113:	data_out=16'ha00;
17'h17114:	data_out=16'ha00;
17'h17115:	data_out=16'ha00;
17'h17116:	data_out=16'ha00;
17'h17117:	data_out=16'ha00;
17'h17118:	data_out=16'h136;
17'h17119:	data_out=16'ha00;
17'h1711a:	data_out=16'ha00;
17'h1711b:	data_out=16'ha00;
17'h1711c:	data_out=16'ha00;
17'h1711d:	data_out=16'h917;
17'h1711e:	data_out=16'ha00;
17'h1711f:	data_out=16'h9ff;
17'h17120:	data_out=16'ha00;
17'h17121:	data_out=16'ha00;
17'h17122:	data_out=16'ha00;
17'h17123:	data_out=16'h9ff;
17'h17124:	data_out=16'ha00;
17'h17125:	data_out=16'ha00;
17'h17126:	data_out=16'ha00;
17'h17127:	data_out=16'ha00;
17'h17128:	data_out=16'ha00;
17'h17129:	data_out=16'ha00;
17'h1712a:	data_out=16'h8b5;
17'h1712b:	data_out=16'ha00;
17'h1712c:	data_out=16'ha00;
17'h1712d:	data_out=16'ha00;
17'h1712e:	data_out=16'h919;
17'h1712f:	data_out=16'ha00;
17'h17130:	data_out=16'ha00;
17'h17131:	data_out=16'h9ff;
17'h17132:	data_out=16'ha00;
17'h17133:	data_out=16'ha00;
17'h17134:	data_out=16'h43d;
17'h17135:	data_out=16'ha00;
17'h17136:	data_out=16'ha00;
17'h17137:	data_out=16'ha00;
17'h17138:	data_out=16'ha00;
17'h17139:	data_out=16'ha00;
17'h1713a:	data_out=16'h83e8;
17'h1713b:	data_out=16'ha00;
17'h1713c:	data_out=16'ha00;
17'h1713d:	data_out=16'ha00;
17'h1713e:	data_out=16'ha00;
17'h1713f:	data_out=16'ha00;
17'h17140:	data_out=16'ha00;
17'h17141:	data_out=16'ha00;
17'h17142:	data_out=16'ha00;
17'h17143:	data_out=16'h9fd;
17'h17144:	data_out=16'h9ff;
17'h17145:	data_out=16'ha00;
17'h17146:	data_out=16'ha00;
17'h17147:	data_out=16'h72b;
17'h17148:	data_out=16'h9df;
17'h17149:	data_out=16'ha00;
17'h1714a:	data_out=16'h64a;
17'h1714b:	data_out=16'ha00;
17'h1714c:	data_out=16'ha00;
17'h1714d:	data_out=16'ha00;
17'h1714e:	data_out=16'ha00;
17'h1714f:	data_out=16'ha00;
17'h17150:	data_out=16'ha00;
17'h17151:	data_out=16'h9f4;
17'h17152:	data_out=16'h9f9;
17'h17153:	data_out=16'ha00;
17'h17154:	data_out=16'ha00;
17'h17155:	data_out=16'ha00;
17'h17156:	data_out=16'ha00;
17'h17157:	data_out=16'h9ff;
17'h17158:	data_out=16'ha00;
17'h17159:	data_out=16'ha00;
17'h1715a:	data_out=16'ha00;
17'h1715b:	data_out=16'ha00;
17'h1715c:	data_out=16'ha00;
17'h1715d:	data_out=16'ha00;
17'h1715e:	data_out=16'ha00;
17'h1715f:	data_out=16'h3b4;
17'h17160:	data_out=16'ha00;
17'h17161:	data_out=16'ha00;
17'h17162:	data_out=16'ha00;
17'h17163:	data_out=16'ha00;
17'h17164:	data_out=16'h926;
17'h17165:	data_out=16'ha00;
17'h17166:	data_out=16'ha00;
17'h17167:	data_out=16'h94f;
17'h17168:	data_out=16'ha00;
17'h17169:	data_out=16'ha00;
17'h1716a:	data_out=16'ha00;
17'h1716b:	data_out=16'ha00;
17'h1716c:	data_out=16'h86f0;
17'h1716d:	data_out=16'ha00;
17'h1716e:	data_out=16'ha00;
17'h1716f:	data_out=16'ha00;
17'h17170:	data_out=16'ha00;
17'h17171:	data_out=16'h80a5;
17'h17172:	data_out=16'ha00;
17'h17173:	data_out=16'ha00;
17'h17174:	data_out=16'ha00;
17'h17175:	data_out=16'ha00;
17'h17176:	data_out=16'ha00;
17'h17177:	data_out=16'ha00;
17'h17178:	data_out=16'ha00;
17'h17179:	data_out=16'h9fd;
17'h1717a:	data_out=16'ha00;
17'h1717b:	data_out=16'ha00;
17'h1717c:	data_out=16'h84bb;
17'h1717d:	data_out=16'h85d;
17'h1717e:	data_out=16'ha00;
17'h1717f:	data_out=16'h9c7;
17'h17180:	data_out=16'h930;
17'h17181:	data_out=16'h87f;
17'h17182:	data_out=16'ha00;
17'h17183:	data_out=16'ha00;
17'h17184:	data_out=16'ha00;
17'h17185:	data_out=16'ha00;
17'h17186:	data_out=16'ha00;
17'h17187:	data_out=16'h908;
17'h17188:	data_out=16'ha00;
17'h17189:	data_out=16'ha00;
17'h1718a:	data_out=16'ha00;
17'h1718b:	data_out=16'h9ff;
17'h1718c:	data_out=16'ha00;
17'h1718d:	data_out=16'h9fa;
17'h1718e:	data_out=16'ha00;
17'h1718f:	data_out=16'ha00;
17'h17190:	data_out=16'ha00;
17'h17191:	data_out=16'ha00;
17'h17192:	data_out=16'h8c1;
17'h17193:	data_out=16'ha00;
17'h17194:	data_out=16'ha00;
17'h17195:	data_out=16'ha00;
17'h17196:	data_out=16'ha00;
17'h17197:	data_out=16'ha00;
17'h17198:	data_out=16'h2ea;
17'h17199:	data_out=16'ha00;
17'h1719a:	data_out=16'ha00;
17'h1719b:	data_out=16'ha00;
17'h1719c:	data_out=16'ha00;
17'h1719d:	data_out=16'ha00;
17'h1719e:	data_out=16'ha00;
17'h1719f:	data_out=16'ha00;
17'h171a0:	data_out=16'ha00;
17'h171a1:	data_out=16'ha00;
17'h171a2:	data_out=16'ha00;
17'h171a3:	data_out=16'ha00;
17'h171a4:	data_out=16'ha00;
17'h171a5:	data_out=16'ha00;
17'h171a6:	data_out=16'ha00;
17'h171a7:	data_out=16'ha00;
17'h171a8:	data_out=16'ha00;
17'h171a9:	data_out=16'ha00;
17'h171aa:	data_out=16'h74f;
17'h171ab:	data_out=16'ha00;
17'h171ac:	data_out=16'ha00;
17'h171ad:	data_out=16'ha00;
17'h171ae:	data_out=16'h940;
17'h171af:	data_out=16'ha00;
17'h171b0:	data_out=16'ha00;
17'h171b1:	data_out=16'ha00;
17'h171b2:	data_out=16'ha00;
17'h171b3:	data_out=16'ha00;
17'h171b4:	data_out=16'h5b4;
17'h171b5:	data_out=16'ha00;
17'h171b6:	data_out=16'ha00;
17'h171b7:	data_out=16'ha00;
17'h171b8:	data_out=16'ha00;
17'h171b9:	data_out=16'ha00;
17'h171ba:	data_out=16'h837d;
17'h171bb:	data_out=16'ha00;
17'h171bc:	data_out=16'ha00;
17'h171bd:	data_out=16'ha00;
17'h171be:	data_out=16'ha00;
17'h171bf:	data_out=16'ha00;
17'h171c0:	data_out=16'ha00;
17'h171c1:	data_out=16'ha00;
17'h171c2:	data_out=16'ha00;
17'h171c3:	data_out=16'h9ff;
17'h171c4:	data_out=16'ha00;
17'h171c5:	data_out=16'ha00;
17'h171c6:	data_out=16'ha00;
17'h171c7:	data_out=16'h6c9;
17'h171c8:	data_out=16'h9fa;
17'h171c9:	data_out=16'ha00;
17'h171ca:	data_out=16'h5fe;
17'h171cb:	data_out=16'ha00;
17'h171cc:	data_out=16'ha00;
17'h171cd:	data_out=16'ha00;
17'h171ce:	data_out=16'ha00;
17'h171cf:	data_out=16'ha00;
17'h171d0:	data_out=16'ha00;
17'h171d1:	data_out=16'ha00;
17'h171d2:	data_out=16'ha00;
17'h171d3:	data_out=16'ha00;
17'h171d4:	data_out=16'ha00;
17'h171d5:	data_out=16'ha00;
17'h171d6:	data_out=16'ha00;
17'h171d7:	data_out=16'ha00;
17'h171d8:	data_out=16'ha00;
17'h171d9:	data_out=16'ha00;
17'h171da:	data_out=16'ha00;
17'h171db:	data_out=16'ha00;
17'h171dc:	data_out=16'ha00;
17'h171dd:	data_out=16'ha00;
17'h171de:	data_out=16'ha00;
17'h171df:	data_out=16'h50e;
17'h171e0:	data_out=16'ha00;
17'h171e1:	data_out=16'ha00;
17'h171e2:	data_out=16'ha00;
17'h171e3:	data_out=16'ha00;
17'h171e4:	data_out=16'h96c;
17'h171e5:	data_out=16'ha00;
17'h171e6:	data_out=16'ha00;
17'h171e7:	data_out=16'h8a9;
17'h171e8:	data_out=16'ha00;
17'h171e9:	data_out=16'ha00;
17'h171ea:	data_out=16'ha00;
17'h171eb:	data_out=16'ha00;
17'h171ec:	data_out=16'h770;
17'h171ed:	data_out=16'ha00;
17'h171ee:	data_out=16'ha00;
17'h171ef:	data_out=16'ha00;
17'h171f0:	data_out=16'ha00;
17'h171f1:	data_out=16'h8182;
17'h171f2:	data_out=16'ha00;
17'h171f3:	data_out=16'ha00;
17'h171f4:	data_out=16'ha00;
17'h171f5:	data_out=16'ha00;
17'h171f6:	data_out=16'ha00;
17'h171f7:	data_out=16'ha00;
17'h171f8:	data_out=16'ha00;
17'h171f9:	data_out=16'h9ff;
17'h171fa:	data_out=16'ha00;
17'h171fb:	data_out=16'ha00;
17'h171fc:	data_out=16'h8429;
17'h171fd:	data_out=16'h8a9;
17'h171fe:	data_out=16'ha00;
17'h171ff:	data_out=16'h9fa;
17'h17200:	data_out=16'h985;
17'h17201:	data_out=16'h850;
17'h17202:	data_out=16'ha00;
17'h17203:	data_out=16'ha00;
17'h17204:	data_out=16'ha00;
17'h17205:	data_out=16'ha00;
17'h17206:	data_out=16'ha00;
17'h17207:	data_out=16'h9ab;
17'h17208:	data_out=16'ha00;
17'h17209:	data_out=16'ha00;
17'h1720a:	data_out=16'ha00;
17'h1720b:	data_out=16'ha00;
17'h1720c:	data_out=16'ha00;
17'h1720d:	data_out=16'ha00;
17'h1720e:	data_out=16'ha00;
17'h1720f:	data_out=16'ha00;
17'h17210:	data_out=16'ha00;
17'h17211:	data_out=16'ha00;
17'h17212:	data_out=16'h7cb;
17'h17213:	data_out=16'ha00;
17'h17214:	data_out=16'ha00;
17'h17215:	data_out=16'ha00;
17'h17216:	data_out=16'ha00;
17'h17217:	data_out=16'ha00;
17'h17218:	data_out=16'h235;
17'h17219:	data_out=16'ha00;
17'h1721a:	data_out=16'ha00;
17'h1721b:	data_out=16'ha00;
17'h1721c:	data_out=16'ha00;
17'h1721d:	data_out=16'ha00;
17'h1721e:	data_out=16'ha00;
17'h1721f:	data_out=16'ha00;
17'h17220:	data_out=16'ha00;
17'h17221:	data_out=16'ha00;
17'h17222:	data_out=16'ha00;
17'h17223:	data_out=16'ha00;
17'h17224:	data_out=16'ha00;
17'h17225:	data_out=16'ha00;
17'h17226:	data_out=16'ha00;
17'h17227:	data_out=16'ha00;
17'h17228:	data_out=16'ha00;
17'h17229:	data_out=16'ha00;
17'h1722a:	data_out=16'h754;
17'h1722b:	data_out=16'ha00;
17'h1722c:	data_out=16'ha00;
17'h1722d:	data_out=16'ha00;
17'h1722e:	data_out=16'h855;
17'h1722f:	data_out=16'ha00;
17'h17230:	data_out=16'ha00;
17'h17231:	data_out=16'ha00;
17'h17232:	data_out=16'ha00;
17'h17233:	data_out=16'ha00;
17'h17234:	data_out=16'h5ba;
17'h17235:	data_out=16'ha00;
17'h17236:	data_out=16'ha00;
17'h17237:	data_out=16'ha00;
17'h17238:	data_out=16'ha00;
17'h17239:	data_out=16'ha00;
17'h1723a:	data_out=16'h4c0;
17'h1723b:	data_out=16'ha00;
17'h1723c:	data_out=16'ha00;
17'h1723d:	data_out=16'ha00;
17'h1723e:	data_out=16'ha00;
17'h1723f:	data_out=16'ha00;
17'h17240:	data_out=16'ha00;
17'h17241:	data_out=16'ha00;
17'h17242:	data_out=16'ha00;
17'h17243:	data_out=16'h9ff;
17'h17244:	data_out=16'ha00;
17'h17245:	data_out=16'ha00;
17'h17246:	data_out=16'ha00;
17'h17247:	data_out=16'h81b;
17'h17248:	data_out=16'h7ef;
17'h17249:	data_out=16'ha00;
17'h1724a:	data_out=16'h3fc;
17'h1724b:	data_out=16'ha00;
17'h1724c:	data_out=16'ha00;
17'h1724d:	data_out=16'ha00;
17'h1724e:	data_out=16'h9ff;
17'h1724f:	data_out=16'ha00;
17'h17250:	data_out=16'ha00;
17'h17251:	data_out=16'ha00;
17'h17252:	data_out=16'ha00;
17'h17253:	data_out=16'ha00;
17'h17254:	data_out=16'ha00;
17'h17255:	data_out=16'ha00;
17'h17256:	data_out=16'ha00;
17'h17257:	data_out=16'ha00;
17'h17258:	data_out=16'ha00;
17'h17259:	data_out=16'ha00;
17'h1725a:	data_out=16'ha00;
17'h1725b:	data_out=16'ha00;
17'h1725c:	data_out=16'ha00;
17'h1725d:	data_out=16'ha00;
17'h1725e:	data_out=16'ha00;
17'h1725f:	data_out=16'h2e3;
17'h17260:	data_out=16'ha00;
17'h17261:	data_out=16'ha00;
17'h17262:	data_out=16'ha00;
17'h17263:	data_out=16'ha00;
17'h17264:	data_out=16'h9fb;
17'h17265:	data_out=16'ha00;
17'h17266:	data_out=16'ha00;
17'h17267:	data_out=16'ha00;
17'h17268:	data_out=16'ha00;
17'h17269:	data_out=16'ha00;
17'h1726a:	data_out=16'ha00;
17'h1726b:	data_out=16'ha00;
17'h1726c:	data_out=16'h92;
17'h1726d:	data_out=16'ha00;
17'h1726e:	data_out=16'ha00;
17'h1726f:	data_out=16'ha00;
17'h17270:	data_out=16'ha00;
17'h17271:	data_out=16'h84e4;
17'h17272:	data_out=16'ha00;
17'h17273:	data_out=16'ha00;
17'h17274:	data_out=16'ha00;
17'h17275:	data_out=16'ha00;
17'h17276:	data_out=16'ha00;
17'h17277:	data_out=16'ha00;
17'h17278:	data_out=16'ha00;
17'h17279:	data_out=16'h9fe;
17'h1727a:	data_out=16'ha00;
17'h1727b:	data_out=16'ha00;
17'h1727c:	data_out=16'h877d;
17'h1727d:	data_out=16'h832;
17'h1727e:	data_out=16'ha00;
17'h1727f:	data_out=16'h994;
17'h17280:	data_out=16'h9b1;
17'h17281:	data_out=16'h9e9;
17'h17282:	data_out=16'ha00;
17'h17283:	data_out=16'ha00;
17'h17284:	data_out=16'ha00;
17'h17285:	data_out=16'ha00;
17'h17286:	data_out=16'ha00;
17'h17287:	data_out=16'h9c0;
17'h17288:	data_out=16'ha00;
17'h17289:	data_out=16'ha00;
17'h1728a:	data_out=16'h9ef;
17'h1728b:	data_out=16'ha00;
17'h1728c:	data_out=16'ha00;
17'h1728d:	data_out=16'ha00;
17'h1728e:	data_out=16'ha00;
17'h1728f:	data_out=16'h9f0;
17'h17290:	data_out=16'ha00;
17'h17291:	data_out=16'ha00;
17'h17292:	data_out=16'h9b1;
17'h17293:	data_out=16'ha00;
17'h17294:	data_out=16'ha00;
17'h17295:	data_out=16'ha00;
17'h17296:	data_out=16'ha00;
17'h17297:	data_out=16'ha00;
17'h17298:	data_out=16'hce;
17'h17299:	data_out=16'ha00;
17'h1729a:	data_out=16'ha00;
17'h1729b:	data_out=16'ha00;
17'h1729c:	data_out=16'ha00;
17'h1729d:	data_out=16'h9f3;
17'h1729e:	data_out=16'ha00;
17'h1729f:	data_out=16'h9f3;
17'h172a0:	data_out=16'h9f3;
17'h172a1:	data_out=16'ha00;
17'h172a2:	data_out=16'ha00;
17'h172a3:	data_out=16'ha00;
17'h172a4:	data_out=16'ha00;
17'h172a5:	data_out=16'ha00;
17'h172a6:	data_out=16'ha00;
17'h172a7:	data_out=16'ha00;
17'h172a8:	data_out=16'ha00;
17'h172a9:	data_out=16'ha00;
17'h172aa:	data_out=16'h95a;
17'h172ab:	data_out=16'ha00;
17'h172ac:	data_out=16'ha00;
17'h172ad:	data_out=16'ha00;
17'h172ae:	data_out=16'h9fd;
17'h172af:	data_out=16'ha00;
17'h172b0:	data_out=16'ha00;
17'h172b1:	data_out=16'h8cd;
17'h172b2:	data_out=16'ha00;
17'h172b3:	data_out=16'ha00;
17'h172b4:	data_out=16'h7cd;
17'h172b5:	data_out=16'ha00;
17'h172b6:	data_out=16'h9fc;
17'h172b7:	data_out=16'ha00;
17'h172b8:	data_out=16'ha00;
17'h172b9:	data_out=16'ha00;
17'h172ba:	data_out=16'ha00;
17'h172bb:	data_out=16'ha00;
17'h172bc:	data_out=16'ha00;
17'h172bd:	data_out=16'ha00;
17'h172be:	data_out=16'ha00;
17'h172bf:	data_out=16'ha00;
17'h172c0:	data_out=16'ha00;
17'h172c1:	data_out=16'ha00;
17'h172c2:	data_out=16'ha00;
17'h172c3:	data_out=16'h9ff;
17'h172c4:	data_out=16'ha00;
17'h172c5:	data_out=16'ha00;
17'h172c6:	data_out=16'ha00;
17'h172c7:	data_out=16'h9bf;
17'h172c8:	data_out=16'h9f8;
17'h172c9:	data_out=16'ha00;
17'h172ca:	data_out=16'h872;
17'h172cb:	data_out=16'ha00;
17'h172cc:	data_out=16'ha00;
17'h172cd:	data_out=16'ha00;
17'h172ce:	data_out=16'h9ff;
17'h172cf:	data_out=16'ha00;
17'h172d0:	data_out=16'ha00;
17'h172d1:	data_out=16'ha00;
17'h172d2:	data_out=16'ha00;
17'h172d3:	data_out=16'h9fb;
17'h172d4:	data_out=16'h9e6;
17'h172d5:	data_out=16'ha00;
17'h172d6:	data_out=16'ha00;
17'h172d7:	data_out=16'ha00;
17'h172d8:	data_out=16'ha00;
17'h172d9:	data_out=16'ha00;
17'h172da:	data_out=16'ha00;
17'h172db:	data_out=16'ha00;
17'h172dc:	data_out=16'ha00;
17'h172dd:	data_out=16'h9ff;
17'h172de:	data_out=16'ha00;
17'h172df:	data_out=16'h5ed;
17'h172e0:	data_out=16'ha00;
17'h172e1:	data_out=16'ha00;
17'h172e2:	data_out=16'ha00;
17'h172e3:	data_out=16'ha00;
17'h172e4:	data_out=16'h9f1;
17'h172e5:	data_out=16'ha00;
17'h172e6:	data_out=16'ha00;
17'h172e7:	data_out=16'h9f9;
17'h172e8:	data_out=16'ha00;
17'h172e9:	data_out=16'ha00;
17'h172ea:	data_out=16'ha00;
17'h172eb:	data_out=16'ha00;
17'h172ec:	data_out=16'h3c4;
17'h172ed:	data_out=16'ha00;
17'h172ee:	data_out=16'ha00;
17'h172ef:	data_out=16'ha00;
17'h172f0:	data_out=16'ha00;
17'h172f1:	data_out=16'h81dd;
17'h172f2:	data_out=16'ha00;
17'h172f3:	data_out=16'ha00;
17'h172f4:	data_out=16'ha00;
17'h172f5:	data_out=16'ha00;
17'h172f6:	data_out=16'ha00;
17'h172f7:	data_out=16'ha00;
17'h172f8:	data_out=16'ha00;
17'h172f9:	data_out=16'h9fa;
17'h172fa:	data_out=16'ha00;
17'h172fb:	data_out=16'ha00;
17'h172fc:	data_out=16'h8775;
17'h172fd:	data_out=16'h7bb;
17'h172fe:	data_out=16'ha00;
17'h172ff:	data_out=16'h90e;
17'h17300:	data_out=16'h9ef;
17'h17301:	data_out=16'h9b5;
17'h17302:	data_out=16'ha00;
17'h17303:	data_out=16'ha00;
17'h17304:	data_out=16'h8e7;
17'h17305:	data_out=16'h943;
17'h17306:	data_out=16'ha00;
17'h17307:	data_out=16'h950;
17'h17308:	data_out=16'ha00;
17'h17309:	data_out=16'ha00;
17'h1730a:	data_out=16'h92d;
17'h1730b:	data_out=16'ha00;
17'h1730c:	data_out=16'ha00;
17'h1730d:	data_out=16'ha00;
17'h1730e:	data_out=16'ha00;
17'h1730f:	data_out=16'h9f1;
17'h17310:	data_out=16'ha00;
17'h17311:	data_out=16'h9fd;
17'h17312:	data_out=16'h9f8;
17'h17313:	data_out=16'ha00;
17'h17314:	data_out=16'ha00;
17'h17315:	data_out=16'h9c9;
17'h17316:	data_out=16'h9fb;
17'h17317:	data_out=16'ha00;
17'h17318:	data_out=16'h83e9;
17'h17319:	data_out=16'ha00;
17'h1731a:	data_out=16'h95e;
17'h1731b:	data_out=16'ha00;
17'h1731c:	data_out=16'ha00;
17'h1731d:	data_out=16'h9ed;
17'h1731e:	data_out=16'ha00;
17'h1731f:	data_out=16'h927;
17'h17320:	data_out=16'h9ed;
17'h17321:	data_out=16'ha00;
17'h17322:	data_out=16'ha00;
17'h17323:	data_out=16'h2ca;
17'h17324:	data_out=16'h2b8;
17'h17325:	data_out=16'ha00;
17'h17326:	data_out=16'ha00;
17'h17327:	data_out=16'h9f8;
17'h17328:	data_out=16'ha00;
17'h17329:	data_out=16'ha00;
17'h1732a:	data_out=16'h9be;
17'h1732b:	data_out=16'h9ff;
17'h1732c:	data_out=16'h9f7;
17'h1732d:	data_out=16'ha00;
17'h1732e:	data_out=16'h9ff;
17'h1732f:	data_out=16'ha00;
17'h17330:	data_out=16'ha00;
17'h17331:	data_out=16'h831;
17'h17332:	data_out=16'h9fb;
17'h17333:	data_out=16'ha00;
17'h17334:	data_out=16'h991;
17'h17335:	data_out=16'h9fd;
17'h17336:	data_out=16'h9fc;
17'h17337:	data_out=16'ha00;
17'h17338:	data_out=16'ha00;
17'h17339:	data_out=16'ha00;
17'h1733a:	data_out=16'ha00;
17'h1733b:	data_out=16'h99a;
17'h1733c:	data_out=16'ha00;
17'h1733d:	data_out=16'h9fa;
17'h1733e:	data_out=16'ha00;
17'h1733f:	data_out=16'h93e;
17'h17340:	data_out=16'h9fb;
17'h17341:	data_out=16'ha00;
17'h17342:	data_out=16'ha00;
17'h17343:	data_out=16'ha00;
17'h17344:	data_out=16'h923;
17'h17345:	data_out=16'h9c7;
17'h17346:	data_out=16'ha00;
17'h17347:	data_out=16'h9e1;
17'h17348:	data_out=16'h9fd;
17'h17349:	data_out=16'ha00;
17'h1734a:	data_out=16'h942;
17'h1734b:	data_out=16'ha00;
17'h1734c:	data_out=16'ha00;
17'h1734d:	data_out=16'ha00;
17'h1734e:	data_out=16'ha00;
17'h1734f:	data_out=16'ha00;
17'h17350:	data_out=16'ha00;
17'h17351:	data_out=16'h9f8;
17'h17352:	data_out=16'h66b;
17'h17353:	data_out=16'h9fa;
17'h17354:	data_out=16'h9f5;
17'h17355:	data_out=16'ha00;
17'h17356:	data_out=16'ha00;
17'h17357:	data_out=16'h9fd;
17'h17358:	data_out=16'ha00;
17'h17359:	data_out=16'h9f7;
17'h1735a:	data_out=16'ha00;
17'h1735b:	data_out=16'h9ca;
17'h1735c:	data_out=16'ha00;
17'h1735d:	data_out=16'ha00;
17'h1735e:	data_out=16'ha00;
17'h1735f:	data_out=16'h5dc;
17'h17360:	data_out=16'ha00;
17'h17361:	data_out=16'h9f9;
17'h17362:	data_out=16'ha00;
17'h17363:	data_out=16'ha00;
17'h17364:	data_out=16'ha00;
17'h17365:	data_out=16'h9f8;
17'h17366:	data_out=16'ha00;
17'h17367:	data_out=16'h9f9;
17'h17368:	data_out=16'ha00;
17'h17369:	data_out=16'ha00;
17'h1736a:	data_out=16'ha00;
17'h1736b:	data_out=16'h9d8;
17'h1736c:	data_out=16'h890;
17'h1736d:	data_out=16'ha00;
17'h1736e:	data_out=16'ha00;
17'h1736f:	data_out=16'h9f7;
17'h17370:	data_out=16'ha00;
17'h17371:	data_out=16'h88c9;
17'h17372:	data_out=16'h9b3;
17'h17373:	data_out=16'h9d1;
17'h17374:	data_out=16'ha00;
17'h17375:	data_out=16'h9ff;
17'h17376:	data_out=16'ha00;
17'h17377:	data_out=16'ha00;
17'h17378:	data_out=16'ha00;
17'h17379:	data_out=16'h9fb;
17'h1737a:	data_out=16'ha00;
17'h1737b:	data_out=16'ha00;
17'h1737c:	data_out=16'h8a00;
17'h1737d:	data_out=16'h694;
17'h1737e:	data_out=16'ha00;
17'h1737f:	data_out=16'h8d5;
17'h17380:	data_out=16'ha00;
17'h17381:	data_out=16'h9de;
17'h17382:	data_out=16'ha00;
17'h17383:	data_out=16'ha00;
17'h17384:	data_out=16'h979;
17'h17385:	data_out=16'h9d6;
17'h17386:	data_out=16'h9f8;
17'h17387:	data_out=16'h985;
17'h17388:	data_out=16'ha00;
17'h17389:	data_out=16'ha00;
17'h1738a:	data_out=16'h971;
17'h1738b:	data_out=16'ha00;
17'h1738c:	data_out=16'ha00;
17'h1738d:	data_out=16'ha00;
17'h1738e:	data_out=16'h60a;
17'h1738f:	data_out=16'h9f9;
17'h17390:	data_out=16'ha00;
17'h17391:	data_out=16'h9f7;
17'h17392:	data_out=16'ha00;
17'h17393:	data_out=16'ha00;
17'h17394:	data_out=16'ha00;
17'h17395:	data_out=16'h9fa;
17'h17396:	data_out=16'h9fe;
17'h17397:	data_out=16'ha00;
17'h17398:	data_out=16'h8061;
17'h17399:	data_out=16'h9fc;
17'h1739a:	data_out=16'h9cb;
17'h1739b:	data_out=16'ha00;
17'h1739c:	data_out=16'ha00;
17'h1739d:	data_out=16'h9fb;
17'h1739e:	data_out=16'ha00;
17'h1739f:	data_out=16'h561;
17'h173a0:	data_out=16'h9ff;
17'h173a1:	data_out=16'h63f;
17'h173a2:	data_out=16'ha00;
17'h173a3:	data_out=16'h8a00;
17'h173a4:	data_out=16'h8a00;
17'h173a5:	data_out=16'h9f9;
17'h173a6:	data_out=16'ha00;
17'h173a7:	data_out=16'h9fb;
17'h173a8:	data_out=16'h720;
17'h173a9:	data_out=16'ha00;
17'h173aa:	data_out=16'h9dc;
17'h173ab:	data_out=16'h9ff;
17'h173ac:	data_out=16'h9fb;
17'h173ad:	data_out=16'ha00;
17'h173ae:	data_out=16'h9f8;
17'h173af:	data_out=16'ha00;
17'h173b0:	data_out=16'ha00;
17'h173b1:	data_out=16'h958;
17'h173b2:	data_out=16'h9ef;
17'h173b3:	data_out=16'ha00;
17'h173b4:	data_out=16'h9d0;
17'h173b5:	data_out=16'h9f4;
17'h173b6:	data_out=16'ha00;
17'h173b7:	data_out=16'ha00;
17'h173b8:	data_out=16'ha00;
17'h173b9:	data_out=16'ha00;
17'h173ba:	data_out=16'h9fc;
17'h173bb:	data_out=16'h9d7;
17'h173bc:	data_out=16'ha00;
17'h173bd:	data_out=16'h9ff;
17'h173be:	data_out=16'h72d;
17'h173bf:	data_out=16'h9d3;
17'h173c0:	data_out=16'h9ef;
17'h173c1:	data_out=16'ha00;
17'h173c2:	data_out=16'ha00;
17'h173c3:	data_out=16'h9fa;
17'h173c4:	data_out=16'h9c7;
17'h173c5:	data_out=16'h9fa;
17'h173c6:	data_out=16'ha00;
17'h173c7:	data_out=16'h9e3;
17'h173c8:	data_out=16'h9ff;
17'h173c9:	data_out=16'ha00;
17'h173ca:	data_out=16'h9ed;
17'h173cb:	data_out=16'ha00;
17'h173cc:	data_out=16'h9fc;
17'h173cd:	data_out=16'ha00;
17'h173ce:	data_out=16'ha00;
17'h173cf:	data_out=16'h9fe;
17'h173d0:	data_out=16'ha00;
17'h173d1:	data_out=16'h9fc;
17'h173d2:	data_out=16'h892e;
17'h173d3:	data_out=16'h9ff;
17'h173d4:	data_out=16'h9ff;
17'h173d5:	data_out=16'ha00;
17'h173d6:	data_out=16'ha00;
17'h173d7:	data_out=16'h9bb;
17'h173d8:	data_out=16'ha00;
17'h173d9:	data_out=16'h9e8;
17'h173da:	data_out=16'ha00;
17'h173db:	data_out=16'h9ee;
17'h173dc:	data_out=16'ha00;
17'h173dd:	data_out=16'ha00;
17'h173de:	data_out=16'ha00;
17'h173df:	data_out=16'h9fe;
17'h173e0:	data_out=16'ha00;
17'h173e1:	data_out=16'h9ef;
17'h173e2:	data_out=16'ha00;
17'h173e3:	data_out=16'ha00;
17'h173e4:	data_out=16'ha00;
17'h173e5:	data_out=16'h9eb;
17'h173e6:	data_out=16'h9fd;
17'h173e7:	data_out=16'h9fc;
17'h173e8:	data_out=16'h67b;
17'h173e9:	data_out=16'ha00;
17'h173ea:	data_out=16'h5e0;
17'h173eb:	data_out=16'h9f1;
17'h173ec:	data_out=16'ha00;
17'h173ed:	data_out=16'ha00;
17'h173ee:	data_out=16'h5e0;
17'h173ef:	data_out=16'h9f3;
17'h173f0:	data_out=16'h5f7;
17'h173f1:	data_out=16'h39e;
17'h173f2:	data_out=16'h9e6;
17'h173f3:	data_out=16'h9e8;
17'h173f4:	data_out=16'ha00;
17'h173f5:	data_out=16'h9f9;
17'h173f6:	data_out=16'ha00;
17'h173f7:	data_out=16'ha00;
17'h173f8:	data_out=16'h9ff;
17'h173f9:	data_out=16'ha00;
17'h173fa:	data_out=16'ha00;
17'h173fb:	data_out=16'h731;
17'h173fc:	data_out=16'h837b;
17'h173fd:	data_out=16'h857;
17'h173fe:	data_out=16'ha00;
17'h173ff:	data_out=16'h9a5;
17'h17400:	data_out=16'ha00;
17'h17401:	data_out=16'h9fc;
17'h17402:	data_out=16'h9fe;
17'h17403:	data_out=16'ha00;
17'h17404:	data_out=16'h9e6;
17'h17405:	data_out=16'h9f5;
17'h17406:	data_out=16'h9ef;
17'h17407:	data_out=16'h9c0;
17'h17408:	data_out=16'ha00;
17'h17409:	data_out=16'h9f4;
17'h1740a:	data_out=16'h9a8;
17'h1740b:	data_out=16'ha00;
17'h1740c:	data_out=16'ha00;
17'h1740d:	data_out=16'ha00;
17'h1740e:	data_out=16'h49a;
17'h1740f:	data_out=16'h9f7;
17'h17410:	data_out=16'ha00;
17'h17411:	data_out=16'h9f9;
17'h17412:	data_out=16'ha00;
17'h17413:	data_out=16'ha00;
17'h17414:	data_out=16'ha00;
17'h17415:	data_out=16'h9fb;
17'h17416:	data_out=16'h9fb;
17'h17417:	data_out=16'ha00;
17'h17418:	data_out=16'h812c;
17'h17419:	data_out=16'h9ff;
17'h1741a:	data_out=16'h9f4;
17'h1741b:	data_out=16'ha00;
17'h1741c:	data_out=16'ha00;
17'h1741d:	data_out=16'h9fe;
17'h1741e:	data_out=16'ha00;
17'h1741f:	data_out=16'h497;
17'h17420:	data_out=16'ha00;
17'h17421:	data_out=16'h4c5;
17'h17422:	data_out=16'ha00;
17'h17423:	data_out=16'h89ff;
17'h17424:	data_out=16'h89ff;
17'h17425:	data_out=16'h9ad;
17'h17426:	data_out=16'ha00;
17'h17427:	data_out=16'h9fd;
17'h17428:	data_out=16'h582;
17'h17429:	data_out=16'ha00;
17'h1742a:	data_out=16'h9ef;
17'h1742b:	data_out=16'ha00;
17'h1742c:	data_out=16'h9fa;
17'h1742d:	data_out=16'ha00;
17'h1742e:	data_out=16'h9f8;
17'h1742f:	data_out=16'ha00;
17'h17430:	data_out=16'ha00;
17'h17431:	data_out=16'h9e3;
17'h17432:	data_out=16'h9f4;
17'h17433:	data_out=16'ha00;
17'h17434:	data_out=16'h9fc;
17'h17435:	data_out=16'h9f2;
17'h17436:	data_out=16'ha00;
17'h17437:	data_out=16'h9ff;
17'h17438:	data_out=16'ha00;
17'h17439:	data_out=16'ha00;
17'h1743a:	data_out=16'h9f3;
17'h1743b:	data_out=16'h9f0;
17'h1743c:	data_out=16'ha00;
17'h1743d:	data_out=16'h9f9;
17'h1743e:	data_out=16'h58d;
17'h1743f:	data_out=16'h9f5;
17'h17440:	data_out=16'h9f1;
17'h17441:	data_out=16'ha00;
17'h17442:	data_out=16'ha00;
17'h17443:	data_out=16'h361;
17'h17444:	data_out=16'h9f3;
17'h17445:	data_out=16'h9fb;
17'h17446:	data_out=16'ha00;
17'h17447:	data_out=16'h9ea;
17'h17448:	data_out=16'ha00;
17'h17449:	data_out=16'h9f9;
17'h1744a:	data_out=16'h9fe;
17'h1744b:	data_out=16'ha00;
17'h1744c:	data_out=16'h9f6;
17'h1744d:	data_out=16'ha00;
17'h1744e:	data_out=16'ha00;
17'h1744f:	data_out=16'h9f9;
17'h17450:	data_out=16'ha00;
17'h17451:	data_out=16'h97b;
17'h17452:	data_out=16'h89ff;
17'h17453:	data_out=16'ha00;
17'h17454:	data_out=16'ha00;
17'h17455:	data_out=16'ha00;
17'h17456:	data_out=16'ha00;
17'h17457:	data_out=16'h429;
17'h17458:	data_out=16'ha00;
17'h17459:	data_out=16'h9ec;
17'h1745a:	data_out=16'ha00;
17'h1745b:	data_out=16'h9f4;
17'h1745c:	data_out=16'ha00;
17'h1745d:	data_out=16'ha00;
17'h1745e:	data_out=16'ha00;
17'h1745f:	data_out=16'h9ff;
17'h17460:	data_out=16'ha00;
17'h17461:	data_out=16'h9f4;
17'h17462:	data_out=16'ha00;
17'h17463:	data_out=16'ha00;
17'h17464:	data_out=16'ha00;
17'h17465:	data_out=16'h9ef;
17'h17466:	data_out=16'h9fe;
17'h17467:	data_out=16'h9fe;
17'h17468:	data_out=16'h4f4;
17'h17469:	data_out=16'ha00;
17'h1746a:	data_out=16'h473;
17'h1746b:	data_out=16'h9f5;
17'h1746c:	data_out=16'ha00;
17'h1746d:	data_out=16'ha00;
17'h1746e:	data_out=16'h473;
17'h1746f:	data_out=16'h9f9;
17'h17470:	data_out=16'h48a;
17'h17471:	data_out=16'h785;
17'h17472:	data_out=16'h9ee;
17'h17473:	data_out=16'h9f1;
17'h17474:	data_out=16'ha00;
17'h17475:	data_out=16'h9fb;
17'h17476:	data_out=16'ha00;
17'h17477:	data_out=16'ha00;
17'h17478:	data_out=16'h9f7;
17'h17479:	data_out=16'h9ff;
17'h1747a:	data_out=16'ha00;
17'h1747b:	data_out=16'h591;
17'h1747c:	data_out=16'h814a;
17'h1747d:	data_out=16'h90f;
17'h1747e:	data_out=16'ha00;
17'h1747f:	data_out=16'h9ef;
17'h17480:	data_out=16'ha00;
17'h17481:	data_out=16'ha00;
17'h17482:	data_out=16'ha00;
17'h17483:	data_out=16'h9fe;
17'h17484:	data_out=16'h9ed;
17'h17485:	data_out=16'h9fc;
17'h17486:	data_out=16'h963;
17'h17487:	data_out=16'h9d2;
17'h17488:	data_out=16'ha00;
17'h17489:	data_out=16'h959;
17'h1748a:	data_out=16'h9b2;
17'h1748b:	data_out=16'ha00;
17'h1748c:	data_out=16'ha00;
17'h1748d:	data_out=16'h9fd;
17'h1748e:	data_out=16'h2fe;
17'h1748f:	data_out=16'ha00;
17'h17490:	data_out=16'ha00;
17'h17491:	data_out=16'h9fe;
17'h17492:	data_out=16'ha00;
17'h17493:	data_out=16'h9fb;
17'h17494:	data_out=16'h9fd;
17'h17495:	data_out=16'h9fc;
17'h17496:	data_out=16'h9fb;
17'h17497:	data_out=16'h9ff;
17'h17498:	data_out=16'h81a5;
17'h17499:	data_out=16'ha00;
17'h1749a:	data_out=16'h9fc;
17'h1749b:	data_out=16'ha00;
17'h1749c:	data_out=16'ha00;
17'h1749d:	data_out=16'ha00;
17'h1749e:	data_out=16'ha00;
17'h1749f:	data_out=16'h8446;
17'h174a0:	data_out=16'ha00;
17'h174a1:	data_out=16'h31b;
17'h174a2:	data_out=16'ha00;
17'h174a3:	data_out=16'h89ff;
17'h174a4:	data_out=16'h89ff;
17'h174a5:	data_out=16'h89c;
17'h174a6:	data_out=16'h9fb;
17'h174a7:	data_out=16'ha00;
17'h174a8:	data_out=16'h3a9;
17'h174a9:	data_out=16'ha00;
17'h174aa:	data_out=16'h9fe;
17'h174ab:	data_out=16'ha00;
17'h174ac:	data_out=16'h9fa;
17'h174ad:	data_out=16'ha00;
17'h174ae:	data_out=16'ha00;
17'h174af:	data_out=16'ha00;
17'h174b0:	data_out=16'ha00;
17'h174b1:	data_out=16'h9f9;
17'h174b2:	data_out=16'h9fb;
17'h174b3:	data_out=16'ha00;
17'h174b4:	data_out=16'ha00;
17'h174b5:	data_out=16'h9fb;
17'h174b6:	data_out=16'ha00;
17'h174b7:	data_out=16'ha00;
17'h174b8:	data_out=16'ha00;
17'h174b9:	data_out=16'ha00;
17'h174ba:	data_out=16'h238;
17'h174bb:	data_out=16'h9fb;
17'h174bc:	data_out=16'ha00;
17'h174bd:	data_out=16'ha00;
17'h174be:	data_out=16'h3b2;
17'h174bf:	data_out=16'h9fc;
17'h174c0:	data_out=16'h9f6;
17'h174c1:	data_out=16'ha00;
17'h174c2:	data_out=16'ha00;
17'h174c3:	data_out=16'h8351;
17'h174c4:	data_out=16'h9fc;
17'h174c5:	data_out=16'h9fc;
17'h174c6:	data_out=16'ha00;
17'h174c7:	data_out=16'h498;
17'h174c8:	data_out=16'ha00;
17'h174c9:	data_out=16'h92e;
17'h174ca:	data_out=16'ha00;
17'h174cb:	data_out=16'ha00;
17'h174cc:	data_out=16'h9dc;
17'h174cd:	data_out=16'ha00;
17'h174ce:	data_out=16'ha00;
17'h174cf:	data_out=16'h615;
17'h174d0:	data_out=16'h9fe;
17'h174d1:	data_out=16'h905;
17'h174d2:	data_out=16'h89ff;
17'h174d3:	data_out=16'ha00;
17'h174d4:	data_out=16'ha00;
17'h174d5:	data_out=16'h9fb;
17'h174d6:	data_out=16'h9fc;
17'h174d7:	data_out=16'h80f6;
17'h174d8:	data_out=16'ha00;
17'h174d9:	data_out=16'h9f0;
17'h174da:	data_out=16'ha00;
17'h174db:	data_out=16'h9fd;
17'h174dc:	data_out=16'ha00;
17'h174dd:	data_out=16'ha00;
17'h174de:	data_out=16'ha00;
17'h174df:	data_out=16'ha00;
17'h174e0:	data_out=16'h9fc;
17'h174e1:	data_out=16'h9fa;
17'h174e2:	data_out=16'ha00;
17'h174e3:	data_out=16'ha00;
17'h174e4:	data_out=16'ha00;
17'h174e5:	data_out=16'h9f6;
17'h174e6:	data_out=16'h848;
17'h174e7:	data_out=16'ha00;
17'h174e8:	data_out=16'h33b;
17'h174e9:	data_out=16'ha00;
17'h174ea:	data_out=16'h2de;
17'h174eb:	data_out=16'h9fa;
17'h174ec:	data_out=16'ha00;
17'h174ed:	data_out=16'ha00;
17'h174ee:	data_out=16'h2df;
17'h174ef:	data_out=16'h9ff;
17'h174f0:	data_out=16'h2f1;
17'h174f1:	data_out=16'h5c4;
17'h174f2:	data_out=16'h9f2;
17'h174f3:	data_out=16'h9f6;
17'h174f4:	data_out=16'ha00;
17'h174f5:	data_out=16'h9fc;
17'h174f6:	data_out=16'ha00;
17'h174f7:	data_out=16'ha00;
17'h174f8:	data_out=16'h861;
17'h174f9:	data_out=16'ha00;
17'h174fa:	data_out=16'ha00;
17'h174fb:	data_out=16'h3b5;
17'h174fc:	data_out=16'h8061;
17'h174fd:	data_out=16'h467;
17'h174fe:	data_out=16'h9ec;
17'h174ff:	data_out=16'h9fc;
17'h17500:	data_out=16'ha00;
17'h17501:	data_out=16'ha00;
17'h17502:	data_out=16'ha00;
17'h17503:	data_out=16'h9fc;
17'h17504:	data_out=16'h987;
17'h17505:	data_out=16'h9e4;
17'h17506:	data_out=16'h66a;
17'h17507:	data_out=16'h13d;
17'h17508:	data_out=16'ha00;
17'h17509:	data_out=16'h76a;
17'h1750a:	data_out=16'h968;
17'h1750b:	data_out=16'ha00;
17'h1750c:	data_out=16'ha00;
17'h1750d:	data_out=16'h9fa;
17'h1750e:	data_out=16'h18b;
17'h1750f:	data_out=16'h9fe;
17'h17510:	data_out=16'h9fd;
17'h17511:	data_out=16'h9f2;
17'h17512:	data_out=16'ha00;
17'h17513:	data_out=16'h9f9;
17'h17514:	data_out=16'h9ff;
17'h17515:	data_out=16'h7a0;
17'h17516:	data_out=16'h9fa;
17'h17517:	data_out=16'ha00;
17'h17518:	data_out=16'h8303;
17'h17519:	data_out=16'ha00;
17'h1751a:	data_out=16'h9dd;
17'h1751b:	data_out=16'ha00;
17'h1751c:	data_out=16'ha00;
17'h1751d:	data_out=16'ha00;
17'h1751e:	data_out=16'ha00;
17'h1751f:	data_out=16'h89d2;
17'h17520:	data_out=16'ha00;
17'h17521:	data_out=16'h1a7;
17'h17522:	data_out=16'ha00;
17'h17523:	data_out=16'h8a00;
17'h17524:	data_out=16'h8a00;
17'h17525:	data_out=16'h80c;
17'h17526:	data_out=16'h9f5;
17'h17527:	data_out=16'ha00;
17'h17528:	data_out=16'h21d;
17'h17529:	data_out=16'ha00;
17'h1752a:	data_out=16'h9ff;
17'h1752b:	data_out=16'ha00;
17'h1752c:	data_out=16'h9ee;
17'h1752d:	data_out=16'ha00;
17'h1752e:	data_out=16'h9ff;
17'h1752f:	data_out=16'ha00;
17'h17530:	data_out=16'ha00;
17'h17531:	data_out=16'h9be;
17'h17532:	data_out=16'h9df;
17'h17533:	data_out=16'ha00;
17'h17534:	data_out=16'ha00;
17'h17535:	data_out=16'h9e3;
17'h17536:	data_out=16'ha00;
17'h17537:	data_out=16'ha00;
17'h17538:	data_out=16'ha00;
17'h17539:	data_out=16'ha00;
17'h1753a:	data_out=16'h165;
17'h1753b:	data_out=16'h9cf;
17'h1753c:	data_out=16'ha00;
17'h1753d:	data_out=16'h9fe;
17'h1753e:	data_out=16'h224;
17'h1753f:	data_out=16'h9e3;
17'h17540:	data_out=16'h9db;
17'h17541:	data_out=16'ha00;
17'h17542:	data_out=16'ha00;
17'h17543:	data_out=16'h805f;
17'h17544:	data_out=16'h9dc;
17'h17545:	data_out=16'h850;
17'h17546:	data_out=16'ha00;
17'h17547:	data_out=16'h8132;
17'h17548:	data_out=16'ha00;
17'h17549:	data_out=16'h91e;
17'h1754a:	data_out=16'ha00;
17'h1754b:	data_out=16'ha00;
17'h1754c:	data_out=16'h99e;
17'h1754d:	data_out=16'ha00;
17'h1754e:	data_out=16'ha00;
17'h1754f:	data_out=16'hec;
17'h17550:	data_out=16'h9fe;
17'h17551:	data_out=16'h95a;
17'h17552:	data_out=16'h8a00;
17'h17553:	data_out=16'ha00;
17'h17554:	data_out=16'ha00;
17'h17555:	data_out=16'h9f6;
17'h17556:	data_out=16'h9fc;
17'h17557:	data_out=16'h805e;
17'h17558:	data_out=16'ha00;
17'h17559:	data_out=16'h9a7;
17'h1755a:	data_out=16'ha00;
17'h1755b:	data_out=16'h9df;
17'h1755c:	data_out=16'ha00;
17'h1755d:	data_out=16'ha00;
17'h1755e:	data_out=16'ha00;
17'h1755f:	data_out=16'h8b6;
17'h17560:	data_out=16'h9f8;
17'h17561:	data_out=16'h9e2;
17'h17562:	data_out=16'ha00;
17'h17563:	data_out=16'ha00;
17'h17564:	data_out=16'ha00;
17'h17565:	data_out=16'h9c8;
17'h17566:	data_out=16'h5f4;
17'h17567:	data_out=16'h9ff;
17'h17568:	data_out=16'h1c3;
17'h17569:	data_out=16'ha00;
17'h1756a:	data_out=16'h16f;
17'h1756b:	data_out=16'h9ea;
17'h1756c:	data_out=16'h9fe;
17'h1756d:	data_out=16'ha00;
17'h1756e:	data_out=16'h170;
17'h1756f:	data_out=16'h9f4;
17'h17570:	data_out=16'h180;
17'h17571:	data_out=16'h38;
17'h17572:	data_out=16'h9ba;
17'h17573:	data_out=16'h9d5;
17'h17574:	data_out=16'ha00;
17'h17575:	data_out=16'h9e7;
17'h17576:	data_out=16'ha00;
17'h17577:	data_out=16'h9fe;
17'h17578:	data_out=16'h9c0;
17'h17579:	data_out=16'ha00;
17'h1757a:	data_out=16'ha00;
17'h1757b:	data_out=16'h226;
17'h1757c:	data_out=16'h821d;
17'h1757d:	data_out=16'ha5;
17'h1757e:	data_out=16'h9b6;
17'h1757f:	data_out=16'h133;
17'h17580:	data_out=16'h9fc;
17'h17581:	data_out=16'h9fe;
17'h17582:	data_out=16'h9ff;
17'h17583:	data_out=16'h9f9;
17'h17584:	data_out=16'h9f4;
17'h17585:	data_out=16'h9fc;
17'h17586:	data_out=16'h5f1;
17'h17587:	data_out=16'h307;
17'h17588:	data_out=16'ha00;
17'h17589:	data_out=16'h44e;
17'h1758a:	data_out=16'h9eb;
17'h1758b:	data_out=16'ha00;
17'h1758c:	data_out=16'ha00;
17'h1758d:	data_out=16'h9f0;
17'h1758e:	data_out=16'h162;
17'h1758f:	data_out=16'h9fc;
17'h17590:	data_out=16'h9f4;
17'h17591:	data_out=16'h9fb;
17'h17592:	data_out=16'h9ff;
17'h17593:	data_out=16'h9f8;
17'h17594:	data_out=16'ha00;
17'h17595:	data_out=16'h618;
17'h17596:	data_out=16'h9fb;
17'h17597:	data_out=16'ha00;
17'h17598:	data_out=16'h8226;
17'h17599:	data_out=16'h76e;
17'h1759a:	data_out=16'h9fb;
17'h1759b:	data_out=16'ha00;
17'h1759c:	data_out=16'ha00;
17'h1759d:	data_out=16'h9fd;
17'h1759e:	data_out=16'ha00;
17'h1759f:	data_out=16'h8279;
17'h175a0:	data_out=16'h9ff;
17'h175a1:	data_out=16'h179;
17'h175a2:	data_out=16'h9ff;
17'h175a3:	data_out=16'h8a00;
17'h175a4:	data_out=16'h8a00;
17'h175a5:	data_out=16'h8d2;
17'h175a6:	data_out=16'h9f4;
17'h175a7:	data_out=16'h9fe;
17'h175a8:	data_out=16'h1d5;
17'h175a9:	data_out=16'h9fb;
17'h175aa:	data_out=16'h9fa;
17'h175ab:	data_out=16'ha00;
17'h175ac:	data_out=16'h9fa;
17'h175ad:	data_out=16'h9fc;
17'h175ae:	data_out=16'h9fe;
17'h175af:	data_out=16'ha00;
17'h175b0:	data_out=16'ha00;
17'h175b1:	data_out=16'h9fa;
17'h175b2:	data_out=16'h9fb;
17'h175b3:	data_out=16'ha00;
17'h175b4:	data_out=16'h9fe;
17'h175b5:	data_out=16'h9fb;
17'h175b6:	data_out=16'ha00;
17'h175b7:	data_out=16'ha00;
17'h175b8:	data_out=16'ha00;
17'h175b9:	data_out=16'ha00;
17'h175ba:	data_out=16'h80d1;
17'h175bb:	data_out=16'h9fb;
17'h175bc:	data_out=16'ha00;
17'h175bd:	data_out=16'h9fc;
17'h175be:	data_out=16'h1db;
17'h175bf:	data_out=16'h9fb;
17'h175c0:	data_out=16'h9f8;
17'h175c1:	data_out=16'ha00;
17'h175c2:	data_out=16'h9f9;
17'h175c3:	data_out=16'h26d;
17'h175c4:	data_out=16'h9fb;
17'h175c5:	data_out=16'h67e;
17'h175c6:	data_out=16'ha00;
17'h175c7:	data_out=16'h81c5;
17'h175c8:	data_out=16'ha00;
17'h175c9:	data_out=16'h96e;
17'h175ca:	data_out=16'ha00;
17'h175cb:	data_out=16'h9f9;
17'h175cc:	data_out=16'h4f8;
17'h175cd:	data_out=16'ha00;
17'h175ce:	data_out=16'ha00;
17'h175cf:	data_out=16'h8154;
17'h175d0:	data_out=16'h9ff;
17'h175d1:	data_out=16'h9c0;
17'h175d2:	data_out=16'h8a00;
17'h175d3:	data_out=16'ha00;
17'h175d4:	data_out=16'ha00;
17'h175d5:	data_out=16'h9ef;
17'h175d6:	data_out=16'h9fc;
17'h175d7:	data_out=16'h3d8;
17'h175d8:	data_out=16'ha00;
17'h175d9:	data_out=16'h9ed;
17'h175da:	data_out=16'ha00;
17'h175db:	data_out=16'h9fb;
17'h175dc:	data_out=16'ha00;
17'h175dd:	data_out=16'ha00;
17'h175de:	data_out=16'ha00;
17'h175df:	data_out=16'h43a;
17'h175e0:	data_out=16'h9f5;
17'h175e1:	data_out=16'h9fb;
17'h175e2:	data_out=16'h9fb;
17'h175e3:	data_out=16'ha00;
17'h175e4:	data_out=16'h9ff;
17'h175e5:	data_out=16'h9fa;
17'h175e6:	data_out=16'h372;
17'h175e7:	data_out=16'h9fe;
17'h175e8:	data_out=16'h190;
17'h175e9:	data_out=16'ha00;
17'h175ea:	data_out=16'h14d;
17'h175eb:	data_out=16'h9fc;
17'h175ec:	data_out=16'h9f9;
17'h175ed:	data_out=16'ha00;
17'h175ee:	data_out=16'h14e;
17'h175ef:	data_out=16'h9fc;
17'h175f0:	data_out=16'h15a;
17'h175f1:	data_out=16'h82b0;
17'h175f2:	data_out=16'h9f1;
17'h175f3:	data_out=16'h9f8;
17'h175f4:	data_out=16'ha00;
17'h175f5:	data_out=16'h9ff;
17'h175f6:	data_out=16'h5f6;
17'h175f7:	data_out=16'h9f8;
17'h175f8:	data_out=16'h86f;
17'h175f9:	data_out=16'h9ff;
17'h175fa:	data_out=16'ha00;
17'h175fb:	data_out=16'h1dd;
17'h175fc:	data_out=16'h81d8;
17'h175fd:	data_out=16'h428;
17'h175fe:	data_out=16'h961;
17'h175ff:	data_out=16'h2c2;
17'h17600:	data_out=16'h25c;
17'h17601:	data_out=16'h95f;
17'h17602:	data_out=16'h9ff;
17'h17603:	data_out=16'ha00;
17'h17604:	data_out=16'h60d;
17'h17605:	data_out=16'ha00;
17'h17606:	data_out=16'h9e1;
17'h17607:	data_out=16'h84cc;
17'h17608:	data_out=16'ha00;
17'h17609:	data_out=16'h30d;
17'h1760a:	data_out=16'h945;
17'h1760b:	data_out=16'ha00;
17'h1760c:	data_out=16'h973;
17'h1760d:	data_out=16'h670;
17'h1760e:	data_out=16'h260;
17'h1760f:	data_out=16'h907;
17'h17610:	data_out=16'h9fb;
17'h17611:	data_out=16'h9ff;
17'h17612:	data_out=16'h531;
17'h17613:	data_out=16'h9fc;
17'h17614:	data_out=16'ha00;
17'h17615:	data_out=16'h2d5;
17'h17616:	data_out=16'h992;
17'h17617:	data_out=16'ha00;
17'h17618:	data_out=16'h8289;
17'h17619:	data_out=16'h376;
17'h1761a:	data_out=16'h7fa;
17'h1761b:	data_out=16'ha00;
17'h1761c:	data_out=16'ha00;
17'h1761d:	data_out=16'h9fe;
17'h1761e:	data_out=16'ha00;
17'h1761f:	data_out=16'h1dc;
17'h17620:	data_out=16'h7ed;
17'h17621:	data_out=16'h273;
17'h17622:	data_out=16'h994;
17'h17623:	data_out=16'h874c;
17'h17624:	data_out=16'h8749;
17'h17625:	data_out=16'h546;
17'h17626:	data_out=16'h9fa;
17'h17627:	data_out=16'h9ff;
17'h17628:	data_out=16'h2c2;
17'h17629:	data_out=16'h9ea;
17'h1762a:	data_out=16'h341;
17'h1762b:	data_out=16'h804;
17'h1762c:	data_out=16'h874;
17'h1762d:	data_out=16'h9d5;
17'h1762e:	data_out=16'h77a;
17'h1762f:	data_out=16'ha00;
17'h17630:	data_out=16'h9ff;
17'h17631:	data_out=16'h547;
17'h17632:	data_out=16'h9ff;
17'h17633:	data_out=16'ha00;
17'h17634:	data_out=16'h80f4;
17'h17635:	data_out=16'h9fe;
17'h17636:	data_out=16'h965;
17'h17637:	data_out=16'h9ff;
17'h17638:	data_out=16'h8e2;
17'h17639:	data_out=16'ha00;
17'h1763a:	data_out=16'h8a00;
17'h1763b:	data_out=16'h9ff;
17'h1763c:	data_out=16'ha00;
17'h1763d:	data_out=16'h9fc;
17'h1763e:	data_out=16'h2c6;
17'h1763f:	data_out=16'ha00;
17'h17640:	data_out=16'h9fd;
17'h17641:	data_out=16'ha00;
17'h17642:	data_out=16'h9fa;
17'h17643:	data_out=16'h9f7;
17'h17644:	data_out=16'h9ff;
17'h17645:	data_out=16'h326;
17'h17646:	data_out=16'ha00;
17'h17647:	data_out=16'h8954;
17'h17648:	data_out=16'h231;
17'h17649:	data_out=16'h671;
17'h1764a:	data_out=16'h8285;
17'h1764b:	data_out=16'h371;
17'h1764c:	data_out=16'h8852;
17'h1764d:	data_out=16'h97b;
17'h1764e:	data_out=16'h54a;
17'h1764f:	data_out=16'h8a00;
17'h17650:	data_out=16'ha00;
17'h17651:	data_out=16'h9fb;
17'h17652:	data_out=16'h87c4;
17'h17653:	data_out=16'ha00;
17'h17654:	data_out=16'h9fe;
17'h17655:	data_out=16'h9f9;
17'h17656:	data_out=16'ha00;
17'h17657:	data_out=16'h7b1;
17'h17658:	data_out=16'ha00;
17'h17659:	data_out=16'h9f8;
17'h1765a:	data_out=16'ha00;
17'h1765b:	data_out=16'h9ff;
17'h1765c:	data_out=16'ha00;
17'h1765d:	data_out=16'h922;
17'h1765e:	data_out=16'ha00;
17'h1765f:	data_out=16'h852b;
17'h17660:	data_out=16'h8cf;
17'h17661:	data_out=16'h9ff;
17'h17662:	data_out=16'ha00;
17'h17663:	data_out=16'ha00;
17'h17664:	data_out=16'h547;
17'h17665:	data_out=16'ha00;
17'h17666:	data_out=16'h317;
17'h17667:	data_out=16'h38f;
17'h17668:	data_out=16'h28a;
17'h17669:	data_out=16'ha00;
17'h1766a:	data_out=16'h254;
17'h1766b:	data_out=16'h9ff;
17'h1766c:	data_out=16'h10;
17'h1766d:	data_out=16'ha00;
17'h1766e:	data_out=16'h254;
17'h1766f:	data_out=16'ha00;
17'h17670:	data_out=16'h25b;
17'h17671:	data_out=16'h89fe;
17'h17672:	data_out=16'h9fa;
17'h17673:	data_out=16'h9fd;
17'h17674:	data_out=16'ha00;
17'h17675:	data_out=16'ha00;
17'h17676:	data_out=16'h2ca;
17'h17677:	data_out=16'h9f9;
17'h17678:	data_out=16'ha00;
17'h17679:	data_out=16'h45d;
17'h1767a:	data_out=16'ha00;
17'h1767b:	data_out=16'h2c8;
17'h1767c:	data_out=16'h849b;
17'h1767d:	data_out=16'h8f2;
17'h1767e:	data_out=16'h9f3;
17'h1767f:	data_out=16'h81d7;
17'h17680:	data_out=16'h8118;
17'h17681:	data_out=16'hd6;
17'h17682:	data_out=16'h69b;
17'h17683:	data_out=16'h83c;
17'h17684:	data_out=16'h89b2;
17'h17685:	data_out=16'h80de;
17'h17686:	data_out=16'h68;
17'h17687:	data_out=16'h89af;
17'h17688:	data_out=16'h9b7;
17'h17689:	data_out=16'h1f5;
17'h1768a:	data_out=16'h831e;
17'h1768b:	data_out=16'ha00;
17'h1768c:	data_out=16'h856d;
17'h1768d:	data_out=16'h38e;
17'h1768e:	data_out=16'h80b3;
17'h1768f:	data_out=16'h3d5;
17'h17690:	data_out=16'h7aa;
17'h17691:	data_out=16'h883c;
17'h17692:	data_out=16'h525;
17'h17693:	data_out=16'h75d;
17'h17694:	data_out=16'ha00;
17'h17695:	data_out=16'h81d3;
17'h17696:	data_out=16'h8088;
17'h17697:	data_out=16'ha00;
17'h17698:	data_out=16'h812d;
17'h17699:	data_out=16'h80e1;
17'h1769a:	data_out=16'h8895;
17'h1769b:	data_out=16'ha00;
17'h1769c:	data_out=16'h803c;
17'h1769d:	data_out=16'h6d;
17'h1769e:	data_out=16'h82d;
17'h1769f:	data_out=16'h86a0;
17'h176a0:	data_out=16'h185;
17'h176a1:	data_out=16'h80a4;
17'h176a2:	data_out=16'h5a4;
17'h176a3:	data_out=16'h854a;
17'h176a4:	data_out=16'h8548;
17'h176a5:	data_out=16'h27a;
17'h176a6:	data_out=16'h8ce;
17'h176a7:	data_out=16'h1df;
17'h176a8:	data_out=16'h8058;
17'h176a9:	data_out=16'h839;
17'h176aa:	data_out=16'h1b8;
17'h176ab:	data_out=16'h22e;
17'h176ac:	data_out=16'h810e;
17'h176ad:	data_out=16'h9fe;
17'h176ae:	data_out=16'h6de;
17'h176af:	data_out=16'h9ff;
17'h176b0:	data_out=16'h86f8;
17'h176b1:	data_out=16'h8789;
17'h176b2:	data_out=16'h8733;
17'h176b3:	data_out=16'h8ca;
17'h176b4:	data_out=16'h8932;
17'h176b5:	data_out=16'h83e9;
17'h176b6:	data_out=16'h6e1;
17'h176b7:	data_out=16'h6fc;
17'h176b8:	data_out=16'h858b;
17'h176b9:	data_out=16'h82a;
17'h176ba:	data_out=16'h8775;
17'h176bb:	data_out=16'h8558;
17'h176bc:	data_out=16'ha00;
17'h176bd:	data_out=16'h82de;
17'h176be:	data_out=16'h803c;
17'h176bf:	data_out=16'h80e9;
17'h176c0:	data_out=16'h809a;
17'h176c1:	data_out=16'ha00;
17'h176c2:	data_out=16'h1c6;
17'h176c3:	data_out=16'h1b8;
17'h176c4:	data_out=16'h82b5;
17'h176c5:	data_out=16'h81cc;
17'h176c6:	data_out=16'ha00;
17'h176c7:	data_out=16'h888d;
17'h176c8:	data_out=16'h359;
17'h176c9:	data_out=16'h2b5;
17'h176ca:	data_out=16'h8970;
17'h176cb:	data_out=16'h8507;
17'h176cc:	data_out=16'h873e;
17'h176cd:	data_out=16'h5bf;
17'h176ce:	data_out=16'h1de;
17'h176cf:	data_out=16'h88e8;
17'h176d0:	data_out=16'h91;
17'h176d1:	data_out=16'h43d;
17'h176d2:	data_out=16'h8557;
17'h176d3:	data_out=16'h7f5;
17'h176d4:	data_out=16'h7b6;
17'h176d5:	data_out=16'h9f6;
17'h176d6:	data_out=16'h4df;
17'h176d7:	data_out=16'h497;
17'h176d8:	data_out=16'ha00;
17'h176d9:	data_out=16'h800b;
17'h176da:	data_out=16'ha00;
17'h176db:	data_out=16'h8581;
17'h176dc:	data_out=16'h99;
17'h176dd:	data_out=16'h334;
17'h176de:	data_out=16'h9ff;
17'h176df:	data_out=16'h8184;
17'h176e0:	data_out=16'h2c1;
17'h176e1:	data_out=16'h8563;
17'h176e2:	data_out=16'h9ff;
17'h176e3:	data_out=16'h945;
17'h176e4:	data_out=16'h85e8;
17'h176e5:	data_out=16'hb;
17'h176e6:	data_out=16'h8139;
17'h176e7:	data_out=16'h2b5;
17'h176e8:	data_out=16'h808d;
17'h176e9:	data_out=16'h9f1;
17'h176ea:	data_out=16'h80b9;
17'h176eb:	data_out=16'h86cc;
17'h176ec:	data_out=16'h8159;
17'h176ed:	data_out=16'h91f;
17'h176ee:	data_out=16'h80b9;
17'h176ef:	data_out=16'h3d2;
17'h176f0:	data_out=16'h80b5;
17'h176f1:	data_out=16'h8a00;
17'h176f2:	data_out=16'h85aa;
17'h176f3:	data_out=16'h8438;
17'h176f4:	data_out=16'h8703;
17'h176f5:	data_out=16'h9fb;
17'h176f6:	data_out=16'h80c7;
17'h176f7:	data_out=16'h620;
17'h176f8:	data_out=16'h1f5;
17'h176f9:	data_out=16'h29d;
17'h176fa:	data_out=16'ha00;
17'h176fb:	data_out=16'h8038;
17'h176fc:	data_out=16'h8241;
17'h176fd:	data_out=16'h8230;
17'h176fe:	data_out=16'h9f7;
17'h176ff:	data_out=16'h8962;
17'h17700:	data_out=16'h803a;
17'h17701:	data_out=16'hd;
17'h17702:	data_out=16'h34f;
17'h17703:	data_out=16'h2cf;
17'h17704:	data_out=16'h8a00;
17'h17705:	data_out=16'h85bb;
17'h17706:	data_out=16'h82c8;
17'h17707:	data_out=16'h875c;
17'h17708:	data_out=16'h480;
17'h17709:	data_out=16'h117;
17'h1770a:	data_out=16'h84df;
17'h1770b:	data_out=16'h6ee;
17'h1770c:	data_out=16'h873b;
17'h1770d:	data_out=16'h1ea;
17'h1770e:	data_out=16'h80ad;
17'h1770f:	data_out=16'h214;
17'h17710:	data_out=16'h505;
17'h17711:	data_out=16'h8a00;
17'h17712:	data_out=16'h46a;
17'h17713:	data_out=16'h24b;
17'h17714:	data_out=16'h638;
17'h17715:	data_out=16'h8263;
17'h17716:	data_out=16'h829c;
17'h17717:	data_out=16'h814;
17'h17718:	data_out=16'h810a;
17'h17719:	data_out=16'h830e;
17'h1771a:	data_out=16'h8972;
17'h1771b:	data_out=16'ha00;
17'h1771c:	data_out=16'h83c0;
17'h1771d:	data_out=16'h81ed;
17'h1771e:	data_out=16'h550;
17'h1771f:	data_out=16'h8589;
17'h17720:	data_out=16'h149;
17'h17721:	data_out=16'h809e;
17'h17722:	data_out=16'h318;
17'h17723:	data_out=16'h8368;
17'h17724:	data_out=16'h8367;
17'h17725:	data_out=16'h12;
17'h17726:	data_out=16'h429;
17'h17727:	data_out=16'h80ec;
17'h17728:	data_out=16'h808d;
17'h17729:	data_out=16'h53d;
17'h1772a:	data_out=16'h2a9;
17'h1772b:	data_out=16'h8087;
17'h1772c:	data_out=16'h82ed;
17'h1772d:	data_out=16'h768;
17'h1772e:	data_out=16'h6fd;
17'h1772f:	data_out=16'h662;
17'h17730:	data_out=16'h894f;
17'h17731:	data_out=16'h88df;
17'h17732:	data_out=16'h894d;
17'h17733:	data_out=16'h554;
17'h17734:	data_out=16'h870b;
17'h17735:	data_out=16'h8873;
17'h17736:	data_out=16'h58b;
17'h17737:	data_out=16'h35f;
17'h17738:	data_out=16'h8607;
17'h17739:	data_out=16'h551;
17'h1773a:	data_out=16'h81b0;
17'h1773b:	data_out=16'h8821;
17'h1773c:	data_out=16'h92d;
17'h1773d:	data_out=16'h83fb;
17'h1773e:	data_out=16'h8087;
17'h1773f:	data_out=16'h85ca;
17'h17740:	data_out=16'h8304;
17'h17741:	data_out=16'h787;
17'h17742:	data_out=16'h74;
17'h17743:	data_out=16'h819b;
17'h17744:	data_out=16'h86a9;
17'h17745:	data_out=16'h826d;
17'h17746:	data_out=16'h65d;
17'h17747:	data_out=16'h831d;
17'h17748:	data_out=16'h41e;
17'h17749:	data_out=16'h8054;
17'h1774a:	data_out=16'h86e0;
17'h1774b:	data_out=16'h8401;
17'h1774c:	data_out=16'h8377;
17'h1774d:	data_out=16'h33e;
17'h1774e:	data_out=16'h295;
17'h1774f:	data_out=16'h84a4;
17'h17750:	data_out=16'h8170;
17'h17751:	data_out=16'h81f3;
17'h17752:	data_out=16'h83a4;
17'h17753:	data_out=16'h3e6;
17'h17754:	data_out=16'h4c8;
17'h17755:	data_out=16'h865;
17'h17756:	data_out=16'h158;
17'h17757:	data_out=16'h187;
17'h17758:	data_out=16'h786;
17'h17759:	data_out=16'h82f8;
17'h1775a:	data_out=16'ha00;
17'h1775b:	data_out=16'h88c4;
17'h1775c:	data_out=16'h8316;
17'h1775d:	data_out=16'h2d2;
17'h1775e:	data_out=16'h6e5;
17'h1775f:	data_out=16'had;
17'h17760:	data_out=16'h1f;
17'h17761:	data_out=16'h88a7;
17'h17762:	data_out=16'h6cd;
17'h17763:	data_out=16'h589;
17'h17764:	data_out=16'h862a;
17'h17765:	data_out=16'h855a;
17'h17766:	data_out=16'h83c7;
17'h17767:	data_out=16'h29e;
17'h17768:	data_out=16'h809a;
17'h17769:	data_out=16'h51b;
17'h1776a:	data_out=16'h80bf;
17'h1776b:	data_out=16'h88b0;
17'h1776c:	data_out=16'h15b;
17'h1776d:	data_out=16'h57d;
17'h1776e:	data_out=16'h80a6;
17'h1776f:	data_out=16'h82c7;
17'h17770:	data_out=16'h80b3;
17'h17771:	data_out=16'h83cf;
17'h17772:	data_out=16'h8764;
17'h17773:	data_out=16'h8746;
17'h17774:	data_out=16'h8955;
17'h17775:	data_out=16'h806c;
17'h17776:	data_out=16'h81d9;
17'h17777:	data_out=16'hbb;
17'h17778:	data_out=16'h829b;
17'h17779:	data_out=16'h492;
17'h1777a:	data_out=16'h609;
17'h1777b:	data_out=16'h8088;
17'h1777c:	data_out=16'h809a;
17'h1777d:	data_out=16'h84e8;
17'h1777e:	data_out=16'h4ad;
17'h1777f:	data_out=16'h8741;
17'h17780:	data_out=16'h81bc;
17'h17781:	data_out=16'h818f;
17'h17782:	data_out=16'h122;
17'h17783:	data_out=16'h9b;
17'h17784:	data_out=16'h8110;
17'h17785:	data_out=16'h8047;
17'h17786:	data_out=16'h28;
17'h17787:	data_out=16'h80c5;
17'h17788:	data_out=16'h802b;
17'h17789:	data_out=16'h2;
17'h1778a:	data_out=16'h81a0;
17'h1778b:	data_out=16'h801f;
17'h1778c:	data_out=16'h814e;
17'h1778d:	data_out=16'h80a0;
17'h1778e:	data_out=16'h31;
17'h1778f:	data_out=16'h806d;
17'h17790:	data_out=16'h6c;
17'h17791:	data_out=16'h81cc;
17'h17792:	data_out=16'hdd;
17'h17793:	data_out=16'h8007;
17'h17794:	data_out=16'h1ae;
17'h17795:	data_out=16'h8105;
17'h17796:	data_out=16'h80f1;
17'h17797:	data_out=16'h1da;
17'h17798:	data_out=16'h80bd;
17'h17799:	data_out=16'h8132;
17'h1779a:	data_out=16'h818f;
17'h1779b:	data_out=16'h8045;
17'h1779c:	data_out=16'ha1;
17'h1779d:	data_out=16'h8056;
17'h1779e:	data_out=16'h11f;
17'h1779f:	data_out=16'h66;
17'h177a0:	data_out=16'h80ca;
17'h177a1:	data_out=16'h34;
17'h177a2:	data_out=16'hd3;
17'h177a3:	data_out=16'h8159;
17'h177a4:	data_out=16'h8159;
17'h177a5:	data_out=16'h800c;
17'h177a6:	data_out=16'heb;
17'h177a7:	data_out=16'h804d;
17'h177a8:	data_out=16'h3a;
17'h177a9:	data_out=16'h8001;
17'h177aa:	data_out=16'h801b;
17'h177ab:	data_out=16'h8137;
17'h177ac:	data_out=16'h8078;
17'h177ad:	data_out=16'h6a;
17'h177ae:	data_out=16'h14f;
17'h177af:	data_out=16'h8082;
17'h177b0:	data_out=16'h8197;
17'h177b1:	data_out=16'h82e0;
17'h177b2:	data_out=16'h8197;
17'h177b3:	data_out=16'h181;
17'h177b4:	data_out=16'h8243;
17'h177b5:	data_out=16'h81c7;
17'h177b6:	data_out=16'h8098;
17'h177b7:	data_out=16'h12f;
17'h177b8:	data_out=16'h8184;
17'h177b9:	data_out=16'hd0;
17'h177ba:	data_out=16'h4d;
17'h177bb:	data_out=16'h81e7;
17'h177bc:	data_out=16'h1b5;
17'h177bd:	data_out=16'h8091;
17'h177be:	data_out=16'h31;
17'h177bf:	data_out=16'h80dc;
17'h177c0:	data_out=16'h8d;
17'h177c1:	data_out=16'h18f;
17'h177c2:	data_out=16'h814e;
17'h177c3:	data_out=16'h116;
17'h177c4:	data_out=16'h811d;
17'h177c5:	data_out=16'h80c7;
17'h177c6:	data_out=16'h196;
17'h177c7:	data_out=16'h8076;
17'h177c8:	data_out=16'hc0;
17'h177c9:	data_out=16'h2;
17'h177ca:	data_out=16'h81e5;
17'h177cb:	data_out=16'h8263;
17'h177cc:	data_out=16'h81a3;
17'h177cd:	data_out=16'h9b;
17'h177ce:	data_out=16'h80b5;
17'h177cf:	data_out=16'h81e0;
17'h177d0:	data_out=16'ha4;
17'h177d1:	data_out=16'h8009;
17'h177d2:	data_out=16'h815a;
17'h177d3:	data_out=16'h8041;
17'h177d4:	data_out=16'h8122;
17'h177d5:	data_out=16'h22c;
17'h177d6:	data_out=16'h179;
17'h177d7:	data_out=16'h199;
17'h177d8:	data_out=16'h220;
17'h177d9:	data_out=16'h12c;
17'h177da:	data_out=16'h16d;
17'h177db:	data_out=16'h818c;
17'h177dc:	data_out=16'h8164;
17'h177dd:	data_out=16'h8066;
17'h177de:	data_out=16'h80ae;
17'h177df:	data_out=16'h80bb;
17'h177e0:	data_out=16'h8085;
17'h177e1:	data_out=16'h81a5;
17'h177e2:	data_out=16'hed;
17'h177e3:	data_out=16'h173;
17'h177e4:	data_out=16'h814c;
17'h177e5:	data_out=16'h8125;
17'h177e6:	data_out=16'h813b;
17'h177e7:	data_out=16'hc5;
17'h177e8:	data_out=16'h38;
17'h177e9:	data_out=16'h47;
17'h177ea:	data_out=16'h2b;
17'h177eb:	data_out=16'h816c;
17'h177ec:	data_out=16'h80fc;
17'h177ed:	data_out=16'h17c;
17'h177ee:	data_out=16'h3e;
17'h177ef:	data_out=16'h39;
17'h177f0:	data_out=16'h32;
17'h177f1:	data_out=16'h804c;
17'h177f2:	data_out=16'h8038;
17'h177f3:	data_out=16'h8118;
17'h177f4:	data_out=16'h819e;
17'h177f5:	data_out=16'h91;
17'h177f6:	data_out=16'h810d;
17'h177f7:	data_out=16'h7e;
17'h177f8:	data_out=16'h26;
17'h177f9:	data_out=16'h5e;
17'h177fa:	data_out=16'h194;
17'h177fb:	data_out=16'h40;
17'h177fc:	data_out=16'h807f;
17'h177fd:	data_out=16'h8065;
17'h177fe:	data_out=16'he0;
17'h177ff:	data_out=16'h80a3;
17'h17800:	data_out=16'h8029;
17'h17801:	data_out=16'h802b;
17'h17802:	data_out=16'h14;
17'h17803:	data_out=16'h10;
17'h17804:	data_out=16'h8021;
17'h17805:	data_out=16'h802c;
17'h17806:	data_out=16'h8021;
17'h17807:	data_out=16'h8012;
17'h17808:	data_out=16'h800e;
17'h17809:	data_out=16'h8012;
17'h1780a:	data_out=16'h8031;
17'h1780b:	data_out=16'hb;
17'h1780c:	data_out=16'h8024;
17'h1780d:	data_out=16'h8019;
17'h1780e:	data_out=16'h8006;
17'h1780f:	data_out=16'h8020;
17'h17810:	data_out=16'h1b;
17'h17811:	data_out=16'h8028;
17'h17812:	data_out=16'h800b;
17'h17813:	data_out=16'h800e;
17'h17814:	data_out=16'h8001;
17'h17815:	data_out=16'h8025;
17'h17816:	data_out=16'h801d;
17'h17817:	data_out=16'h4;
17'h17818:	data_out=16'h8015;
17'h17819:	data_out=16'h8017;
17'h1781a:	data_out=16'h8032;
17'h1781b:	data_out=16'h8005;
17'h1781c:	data_out=16'h8019;
17'h1781d:	data_out=16'h801f;
17'h1781e:	data_out=16'h800c;
17'h1781f:	data_out=16'h800d;
17'h17820:	data_out=16'h8034;
17'h17821:	data_out=16'h8000;
17'h17822:	data_out=16'h8009;
17'h17823:	data_out=16'h8027;
17'h17824:	data_out=16'h801e;
17'h17825:	data_out=16'h800c;
17'h17826:	data_out=16'hd;
17'h17827:	data_out=16'h8014;
17'h17828:	data_out=16'h8008;
17'h17829:	data_out=16'h8000;
17'h1782a:	data_out=16'h8017;
17'h1782b:	data_out=16'h801a;
17'h1782c:	data_out=16'h801b;
17'h1782d:	data_out=16'h4;
17'h1782e:	data_out=16'h16;
17'h1782f:	data_out=16'h8019;
17'h17830:	data_out=16'h8030;
17'h17831:	data_out=16'h8040;
17'h17832:	data_out=16'h802f;
17'h17833:	data_out=16'h8013;
17'h17834:	data_out=16'h802b;
17'h17835:	data_out=16'h8036;
17'h17836:	data_out=16'h800b;
17'h17837:	data_out=16'h8;
17'h17838:	data_out=16'h803d;
17'h17839:	data_out=16'h8003;
17'h1783a:	data_out=16'h8015;
17'h1783b:	data_out=16'h803f;
17'h1783c:	data_out=16'h2a;
17'h1783d:	data_out=16'h8015;
17'h1783e:	data_out=16'h8007;
17'h1783f:	data_out=16'h8028;
17'h17840:	data_out=16'h8032;
17'h17841:	data_out=16'h6;
17'h17842:	data_out=16'h8004;
17'h17843:	data_out=16'h10;
17'h17844:	data_out=16'h8022;
17'h17845:	data_out=16'h8007;
17'h17846:	data_out=16'h27;
17'h17847:	data_out=16'h8026;
17'h17848:	data_out=16'h800e;
17'h17849:	data_out=16'h8008;
17'h1784a:	data_out=16'h8035;
17'h1784b:	data_out=16'h8024;
17'h1784c:	data_out=16'h8027;
17'h1784d:	data_out=16'h800a;
17'h1784e:	data_out=16'h8035;
17'h1784f:	data_out=16'h8025;
17'h17850:	data_out=16'h8012;
17'h17851:	data_out=16'h8001;
17'h17852:	data_out=16'h8029;
17'h17853:	data_out=16'h802f;
17'h17854:	data_out=16'h8028;
17'h17855:	data_out=16'h1f;
17'h17856:	data_out=16'h8013;
17'h17857:	data_out=16'h1f;
17'h17858:	data_out=16'h33;
17'h17859:	data_out=16'h800e;
17'h1785a:	data_out=16'h2f;
17'h1785b:	data_out=16'h8030;
17'h1785c:	data_out=16'h8028;
17'h1785d:	data_out=16'h8018;
17'h1785e:	data_out=16'h801d;
17'h1785f:	data_out=16'h8004;
17'h17860:	data_out=16'h800a;
17'h17861:	data_out=16'h8035;
17'h17862:	data_out=16'h5;
17'h17863:	data_out=16'h800a;
17'h17864:	data_out=16'h801e;
17'h17865:	data_out=16'h8029;
17'h17866:	data_out=16'h8020;
17'h17867:	data_out=16'ha;
17'h17868:	data_out=16'h1;
17'h17869:	data_out=16'h9;
17'h1786a:	data_out=16'h800d;
17'h1786b:	data_out=16'h8031;
17'h1786c:	data_out=16'h801c;
17'h1786d:	data_out=16'h8015;
17'h1786e:	data_out=16'h0;
17'h1786f:	data_out=16'h8025;
17'h17870:	data_out=16'h800a;
17'h17871:	data_out=16'h8012;
17'h17872:	data_out=16'h8014;
17'h17873:	data_out=16'h8027;
17'h17874:	data_out=16'h802e;
17'h17875:	data_out=16'h8023;
17'h17876:	data_out=16'h801e;
17'h17877:	data_out=16'h800d;
17'h17878:	data_out=16'h8015;
17'h17879:	data_out=16'h800b;
17'h1787a:	data_out=16'h800e;
17'h1787b:	data_out=16'h8002;
17'h1787c:	data_out=16'h8008;
17'h1787d:	data_out=16'h802d;
17'h1787e:	data_out=16'h10;
17'h1787f:	data_out=16'h801f;
17'h17880:	data_out=16'h6;
17'h17881:	data_out=16'h9;
17'h17882:	data_out=16'h8;
17'h17883:	data_out=16'h12;
17'h17884:	data_out=16'h12;
17'h17885:	data_out=16'h12;
17'h17886:	data_out=16'h8;
17'h17887:	data_out=16'hd;
17'h17888:	data_out=16'h4;
17'h17889:	data_out=16'hb;
17'h1788a:	data_out=16'ha;
17'h1788b:	data_out=16'h4;
17'h1788c:	data_out=16'h13;
17'h1788d:	data_out=16'h4;
17'h1788e:	data_out=16'h8003;
17'h1788f:	data_out=16'h10;
17'h17890:	data_out=16'h8001;
17'h17891:	data_out=16'h7;
17'h17892:	data_out=16'hb;
17'h17893:	data_out=16'h10;
17'h17894:	data_out=16'h5;
17'h17895:	data_out=16'hc;
17'h17896:	data_out=16'h2;
17'h17897:	data_out=16'hb;
17'h17898:	data_out=16'h8002;
17'h17899:	data_out=16'h2;
17'h1789a:	data_out=16'hb;
17'h1789b:	data_out=16'h7;
17'h1789c:	data_out=16'h15;
17'h1789d:	data_out=16'h11;
17'h1789e:	data_out=16'h1;
17'h1789f:	data_out=16'h6;
17'h178a0:	data_out=16'ha;
17'h178a1:	data_out=16'h7;
17'h178a2:	data_out=16'h4;
17'h178a3:	data_out=16'h1;
17'h178a4:	data_out=16'h7;
17'h178a5:	data_out=16'h12;
17'h178a6:	data_out=16'hf;
17'h178a7:	data_out=16'h11;
17'h178a8:	data_out=16'h2;
17'h178a9:	data_out=16'h7;
17'h178aa:	data_out=16'h2;
17'h178ab:	data_out=16'h4;
17'h178ac:	data_out=16'hc;
17'h178ad:	data_out=16'h3;
17'h178ae:	data_out=16'h2;
17'h178af:	data_out=16'he;
17'h178b0:	data_out=16'hd;
17'h178b1:	data_out=16'ha;
17'h178b2:	data_out=16'hf;
17'h178b3:	data_out=16'hf;
17'h178b4:	data_out=16'h9;
17'h178b5:	data_out=16'h13;
17'h178b6:	data_out=16'h12;
17'h178b7:	data_out=16'h9;
17'h178b8:	data_out=16'h10;
17'h178b9:	data_out=16'h3;
17'h178ba:	data_out=16'h12;
17'h178bb:	data_out=16'h12;
17'h178bc:	data_out=16'h8001;
17'h178bd:	data_out=16'h3;
17'h178be:	data_out=16'h8001;
17'h178bf:	data_out=16'hb;
17'h178c0:	data_out=16'h12;
17'h178c1:	data_out=16'ha;
17'h178c2:	data_out=16'he;
17'h178c3:	data_out=16'h3;
17'h178c4:	data_out=16'h7;
17'h178c5:	data_out=16'h7;
17'h178c6:	data_out=16'h8001;
17'h178c7:	data_out=16'h12;
17'h178c8:	data_out=16'hf;
17'h178c9:	data_out=16'h4;
17'h178ca:	data_out=16'h6;
17'h178cb:	data_out=16'h12;
17'h178cc:	data_out=16'hb;
17'h178cd:	data_out=16'h3;
17'h178ce:	data_out=16'hd;
17'h178cf:	data_out=16'h14;
17'h178d0:	data_out=16'h12;
17'h178d1:	data_out=16'he;
17'h178d2:	data_out=16'ha;
17'h178d3:	data_out=16'h7;
17'h178d4:	data_out=16'hd;
17'h178d5:	data_out=16'h8;
17'h178d6:	data_out=16'hd;
17'h178d7:	data_out=16'h8;
17'h178d8:	data_out=16'hc;
17'h178d9:	data_out=16'hd;
17'h178da:	data_out=16'h3;
17'h178db:	data_out=16'h12;
17'h178dc:	data_out=16'hf;
17'h178dd:	data_out=16'hd;
17'h178de:	data_out=16'ha;
17'h178df:	data_out=16'h7;
17'h178e0:	data_out=16'h7;
17'h178e1:	data_out=16'h4;
17'h178e2:	data_out=16'hf;
17'h178e3:	data_out=16'h9;
17'h178e4:	data_out=16'he;
17'h178e5:	data_out=16'h2;
17'h178e6:	data_out=16'h8;
17'h178e7:	data_out=16'hd;
17'h178e8:	data_out=16'h8004;
17'h178e9:	data_out=16'h9;
17'h178ea:	data_out=16'h8000;
17'h178eb:	data_out=16'hb;
17'h178ec:	data_out=16'h9;
17'h178ed:	data_out=16'h9;
17'h178ee:	data_out=16'h8002;
17'h178ef:	data_out=16'hd;
17'h178f0:	data_out=16'h5;
17'h178f1:	data_out=16'h8002;
17'h178f2:	data_out=16'hd;
17'h178f3:	data_out=16'h6;
17'h178f4:	data_out=16'h10;
17'h178f5:	data_out=16'hb;
17'h178f6:	data_out=16'h11;
17'h178f7:	data_out=16'he;
17'h178f8:	data_out=16'h5;
17'h178f9:	data_out=16'h6;
17'h178fa:	data_out=16'h6;
17'h178fb:	data_out=16'h8003;
17'h178fc:	data_out=16'hd;
17'h178fd:	data_out=16'h10;
17'h178fe:	data_out=16'he;
17'h178ff:	data_out=16'h6;
17'h17900:	data_out=16'h8007;
17'h17901:	data_out=16'h2;
17'h17902:	data_out=16'h7;
17'h17903:	data_out=16'h6;
17'h17904:	data_out=16'h2;
17'h17905:	data_out=16'h8002;
17'h17906:	data_out=16'h1;
17'h17907:	data_out=16'h5;
17'h17908:	data_out=16'h7;
17'h17909:	data_out=16'h7;
17'h1790a:	data_out=16'h8006;
17'h1790b:	data_out=16'h2;
17'h1790c:	data_out=16'h1;
17'h1790d:	data_out=16'h8002;
17'h1790e:	data_out=16'h8007;
17'h1790f:	data_out=16'h8007;
17'h17910:	data_out=16'h8001;
17'h17911:	data_out=16'h8;
17'h17912:	data_out=16'h8002;
17'h17913:	data_out=16'h8008;
17'h17914:	data_out=16'h1;
17'h17915:	data_out=16'h8006;
17'h17916:	data_out=16'h2;
17'h17917:	data_out=16'h8;
17'h17918:	data_out=16'h8001;
17'h17919:	data_out=16'h8006;
17'h1791a:	data_out=16'h8007;
17'h1791b:	data_out=16'h8001;
17'h1791c:	data_out=16'h8006;
17'h1791d:	data_out=16'h6;
17'h1791e:	data_out=16'h3;
17'h1791f:	data_out=16'h8004;
17'h17920:	data_out=16'h8001;
17'h17921:	data_out=16'h1;
17'h17922:	data_out=16'h8006;
17'h17923:	data_out=16'h8008;
17'h17924:	data_out=16'h8;
17'h17925:	data_out=16'h4;
17'h17926:	data_out=16'h5;
17'h17927:	data_out=16'h6;
17'h17928:	data_out=16'h1;
17'h17929:	data_out=16'h9;
17'h1792a:	data_out=16'h8001;
17'h1792b:	data_out=16'h8008;
17'h1792c:	data_out=16'h8002;
17'h1792d:	data_out=16'h2;
17'h1792e:	data_out=16'h8005;
17'h1792f:	data_out=16'h6;
17'h17930:	data_out=16'h1;
17'h17931:	data_out=16'h1;
17'h17932:	data_out=16'h7;
17'h17933:	data_out=16'h8007;
17'h17934:	data_out=16'h5;
17'h17935:	data_out=16'h1;
17'h17936:	data_out=16'h8008;
17'h17937:	data_out=16'h8006;
17'h17938:	data_out=16'h4;
17'h17939:	data_out=16'h8006;
17'h1793a:	data_out=16'h3;
17'h1793b:	data_out=16'h7;
17'h1793c:	data_out=16'h8;
17'h1793d:	data_out=16'h8003;
17'h1793e:	data_out=16'h8006;
17'h1793f:	data_out=16'h8002;
17'h17940:	data_out=16'h7;
17'h17941:	data_out=16'h8003;
17'h17942:	data_out=16'h8001;
17'h17943:	data_out=16'h6;
17'h17944:	data_out=16'h8009;
17'h17945:	data_out=16'h8005;
17'h17946:	data_out=16'h3;
17'h17947:	data_out=16'h2;
17'h17948:	data_out=16'h8005;
17'h17949:	data_out=16'h8007;
17'h1794a:	data_out=16'h3;
17'h1794b:	data_out=16'h2;
17'h1794c:	data_out=16'h4;
17'h1794d:	data_out=16'h7;
17'h1794e:	data_out=16'h8001;
17'h1794f:	data_out=16'h8004;
17'h17950:	data_out=16'h8001;
17'h17951:	data_out=16'h8003;
17'h17952:	data_out=16'h8002;
17'h17953:	data_out=16'h8005;
17'h17954:	data_out=16'h6;
17'h17955:	data_out=16'h8001;
17'h17956:	data_out=16'h8002;
17'h17957:	data_out=16'h1;
17'h17958:	data_out=16'h2;
17'h17959:	data_out=16'h8008;
17'h1795a:	data_out=16'h8001;
17'h1795b:	data_out=16'h1;
17'h1795c:	data_out=16'h8002;
17'h1795d:	data_out=16'h2;
17'h1795e:	data_out=16'h8;
17'h1795f:	data_out=16'h8004;
17'h17960:	data_out=16'h8;
17'h17961:	data_out=16'h8002;
17'h17962:	data_out=16'h8008;
17'h17963:	data_out=16'h9;
17'h17964:	data_out=16'h2;
17'h17965:	data_out=16'h4;
17'h17966:	data_out=16'h1;
17'h17967:	data_out=16'h6;
17'h17968:	data_out=16'h6;
17'h17969:	data_out=16'h8005;
17'h1796a:	data_out=16'h8002;
17'h1796b:	data_out=16'h1;
17'h1796c:	data_out=16'h8007;
17'h1796d:	data_out=16'h6;
17'h1796e:	data_out=16'h6;
17'h1796f:	data_out=16'h2;
17'h17970:	data_out=16'h8006;
17'h17971:	data_out=16'h8006;
17'h17972:	data_out=16'h6;
17'h17973:	data_out=16'h8009;
17'h17974:	data_out=16'h2;
17'h17975:	data_out=16'h8005;
17'h17976:	data_out=16'h1;
17'h17977:	data_out=16'h8005;
17'h17978:	data_out=16'h8004;
17'h17979:	data_out=16'h9;
17'h1797a:	data_out=16'h5;
17'h1797b:	data_out=16'h3;
17'h1797c:	data_out=16'h2;
17'h1797d:	data_out=16'h3;
17'h1797e:	data_out=16'h8;
17'h1797f:	data_out=16'h1;
17'h17980:	data_out=16'h8008;
17'h17981:	data_out=16'h9;
17'h17982:	data_out=16'h0;
17'h17983:	data_out=16'h3;
17'h17984:	data_out=16'h4;
17'h17985:	data_out=16'h8007;
17'h17986:	data_out=16'h8001;
17'h17987:	data_out=16'h1;
17'h17988:	data_out=16'h8003;
17'h17989:	data_out=16'h7;
17'h1798a:	data_out=16'h8008;
17'h1798b:	data_out=16'h8000;
17'h1798c:	data_out=16'h4;
17'h1798d:	data_out=16'h7;
17'h1798e:	data_out=16'h8008;
17'h1798f:	data_out=16'h6;
17'h17990:	data_out=16'h8008;
17'h17991:	data_out=16'h7;
17'h17992:	data_out=16'h6;
17'h17993:	data_out=16'h4;
17'h17994:	data_out=16'h8006;
17'h17995:	data_out=16'h8002;
17'h17996:	data_out=16'h8;
17'h17997:	data_out=16'h8001;
17'h17998:	data_out=16'h8002;
17'h17999:	data_out=16'h3;
17'h1799a:	data_out=16'h8007;
17'h1799b:	data_out=16'h9;
17'h1799c:	data_out=16'h8003;
17'h1799d:	data_out=16'h8009;
17'h1799e:	data_out=16'h0;
17'h1799f:	data_out=16'h8002;
17'h179a0:	data_out=16'h8009;
17'h179a1:	data_out=16'h8008;
17'h179a2:	data_out=16'h8008;
17'h179a3:	data_out=16'h4;
17'h179a4:	data_out=16'h8007;
17'h179a5:	data_out=16'h0;
17'h179a6:	data_out=16'h8004;
17'h179a7:	data_out=16'h8001;
17'h179a8:	data_out=16'h8002;
17'h179a9:	data_out=16'h8002;
17'h179aa:	data_out=16'h8;
17'h179ab:	data_out=16'h8008;
17'h179ac:	data_out=16'h8004;
17'h179ad:	data_out=16'h8009;
17'h179ae:	data_out=16'h8;
17'h179af:	data_out=16'h8003;
17'h179b0:	data_out=16'h8;
17'h179b1:	data_out=16'h5;
17'h179b2:	data_out=16'h8008;
17'h179b3:	data_out=16'h8008;
17'h179b4:	data_out=16'h8006;
17'h179b5:	data_out=16'h9;
17'h179b6:	data_out=16'h0;
17'h179b7:	data_out=16'h1;
17'h179b8:	data_out=16'h3;
17'h179b9:	data_out=16'h2;
17'h179ba:	data_out=16'h1;
17'h179bb:	data_out=16'h8009;
17'h179bc:	data_out=16'h3;
17'h179bd:	data_out=16'h8008;
17'h179be:	data_out=16'h8001;
17'h179bf:	data_out=16'h3;
17'h179c0:	data_out=16'h8007;
17'h179c1:	data_out=16'h8000;
17'h179c2:	data_out=16'h8001;
17'h179c3:	data_out=16'h8005;
17'h179c4:	data_out=16'h8009;
17'h179c5:	data_out=16'h4;
17'h179c6:	data_out=16'h4;
17'h179c7:	data_out=16'h8002;
17'h179c8:	data_out=16'h8007;
17'h179c9:	data_out=16'h3;
17'h179ca:	data_out=16'h8000;
17'h179cb:	data_out=16'h8003;
17'h179cc:	data_out=16'h3;
17'h179cd:	data_out=16'h8002;
17'h179ce:	data_out=16'h4;
17'h179cf:	data_out=16'h2;
17'h179d0:	data_out=16'h8006;
17'h179d1:	data_out=16'h5;
17'h179d2:	data_out=16'h4;
17'h179d3:	data_out=16'h8002;
17'h179d4:	data_out=16'h5;
17'h179d5:	data_out=16'h8005;
17'h179d6:	data_out=16'h8;
17'h179d7:	data_out=16'h8002;
17'h179d8:	data_out=16'h7;
17'h179d9:	data_out=16'h8000;
17'h179da:	data_out=16'h8001;
17'h179db:	data_out=16'h0;
17'h179dc:	data_out=16'h1;
17'h179dd:	data_out=16'h7;
17'h179de:	data_out=16'h8005;
17'h179df:	data_out=16'h3;
17'h179e0:	data_out=16'h8003;
17'h179e1:	data_out=16'h3;
17'h179e2:	data_out=16'h7;
17'h179e3:	data_out=16'h8002;
17'h179e4:	data_out=16'h8003;
17'h179e5:	data_out=16'h2;
17'h179e6:	data_out=16'h5;
17'h179e7:	data_out=16'h8001;
17'h179e8:	data_out=16'h8005;
17'h179e9:	data_out=16'h8005;
17'h179ea:	data_out=16'h6;
17'h179eb:	data_out=16'h8;
17'h179ec:	data_out=16'h3;
17'h179ed:	data_out=16'h0;
17'h179ee:	data_out=16'h1;
17'h179ef:	data_out=16'h6;
17'h179f0:	data_out=16'h8004;
17'h179f1:	data_out=16'h8004;
17'h179f2:	data_out=16'h8006;
17'h179f3:	data_out=16'h8009;
17'h179f4:	data_out=16'h0;
17'h179f5:	data_out=16'h8007;
17'h179f6:	data_out=16'h8001;
17'h179f7:	data_out=16'h8003;
17'h179f8:	data_out=16'h2;
17'h179f9:	data_out=16'h7;
17'h179fa:	data_out=16'h7;
17'h179fb:	data_out=16'h8006;
17'h179fc:	data_out=16'h4;
17'h179fd:	data_out=16'h8007;
17'h179fe:	data_out=16'h6;
17'h179ff:	data_out=16'h8008;
17'h17a00:	data_out=16'h4;
17'h17a01:	data_out=16'h4;
17'h17a02:	data_out=16'h8001;
17'h17a03:	data_out=16'h8007;
17'h17a04:	data_out=16'h8003;
17'h17a05:	data_out=16'h8005;
17'h17a06:	data_out=16'h1;
17'h17a07:	data_out=16'h1;
17'h17a08:	data_out=16'h8001;
17'h17a09:	data_out=16'h8003;
17'h17a0a:	data_out=16'h0;
17'h17a0b:	data_out=16'h8008;
17'h17a0c:	data_out=16'h7;
17'h17a0d:	data_out=16'h8008;
17'h17a0e:	data_out=16'h8;
17'h17a0f:	data_out=16'h8007;
17'h17a10:	data_out=16'h8003;
17'h17a11:	data_out=16'h8007;
17'h17a12:	data_out=16'h8006;
17'h17a13:	data_out=16'h6;
17'h17a14:	data_out=16'h8005;
17'h17a15:	data_out=16'h1;
17'h17a16:	data_out=16'h8005;
17'h17a17:	data_out=16'h7;
17'h17a18:	data_out=16'h8001;
17'h17a19:	data_out=16'h8007;
17'h17a1a:	data_out=16'h8009;
17'h17a1b:	data_out=16'h8006;
17'h17a1c:	data_out=16'h8006;
17'h17a1d:	data_out=16'h6;
17'h17a1e:	data_out=16'h8005;
17'h17a1f:	data_out=16'h8;
17'h17a20:	data_out=16'h1;
17'h17a21:	data_out=16'h4;
17'h17a22:	data_out=16'h8009;
17'h17a23:	data_out=16'h7;
17'h17a24:	data_out=16'h7;
17'h17a25:	data_out=16'h1;
17'h17a26:	data_out=16'h8001;
17'h17a27:	data_out=16'h8003;
17'h17a28:	data_out=16'h8;
17'h17a29:	data_out=16'h8;
17'h17a2a:	data_out=16'h8001;
17'h17a2b:	data_out=16'h5;
17'h17a2c:	data_out=16'h8009;
17'h17a2d:	data_out=16'h8003;
17'h17a2e:	data_out=16'h8;
17'h17a2f:	data_out=16'h8002;
17'h17a30:	data_out=16'h8001;
17'h17a31:	data_out=16'h8008;
17'h17a32:	data_out=16'h8005;
17'h17a33:	data_out=16'h4;
17'h17a34:	data_out=16'h3;
17'h17a35:	data_out=16'h8001;
17'h17a36:	data_out=16'h1;
17'h17a37:	data_out=16'h8008;
17'h17a38:	data_out=16'h1;
17'h17a39:	data_out=16'h2;
17'h17a3a:	data_out=16'h8004;
17'h17a3b:	data_out=16'h4;
17'h17a3c:	data_out=16'h8001;
17'h17a3d:	data_out=16'h0;
17'h17a3e:	data_out=16'h3;
17'h17a3f:	data_out=16'h8009;
17'h17a40:	data_out=16'h8006;
17'h17a41:	data_out=16'h3;
17'h17a42:	data_out=16'h7;
17'h17a43:	data_out=16'h8007;
17'h17a44:	data_out=16'h8005;
17'h17a45:	data_out=16'h8003;
17'h17a46:	data_out=16'h8001;
17'h17a47:	data_out=16'h8006;
17'h17a48:	data_out=16'h8004;
17'h17a49:	data_out=16'h7;
17'h17a4a:	data_out=16'h8;
17'h17a4b:	data_out=16'h8004;
17'h17a4c:	data_out=16'h8005;
17'h17a4d:	data_out=16'h6;
17'h17a4e:	data_out=16'h3;
17'h17a4f:	data_out=16'h3;
17'h17a50:	data_out=16'h7;
17'h17a51:	data_out=16'h7;
17'h17a52:	data_out=16'h8003;
17'h17a53:	data_out=16'h1;
17'h17a54:	data_out=16'h8004;
17'h17a55:	data_out=16'h8;
17'h17a56:	data_out=16'h3;
17'h17a57:	data_out=16'h6;
17'h17a58:	data_out=16'h8000;
17'h17a59:	data_out=16'h7;
17'h17a5a:	data_out=16'h1;
17'h17a5b:	data_out=16'h8;
17'h17a5c:	data_out=16'h8002;
17'h17a5d:	data_out=16'h8006;
17'h17a5e:	data_out=16'h8;
17'h17a5f:	data_out=16'h2;
17'h17a60:	data_out=16'h6;
17'h17a61:	data_out=16'h6;
17'h17a62:	data_out=16'h4;
17'h17a63:	data_out=16'h8008;
17'h17a64:	data_out=16'h8006;
17'h17a65:	data_out=16'h8007;
17'h17a66:	data_out=16'h8005;
17'h17a67:	data_out=16'h8001;
17'h17a68:	data_out=16'h8009;
17'h17a69:	data_out=16'h8006;
17'h17a6a:	data_out=16'h4;
17'h17a6b:	data_out=16'h8005;
17'h17a6c:	data_out=16'h9;
17'h17a6d:	data_out=16'h8003;
17'h17a6e:	data_out=16'h7;
17'h17a6f:	data_out=16'h7;
17'h17a70:	data_out=16'h8005;
17'h17a71:	data_out=16'h8005;
17'h17a72:	data_out=16'h8001;
17'h17a73:	data_out=16'h1;
17'h17a74:	data_out=16'h8006;
17'h17a75:	data_out=16'h8007;
17'h17a76:	data_out=16'h8002;
17'h17a77:	data_out=16'h3;
17'h17a78:	data_out=16'h8009;
17'h17a79:	data_out=16'h8;
17'h17a7a:	data_out=16'h2;
17'h17a7b:	data_out=16'h8001;
17'h17a7c:	data_out=16'h8007;
17'h17a7d:	data_out=16'h1;
17'h17a7e:	data_out=16'h8009;
17'h17a7f:	data_out=16'h8;
17'h17a80:	data_out=16'h8002;
17'h17a81:	data_out=16'h4;
17'h17a82:	data_out=16'h8008;
17'h17a83:	data_out=16'h0;
17'h17a84:	data_out=16'h7;
17'h17a85:	data_out=16'h8004;
17'h17a86:	data_out=16'h8;
17'h17a87:	data_out=16'h7;
17'h17a88:	data_out=16'h8001;
17'h17a89:	data_out=16'h3;
17'h17a8a:	data_out=16'h8007;
17'h17a8b:	data_out=16'h8002;
17'h17a8c:	data_out=16'h8009;
17'h17a8d:	data_out=16'h8009;
17'h17a8e:	data_out=16'h8003;
17'h17a8f:	data_out=16'h8005;
17'h17a90:	data_out=16'h8004;
17'h17a91:	data_out=16'h5;
17'h17a92:	data_out=16'h5;
17'h17a93:	data_out=16'h8001;
17'h17a94:	data_out=16'h7;
17'h17a95:	data_out=16'h8006;
17'h17a96:	data_out=16'h8008;
17'h17a97:	data_out=16'h8;
17'h17a98:	data_out=16'h8008;
17'h17a99:	data_out=16'h3;
17'h17a9a:	data_out=16'h8003;
17'h17a9b:	data_out=16'h8006;
17'h17a9c:	data_out=16'h8005;
17'h17a9d:	data_out=16'h8003;
17'h17a9e:	data_out=16'h8007;
17'h17a9f:	data_out=16'h1;
17'h17aa0:	data_out=16'h8008;
17'h17aa1:	data_out=16'h8006;
17'h17aa2:	data_out=16'h8007;
17'h17aa3:	data_out=16'h8;
17'h17aa4:	data_out=16'h8001;
17'h17aa5:	data_out=16'h8009;
17'h17aa6:	data_out=16'h6;
17'h17aa7:	data_out=16'h7;
17'h17aa8:	data_out=16'h3;
17'h17aa9:	data_out=16'h8;
17'h17aaa:	data_out=16'h8004;
17'h17aab:	data_out=16'h3;
17'h17aac:	data_out=16'h8;
17'h17aad:	data_out=16'h2;
17'h17aae:	data_out=16'h8;
17'h17aaf:	data_out=16'h8006;
17'h17ab0:	data_out=16'h8002;
17'h17ab1:	data_out=16'h4;
17'h17ab2:	data_out=16'h2;
17'h17ab3:	data_out=16'h8004;
17'h17ab4:	data_out=16'h6;
17'h17ab5:	data_out=16'h3;
17'h17ab6:	data_out=16'h8005;
17'h17ab7:	data_out=16'h7;
17'h17ab8:	data_out=16'h8002;
17'h17ab9:	data_out=16'h1;
17'h17aba:	data_out=16'h8008;
17'h17abb:	data_out=16'h1;
17'h17abc:	data_out=16'h7;
17'h17abd:	data_out=16'h8005;
17'h17abe:	data_out=16'h8006;
17'h17abf:	data_out=16'h9;
17'h17ac0:	data_out=16'h8002;
17'h17ac1:	data_out=16'h8004;
17'h17ac2:	data_out=16'h8;
17'h17ac3:	data_out=16'h7;
17'h17ac4:	data_out=16'h8004;
17'h17ac5:	data_out=16'h5;
17'h17ac6:	data_out=16'h4;
17'h17ac7:	data_out=16'h9;
17'h17ac8:	data_out=16'h3;
17'h17ac9:	data_out=16'h8009;
17'h17aca:	data_out=16'h3;
17'h17acb:	data_out=16'h2;
17'h17acc:	data_out=16'h2;
17'h17acd:	data_out=16'h1;
17'h17ace:	data_out=16'h6;
17'h17acf:	data_out=16'h8009;
17'h17ad0:	data_out=16'h8004;
17'h17ad1:	data_out=16'h8001;
17'h17ad2:	data_out=16'h8003;
17'h17ad3:	data_out=16'h8007;
17'h17ad4:	data_out=16'h8007;
17'h17ad5:	data_out=16'h0;
17'h17ad6:	data_out=16'h8009;
17'h17ad7:	data_out=16'h8000;
17'h17ad8:	data_out=16'h8008;
17'h17ad9:	data_out=16'h8007;
17'h17ada:	data_out=16'h8008;
17'h17adb:	data_out=16'h9;
17'h17adc:	data_out=16'h8003;
17'h17add:	data_out=16'h8005;
17'h17ade:	data_out=16'h8;
17'h17adf:	data_out=16'h4;
17'h17ae0:	data_out=16'h8001;
17'h17ae1:	data_out=16'h7;
17'h17ae2:	data_out=16'h2;
17'h17ae3:	data_out=16'h5;
17'h17ae4:	data_out=16'h2;
17'h17ae5:	data_out=16'h8003;
17'h17ae6:	data_out=16'h4;
17'h17ae7:	data_out=16'h8004;
17'h17ae8:	data_out=16'h8003;
17'h17ae9:	data_out=16'h8002;
17'h17aea:	data_out=16'h8;
17'h17aeb:	data_out=16'h8;
17'h17aec:	data_out=16'h8;
17'h17aed:	data_out=16'h4;
17'h17aee:	data_out=16'h9;
17'h17aef:	data_out=16'h8005;
17'h17af0:	data_out=16'h8007;
17'h17af1:	data_out=16'h8004;
17'h17af2:	data_out=16'h8003;
17'h17af3:	data_out=16'h8004;
17'h17af4:	data_out=16'h6;
17'h17af5:	data_out=16'h8003;
17'h17af6:	data_out=16'h4;
17'h17af7:	data_out=16'h7;
17'h17af8:	data_out=16'h8001;
17'h17af9:	data_out=16'h5;
17'h17afa:	data_out=16'h6;
17'h17afb:	data_out=16'h5;
17'h17afc:	data_out=16'h8009;
17'h17afd:	data_out=16'h5;
17'h17afe:	data_out=16'h0;
17'h17aff:	data_out=16'h8001;
17'h17b00:	data_out=16'h3;
17'h17b01:	data_out=16'h8007;
17'h17b02:	data_out=16'h8005;
17'h17b03:	data_out=16'h8004;
17'h17b04:	data_out=16'h8001;
17'h17b05:	data_out=16'h8;
17'h17b06:	data_out=16'h2;
17'h17b07:	data_out=16'h5;
17'h17b08:	data_out=16'h8003;
17'h17b09:	data_out=16'h0;
17'h17b0a:	data_out=16'h4;
17'h17b0b:	data_out=16'h8004;
17'h17b0c:	data_out=16'h8005;
17'h17b0d:	data_out=16'h4;
17'h17b0e:	data_out=16'h8000;
17'h17b0f:	data_out=16'h8002;
17'h17b10:	data_out=16'h9;
17'h17b11:	data_out=16'h6;
17'h17b12:	data_out=16'h2;
17'h17b13:	data_out=16'h5;
17'h17b14:	data_out=16'h8007;
17'h17b15:	data_out=16'h8003;
17'h17b16:	data_out=16'h3;
17'h17b17:	data_out=16'h1;
17'h17b18:	data_out=16'h8006;
17'h17b19:	data_out=16'h8000;
17'h17b1a:	data_out=16'h8003;
17'h17b1b:	data_out=16'h8006;
17'h17b1c:	data_out=16'h8004;
17'h17b1d:	data_out=16'h7;
17'h17b1e:	data_out=16'h2;
17'h17b1f:	data_out=16'h8;
17'h17b20:	data_out=16'h8;
17'h17b21:	data_out=16'h6;
17'h17b22:	data_out=16'h8005;
17'h17b23:	data_out=16'h8002;
17'h17b24:	data_out=16'h5;
17'h17b25:	data_out=16'h5;
17'h17b26:	data_out=16'h8006;
17'h17b27:	data_out=16'h8007;
17'h17b28:	data_out=16'h8004;
17'h17b29:	data_out=16'h7;
17'h17b2a:	data_out=16'h8002;
17'h17b2b:	data_out=16'h0;
17'h17b2c:	data_out=16'h1;
17'h17b2d:	data_out=16'h7;
17'h17b2e:	data_out=16'h7;
17'h17b2f:	data_out=16'h1;
17'h17b30:	data_out=16'h3;
17'h17b31:	data_out=16'h0;
17'h17b32:	data_out=16'h8003;
17'h17b33:	data_out=16'h6;
17'h17b34:	data_out=16'h7;
17'h17b35:	data_out=16'h9;
17'h17b36:	data_out=16'h8002;
17'h17b37:	data_out=16'h8009;
17'h17b38:	data_out=16'h8001;
17'h17b39:	data_out=16'h4;
17'h17b3a:	data_out=16'h8006;
17'h17b3b:	data_out=16'h4;
17'h17b3c:	data_out=16'h2;
17'h17b3d:	data_out=16'h5;
17'h17b3e:	data_out=16'h2;
17'h17b3f:	data_out=16'h1;
17'h17b40:	data_out=16'h2;
17'h17b41:	data_out=16'h6;
17'h17b42:	data_out=16'h8;
17'h17b43:	data_out=16'h8001;
17'h17b44:	data_out=16'h2;
17'h17b45:	data_out=16'h8007;
17'h17b46:	data_out=16'h1;
17'h17b47:	data_out=16'h7;
17'h17b48:	data_out=16'h9;
17'h17b49:	data_out=16'h8;
17'h17b4a:	data_out=16'h8002;
17'h17b4b:	data_out=16'h1;
17'h17b4c:	data_out=16'h6;
17'h17b4d:	data_out=16'h8004;
17'h17b4e:	data_out=16'h8007;
17'h17b4f:	data_out=16'h8000;
17'h17b50:	data_out=16'h6;
17'h17b51:	data_out=16'h8001;
17'h17b52:	data_out=16'h8004;
17'h17b53:	data_out=16'h3;
17'h17b54:	data_out=16'h8002;
17'h17b55:	data_out=16'h3;
17'h17b56:	data_out=16'h4;
17'h17b57:	data_out=16'h6;
17'h17b58:	data_out=16'h8001;
17'h17b59:	data_out=16'h7;
17'h17b5a:	data_out=16'h1;
17'h17b5b:	data_out=16'h8009;
17'h17b5c:	data_out=16'h3;
17'h17b5d:	data_out=16'h8006;
17'h17b5e:	data_out=16'h1;
17'h17b5f:	data_out=16'h8004;
17'h17b60:	data_out=16'h9;
17'h17b61:	data_out=16'h0;
17'h17b62:	data_out=16'h4;
17'h17b63:	data_out=16'h2;
17'h17b64:	data_out=16'h2;
17'h17b65:	data_out=16'h8005;
17'h17b66:	data_out=16'h0;
17'h17b67:	data_out=16'h2;
17'h17b68:	data_out=16'h8006;
17'h17b69:	data_out=16'h8;
17'h17b6a:	data_out=16'h8007;
17'h17b6b:	data_out=16'h9;
17'h17b6c:	data_out=16'h8005;
17'h17b6d:	data_out=16'h8005;
17'h17b6e:	data_out=16'h8001;
17'h17b6f:	data_out=16'h8009;
17'h17b70:	data_out=16'h3;
17'h17b71:	data_out=16'h5;
17'h17b72:	data_out=16'h4;
17'h17b73:	data_out=16'h8008;
17'h17b74:	data_out=16'h8001;
17'h17b75:	data_out=16'h8002;
17'h17b76:	data_out=16'h7;
17'h17b77:	data_out=16'h7;
17'h17b78:	data_out=16'h8005;
17'h17b79:	data_out=16'h8002;
17'h17b7a:	data_out=16'h7;
17'h17b7b:	data_out=16'h7;
17'h17b7c:	data_out=16'h1;
17'h17b7d:	data_out=16'h8001;
17'h17b7e:	data_out=16'h8006;
17'h17b7f:	data_out=16'h1;
17'h17b80:	data_out=16'h9;
17'h17b81:	data_out=16'h6;
17'h17b82:	data_out=16'h8006;
17'h17b83:	data_out=16'h2;
17'h17b84:	data_out=16'h8008;
17'h17b85:	data_out=16'h3;
17'h17b86:	data_out=16'h8006;
17'h17b87:	data_out=16'h8004;
17'h17b88:	data_out=16'h2;
17'h17b89:	data_out=16'h8003;
17'h17b8a:	data_out=16'h8004;
17'h17b8b:	data_out=16'h6;
17'h17b8c:	data_out=16'h1;
17'h17b8d:	data_out=16'h4;
17'h17b8e:	data_out=16'h6;
17'h17b8f:	data_out=16'h8006;
17'h17b90:	data_out=16'h8000;
17'h17b91:	data_out=16'h1;
17'h17b92:	data_out=16'h8005;
17'h17b93:	data_out=16'h8;
17'h17b94:	data_out=16'h8;
17'h17b95:	data_out=16'h8007;
17'h17b96:	data_out=16'h5;
17'h17b97:	data_out=16'h8006;
17'h17b98:	data_out=16'h0;
17'h17b99:	data_out=16'h3;
17'h17b9a:	data_out=16'h8008;
17'h17b9b:	data_out=16'h8007;
17'h17b9c:	data_out=16'h8007;
17'h17b9d:	data_out=16'h8005;
17'h17b9e:	data_out=16'h3;
17'h17b9f:	data_out=16'h8008;
17'h17ba0:	data_out=16'h8008;
17'h17ba1:	data_out=16'h6;
17'h17ba2:	data_out=16'h3;
17'h17ba3:	data_out=16'h8007;
17'h17ba4:	data_out=16'h1;
17'h17ba5:	data_out=16'h6;
17'h17ba6:	data_out=16'h8002;
17'h17ba7:	data_out=16'h8007;
17'h17ba8:	data_out=16'h8007;
17'h17ba9:	data_out=16'h3;
17'h17baa:	data_out=16'h8;
17'h17bab:	data_out=16'h3;
17'h17bac:	data_out=16'h8002;
17'h17bad:	data_out=16'h5;
17'h17bae:	data_out=16'h7;
17'h17baf:	data_out=16'h7;
17'h17bb0:	data_out=16'h8003;
17'h17bb1:	data_out=16'h8007;
17'h17bb2:	data_out=16'h5;
17'h17bb3:	data_out=16'h8005;
17'h17bb4:	data_out=16'h8005;
17'h17bb5:	data_out=16'h1;
17'h17bb6:	data_out=16'h8002;
17'h17bb7:	data_out=16'h5;
17'h17bb8:	data_out=16'h8005;
17'h17bb9:	data_out=16'h8001;
17'h17bba:	data_out=16'h6;
17'h17bbb:	data_out=16'h8003;
17'h17bbc:	data_out=16'h3;
17'h17bbd:	data_out=16'h0;
17'h17bbe:	data_out=16'h8002;
17'h17bbf:	data_out=16'h4;
17'h17bc0:	data_out=16'h8002;
17'h17bc1:	data_out=16'h8009;
17'h17bc2:	data_out=16'h7;
17'h17bc3:	data_out=16'h8;
17'h17bc4:	data_out=16'h7;
17'h17bc5:	data_out=16'h8004;
17'h17bc6:	data_out=16'h8008;
17'h17bc7:	data_out=16'h8009;
17'h17bc8:	data_out=16'h8;
17'h17bc9:	data_out=16'h8009;
17'h17bca:	data_out=16'h4;
17'h17bcb:	data_out=16'h8003;
17'h17bcc:	data_out=16'h5;
17'h17bcd:	data_out=16'h2;
17'h17bce:	data_out=16'h8006;
17'h17bcf:	data_out=16'h8007;
17'h17bd0:	data_out=16'h4;
17'h17bd1:	data_out=16'h9;
17'h17bd2:	data_out=16'h8003;
17'h17bd3:	data_out=16'h8;
17'h17bd4:	data_out=16'h1;
17'h17bd5:	data_out=16'h5;
17'h17bd6:	data_out=16'h3;
17'h17bd7:	data_out=16'h5;
17'h17bd8:	data_out=16'h8005;
17'h17bd9:	data_out=16'h1;
17'h17bda:	data_out=16'h8007;
17'h17bdb:	data_out=16'h7;
17'h17bdc:	data_out=16'h8008;
17'h17bdd:	data_out=16'h8000;
17'h17bde:	data_out=16'h2;
17'h17bdf:	data_out=16'h8001;
17'h17be0:	data_out=16'h0;
17'h17be1:	data_out=16'h8000;
17'h17be2:	data_out=16'h8003;
17'h17be3:	data_out=16'h8002;
17'h17be4:	data_out=16'h5;
17'h17be5:	data_out=16'h8002;
17'h17be6:	data_out=16'h8002;
17'h17be7:	data_out=16'h4;
17'h17be8:	data_out=16'h8002;
17'h17be9:	data_out=16'h8008;
17'h17bea:	data_out=16'h8008;
17'h17beb:	data_out=16'h8005;
17'h17bec:	data_out=16'h3;
17'h17bed:	data_out=16'h8005;
17'h17bee:	data_out=16'h8004;
17'h17bef:	data_out=16'h8002;
17'h17bf0:	data_out=16'h8005;
17'h17bf1:	data_out=16'h3;
17'h17bf2:	data_out=16'h8004;
17'h17bf3:	data_out=16'h5;
17'h17bf4:	data_out=16'h8002;
17'h17bf5:	data_out=16'h9;
17'h17bf6:	data_out=16'h1;
17'h17bf7:	data_out=16'h2;
17'h17bf8:	data_out=16'h0;
17'h17bf9:	data_out=16'h3;
17'h17bfa:	data_out=16'h8000;
17'h17bfb:	data_out=16'h1;
17'h17bfc:	data_out=16'h8006;
17'h17bfd:	data_out=16'h8007;
17'h17bfe:	data_out=16'h9;
17'h17bff:	data_out=16'h3;
17'h17c00:	data_out=16'h19;
17'h17c01:	data_out=16'h1f;
17'h17c02:	data_out=16'h18;
17'h17c03:	data_out=16'h1e;
17'h17c04:	data_out=16'h30;
17'h17c05:	data_out=16'h2c;
17'h17c06:	data_out=16'h5;
17'h17c07:	data_out=16'h1c;
17'h17c08:	data_out=16'h1c;
17'h17c09:	data_out=16'hb;
17'h17c0a:	data_out=16'h1e;
17'h17c0b:	data_out=16'hb;
17'h17c0c:	data_out=16'h2e;
17'h17c0d:	data_out=16'h1e;
17'h17c0e:	data_out=16'h8;
17'h17c0f:	data_out=16'h22;
17'h17c10:	data_out=16'h13;
17'h17c11:	data_out=16'h2c;
17'h17c12:	data_out=16'h24;
17'h17c13:	data_out=16'h1d;
17'h17c14:	data_out=16'h1f;
17'h17c15:	data_out=16'ha;
17'h17c16:	data_out=16'h19;
17'h17c17:	data_out=16'h16;
17'h17c18:	data_out=16'he;
17'h17c19:	data_out=16'h14;
17'h17c1a:	data_out=16'h2b;
17'h17c1b:	data_out=16'h20;
17'h17c1c:	data_out=16'h3a;
17'h17c1d:	data_out=16'h3b;
17'h17c1e:	data_out=16'h26;
17'h17c1f:	data_out=16'h1d;
17'h17c20:	data_out=16'h2f;
17'h17c21:	data_out=16'h8;
17'h17c22:	data_out=16'h26;
17'h17c23:	data_out=16'h14;
17'h17c24:	data_out=16'h14;
17'h17c25:	data_out=16'h1e;
17'h17c26:	data_out=16'hc;
17'h17c27:	data_out=16'h36;
17'h17c28:	data_out=16'h3;
17'h17c29:	data_out=16'h19;
17'h17c2a:	data_out=16'h21;
17'h17c2b:	data_out=16'h17;
17'h17c2c:	data_out=16'h18;
17'h17c2d:	data_out=16'hd;
17'h17c2e:	data_out=16'h18;
17'h17c2f:	data_out=16'h2a;
17'h17c30:	data_out=16'h20;
17'h17c31:	data_out=16'h20;
17'h17c32:	data_out=16'h26;
17'h17c33:	data_out=16'h24;
17'h17c34:	data_out=16'h1f;
17'h17c35:	data_out=16'h32;
17'h17c36:	data_out=16'h1b;
17'h17c37:	data_out=16'h24;
17'h17c38:	data_out=16'h14;
17'h17c39:	data_out=16'h1d;
17'h17c3a:	data_out=16'h28;
17'h17c3b:	data_out=16'h1d;
17'h17c3c:	data_out=16'h25;
17'h17c3d:	data_out=16'h28;
17'h17c3e:	data_out=16'h10;
17'h17c3f:	data_out=16'h20;
17'h17c40:	data_out=16'h36;
17'h17c41:	data_out=16'h2c;
17'h17c42:	data_out=16'h15;
17'h17c43:	data_out=16'ha;
17'h17c44:	data_out=16'h2b;
17'h17c45:	data_out=16'h8;
17'h17c46:	data_out=16'h22;
17'h17c47:	data_out=16'h29;
17'h17c48:	data_out=16'h1f;
17'h17c49:	data_out=16'h2b;
17'h17c4a:	data_out=16'h35;
17'h17c4b:	data_out=16'h25;
17'h17c4c:	data_out=16'h2c;
17'h17c4d:	data_out=16'h1e;
17'h17c4e:	data_out=16'h30;
17'h17c4f:	data_out=16'h2c;
17'h17c50:	data_out=16'h2a;
17'h17c51:	data_out=16'h1f;
17'h17c52:	data_out=16'hd;
17'h17c53:	data_out=16'h4c;
17'h17c54:	data_out=16'h2e;
17'h17c55:	data_out=16'h14;
17'h17c56:	data_out=16'h1b;
17'h17c57:	data_out=16'h12;
17'h17c58:	data_out=16'h18;
17'h17c59:	data_out=16'h2e;
17'h17c5a:	data_out=16'he;
17'h17c5b:	data_out=16'h1d;
17'h17c5c:	data_out=16'h24;
17'h17c5d:	data_out=16'h23;
17'h17c5e:	data_out=16'h2d;
17'h17c5f:	data_out=16'hf;
17'h17c60:	data_out=16'h16;
17'h17c61:	data_out=16'h2a;
17'h17c62:	data_out=16'h1e;
17'h17c63:	data_out=16'h1c;
17'h17c64:	data_out=16'h26;
17'h17c65:	data_out=16'h27;
17'h17c66:	data_out=16'h16;
17'h17c67:	data_out=16'h24;
17'h17c68:	data_out=16'h2;
17'h17c69:	data_out=16'h19;
17'h17c6a:	data_out=16'he;
17'h17c6b:	data_out=16'h1c;
17'h17c6c:	data_out=16'h23;
17'h17c6d:	data_out=16'h1f;
17'h17c6e:	data_out=16'hd;
17'h17c6f:	data_out=16'h3a;
17'h17c70:	data_out=16'h8;
17'h17c71:	data_out=16'h14;
17'h17c72:	data_out=16'h1f;
17'h17c73:	data_out=16'h1c;
17'h17c74:	data_out=16'h23;
17'h17c75:	data_out=16'h14;
17'h17c76:	data_out=16'h13;
17'h17c77:	data_out=16'h28;
17'h17c78:	data_out=16'h6;
17'h17c79:	data_out=16'h24;
17'h17c7a:	data_out=16'h1b;
17'h17c7b:	data_out=16'hd;
17'h17c7c:	data_out=16'h1;
17'h17c7d:	data_out=16'hb;
17'h17c7e:	data_out=16'h18;
17'h17c7f:	data_out=16'h23;
17'h17c80:	data_out=16'h126;
17'h17c81:	data_out=16'h16b;
17'h17c82:	data_out=16'hc0;
17'h17c83:	data_out=16'h101;
17'h17c84:	data_out=16'h179;
17'h17c85:	data_out=16'h18e;
17'h17c86:	data_out=16'h9b;
17'h17c87:	data_out=16'h12d;
17'h17c88:	data_out=16'hdc;
17'h17c89:	data_out=16'h74;
17'h17c8a:	data_out=16'h127;
17'h17c8b:	data_out=16'h73;
17'h17c8c:	data_out=16'h153;
17'h17c8d:	data_out=16'hd7;
17'h17c8e:	data_out=16'h39;
17'h17c8f:	data_out=16'h117;
17'h17c90:	data_out=16'h4f;
17'h17c91:	data_out=16'h160;
17'h17c92:	data_out=16'hd5;
17'h17c93:	data_out=16'hf4;
17'h17c94:	data_out=16'hbb;
17'h17c95:	data_out=16'hc3;
17'h17c96:	data_out=16'h129;
17'h17c97:	data_out=16'hc9;
17'h17c98:	data_out=16'h70;
17'h17c99:	data_out=16'hc2;
17'h17c9a:	data_out=16'h183;
17'h17c9b:	data_out=16'he6;
17'h17c9c:	data_out=16'h1ac;
17'h17c9d:	data_out=16'h192;
17'h17c9e:	data_out=16'h11a;
17'h17c9f:	data_out=16'hc6;
17'h17ca0:	data_out=16'h1ce;
17'h17ca1:	data_out=16'h44;
17'h17ca2:	data_out=16'h9b;
17'h17ca3:	data_out=16'h77;
17'h17ca4:	data_out=16'h69;
17'h17ca5:	data_out=16'hb6;
17'h17ca6:	data_out=16'h66;
17'h17ca7:	data_out=16'h1b5;
17'h17ca8:	data_out=16'h37;
17'h17ca9:	data_out=16'hc3;
17'h17caa:	data_out=16'hf2;
17'h17cab:	data_out=16'hb7;
17'h17cac:	data_out=16'hfb;
17'h17cad:	data_out=16'h8e;
17'h17cae:	data_out=16'hb2;
17'h17caf:	data_out=16'h18e;
17'h17cb0:	data_out=16'h1c0;
17'h17cb1:	data_out=16'h14f;
17'h17cb2:	data_out=16'h1c8;
17'h17cb3:	data_out=16'he1;
17'h17cb4:	data_out=16'h123;
17'h17cb5:	data_out=16'h1bf;
17'h17cb6:	data_out=16'hf4;
17'h17cb7:	data_out=16'hc0;
17'h17cb8:	data_out=16'h13d;
17'h17cb9:	data_out=16'hb3;
17'h17cba:	data_out=16'hcd;
17'h17cbb:	data_out=16'h13b;
17'h17cbc:	data_out=16'hb0;
17'h17cbd:	data_out=16'h14b;
17'h17cbe:	data_out=16'h43;
17'h17cbf:	data_out=16'h183;
17'h17cc0:	data_out=16'h150;
17'h17cc1:	data_out=16'he0;
17'h17cc2:	data_out=16'hc1;
17'h17cc3:	data_out=16'h52;
17'h17cc4:	data_out=16'h141;
17'h17cc5:	data_out=16'h90;
17'h17cc6:	data_out=16'h77;
17'h17cc7:	data_out=16'heb;
17'h17cc8:	data_out=16'hb6;
17'h17cc9:	data_out=16'hbe;
17'h17cca:	data_out=16'h193;
17'h17ccb:	data_out=16'h12a;
17'h17ccc:	data_out=16'hec;
17'h17ccd:	data_out=16'hd6;
17'h17cce:	data_out=16'h169;
17'h17ccf:	data_out=16'hf9;
17'h17cd0:	data_out=16'h101;
17'h17cd1:	data_out=16'hc4;
17'h17cd2:	data_out=16'h7f;
17'h17cd3:	data_out=16'h21e;
17'h17cd4:	data_out=16'h1a4;
17'h17cd5:	data_out=16'h29;
17'h17cd6:	data_out=16'ha8;
17'h17cd7:	data_out=16'h4b;
17'h17cd8:	data_out=16'h2e;
17'h17cd9:	data_out=16'h100;
17'h17cda:	data_out=16'h5f;
17'h17cdb:	data_out=16'h16d;
17'h17cdc:	data_out=16'h14d;
17'h17cdd:	data_out=16'h145;
17'h17cde:	data_out=16'h197;
17'h17cdf:	data_out=16'hb0;
17'h17ce0:	data_out=16'h9f;
17'h17ce1:	data_out=16'h190;
17'h17ce2:	data_out=16'hca;
17'h17ce3:	data_out=16'he6;
17'h17ce4:	data_out=16'hfa;
17'h17ce5:	data_out=16'h123;
17'h17ce6:	data_out=16'hb4;
17'h17ce7:	data_out=16'hc7;
17'h17ce8:	data_out=16'h43;
17'h17ce9:	data_out=16'h96;
17'h17cea:	data_out=16'h40;
17'h17ceb:	data_out=16'h188;
17'h17cec:	data_out=16'h119;
17'h17ced:	data_out=16'he6;
17'h17cee:	data_out=16'h3c;
17'h17cef:	data_out=16'h1b6;
17'h17cf0:	data_out=16'h3f;
17'h17cf1:	data_out=16'hd0;
17'h17cf2:	data_out=16'h132;
17'h17cf3:	data_out=16'h190;
17'h17cf4:	data_out=16'h1b4;
17'h17cf5:	data_out=16'h12c;
17'h17cf6:	data_out=16'haa;
17'h17cf7:	data_out=16'hc7;
17'h17cf8:	data_out=16'ha9;
17'h17cf9:	data_out=16'hfe;
17'h17cfa:	data_out=16'hc9;
17'h17cfb:	data_out=16'h49;
17'h17cfc:	data_out=16'h63;
17'h17cfd:	data_out=16'hc9;
17'h17cfe:	data_out=16'h56;
17'h17cff:	data_out=16'h11c;
17'h17d00:	data_out=16'h1d7;
17'h17d01:	data_out=16'h24b;
17'h17d02:	data_out=16'h1b2;
17'h17d03:	data_out=16'h25e;
17'h17d04:	data_out=16'h279;
17'h17d05:	data_out=16'h2b8;
17'h17d06:	data_out=16'h167;
17'h17d07:	data_out=16'h1dc;
17'h17d08:	data_out=16'h1af;
17'h17d09:	data_out=16'h11a;
17'h17d0a:	data_out=16'h1c5;
17'h17d0b:	data_out=16'h166;
17'h17d0c:	data_out=16'h21d;
17'h17d0d:	data_out=16'h1ce;
17'h17d0e:	data_out=16'h96;
17'h17d0f:	data_out=16'h23c;
17'h17d10:	data_out=16'h103;
17'h17d11:	data_out=16'h251;
17'h17d12:	data_out=16'h1ab;
17'h17d13:	data_out=16'h247;
17'h17d14:	data_out=16'h1b0;
17'h17d15:	data_out=16'h16e;
17'h17d16:	data_out=16'h209;
17'h17d17:	data_out=16'h1d6;
17'h17d18:	data_out=16'he3;
17'h17d19:	data_out=16'h130;
17'h17d1a:	data_out=16'h297;
17'h17d1b:	data_out=16'h1d9;
17'h17d1c:	data_out=16'h2d7;
17'h17d1d:	data_out=16'h2ab;
17'h17d1e:	data_out=16'h20c;
17'h17d1f:	data_out=16'h1b5;
17'h17d20:	data_out=16'h2e4;
17'h17d21:	data_out=16'h91;
17'h17d22:	data_out=16'h183;
17'h17d23:	data_out=16'hae;
17'h17d24:	data_out=16'hab;
17'h17d25:	data_out=16'h16b;
17'h17d26:	data_out=16'hf8;
17'h17d27:	data_out=16'h2db;
17'h17d28:	data_out=16'h9a;
17'h17d29:	data_out=16'h1ef;
17'h17d2a:	data_out=16'h1ca;
17'h17d2b:	data_out=16'h19d;
17'h17d2c:	data_out=16'h1e7;
17'h17d2d:	data_out=16'h143;
17'h17d2e:	data_out=16'h189;
17'h17d2f:	data_out=16'h2e8;
17'h17d30:	data_out=16'h287;
17'h17d31:	data_out=16'h1e2;
17'h17d32:	data_out=16'h297;
17'h17d33:	data_out=16'h1cc;
17'h17d34:	data_out=16'h1de;
17'h17d35:	data_out=16'h2a9;
17'h17d36:	data_out=16'h1f3;
17'h17d37:	data_out=16'h1be;
17'h17d38:	data_out=16'h21f;
17'h17d39:	data_out=16'h1c2;
17'h17d3a:	data_out=16'h166;
17'h17d3b:	data_out=16'h1d6;
17'h17d3c:	data_out=16'h1d9;
17'h17d3d:	data_out=16'h278;
17'h17d3e:	data_out=16'ha1;
17'h17d3f:	data_out=16'h2b8;
17'h17d40:	data_out=16'h248;
17'h17d41:	data_out=16'h1d3;
17'h17d42:	data_out=16'h16a;
17'h17d43:	data_out=16'h13f;
17'h17d44:	data_out=16'h218;
17'h17d45:	data_out=16'h12f;
17'h17d46:	data_out=16'h178;
17'h17d47:	data_out=16'h18c;
17'h17d48:	data_out=16'h17e;
17'h17d49:	data_out=16'h170;
17'h17d4a:	data_out=16'h27a;
17'h17d4b:	data_out=16'h1fd;
17'h17d4c:	data_out=16'h1ba;
17'h17d4d:	data_out=16'h197;
17'h17d4e:	data_out=16'h286;
17'h17d4f:	data_out=16'h1b2;
17'h17d50:	data_out=16'h1f8;
17'h17d51:	data_out=16'h1e6;
17'h17d52:	data_out=16'hc9;
17'h17d53:	data_out=16'h321;
17'h17d54:	data_out=16'h2fb;
17'h17d55:	data_out=16'h13c;
17'h17d56:	data_out=16'h15e;
17'h17d57:	data_out=16'hd8;
17'h17d58:	data_out=16'h128;
17'h17d59:	data_out=16'h1e7;
17'h17d5a:	data_out=16'he4;
17'h17d5b:	data_out=16'h264;
17'h17d5c:	data_out=16'h23e;
17'h17d5d:	data_out=16'h24e;
17'h17d5e:	data_out=16'h2de;
17'h17d5f:	data_out=16'h13c;
17'h17d60:	data_out=16'h136;
17'h17d61:	data_out=16'h29b;
17'h17d62:	data_out=16'h18e;
17'h17d63:	data_out=16'h1d2;
17'h17d64:	data_out=16'h19b;
17'h17d65:	data_out=16'h1f3;
17'h17d66:	data_out=16'h11b;
17'h17d67:	data_out=16'h1bf;
17'h17d68:	data_out=16'h95;
17'h17d69:	data_out=16'h158;
17'h17d6a:	data_out=16'h93;
17'h17d6b:	data_out=16'h2bc;
17'h17d6c:	data_out=16'h19b;
17'h17d6d:	data_out=16'h1d5;
17'h17d6e:	data_out=16'h8a;
17'h17d6f:	data_out=16'h2e6;
17'h17d70:	data_out=16'h8c;
17'h17d71:	data_out=16'h15f;
17'h17d72:	data_out=16'h233;
17'h17d73:	data_out=16'h2e0;
17'h17d74:	data_out=16'h285;
17'h17d75:	data_out=16'h22e;
17'h17d76:	data_out=16'h148;
17'h17d77:	data_out=16'h21d;
17'h17d78:	data_out=16'h18f;
17'h17d79:	data_out=16'h1c3;
17'h17d7a:	data_out=16'h1c6;
17'h17d7b:	data_out=16'h9f;
17'h17d7c:	data_out=16'hd7;
17'h17d7d:	data_out=16'h19c;
17'h17d7e:	data_out=16'h130;
17'h17d7f:	data_out=16'h1e1;
17'h17d80:	data_out=16'h251;
17'h17d81:	data_out=16'h274;
17'h17d82:	data_out=16'h2b8;
17'h17d83:	data_out=16'h47b;
17'h17d84:	data_out=16'h21e;
17'h17d85:	data_out=16'h2cb;
17'h17d86:	data_out=16'h202;
17'h17d87:	data_out=16'hb1;
17'h17d88:	data_out=16'h288;
17'h17d89:	data_out=16'h13e;
17'h17d8a:	data_out=16'h16e;
17'h17d8b:	data_out=16'h291;
17'h17d8c:	data_out=16'h2b9;
17'h17d8d:	data_out=16'h2a5;
17'h17d8e:	data_out=16'hf8;
17'h17d8f:	data_out=16'h2f1;
17'h17d90:	data_out=16'h2d7;
17'h17d91:	data_out=16'h245;
17'h17d92:	data_out=16'h1d8;
17'h17d93:	data_out=16'h3c7;
17'h17d94:	data_out=16'h2d0;
17'h17d95:	data_out=16'h17c;
17'h17d96:	data_out=16'h259;
17'h17d97:	data_out=16'h335;
17'h17d98:	data_out=16'hb7;
17'h17d99:	data_out=16'h1a3;
17'h17d9a:	data_out=16'h26b;
17'h17d9b:	data_out=16'h309;
17'h17d9c:	data_out=16'h425;
17'h17d9d:	data_out=16'h31c;
17'h17d9e:	data_out=16'h279;
17'h17d9f:	data_out=16'h17e;
17'h17da0:	data_out=16'h352;
17'h17da1:	data_out=16'hf6;
17'h17da2:	data_out=16'h2a6;
17'h17da3:	data_out=16'h97;
17'h17da4:	data_out=16'h97;
17'h17da5:	data_out=16'h1cd;
17'h17da6:	data_out=16'h16a;
17'h17da7:	data_out=16'h366;
17'h17da8:	data_out=16'h111;
17'h17da9:	data_out=16'h366;
17'h17daa:	data_out=16'h275;
17'h17dab:	data_out=16'h31b;
17'h17dac:	data_out=16'h223;
17'h17dad:	data_out=16'h2a5;
17'h17dae:	data_out=16'h265;
17'h17daf:	data_out=16'h419;
17'h17db0:	data_out=16'h28d;
17'h17db1:	data_out=16'h117;
17'h17db2:	data_out=16'h2aa;
17'h17db3:	data_out=16'h29d;
17'h17db4:	data_out=16'h21b;
17'h17db5:	data_out=16'h2b1;
17'h17db6:	data_out=16'h305;
17'h17db7:	data_out=16'h2be;
17'h17db8:	data_out=16'h298;
17'h17db9:	data_out=16'h28b;
17'h17dba:	data_out=16'h1b0;
17'h17dbb:	data_out=16'h111;
17'h17dbc:	data_out=16'h429;
17'h17dbd:	data_out=16'h313;
17'h17dbe:	data_out=16'h111;
17'h17dbf:	data_out=16'h2ca;
17'h17dc0:	data_out=16'h22b;
17'h17dc1:	data_out=16'h35e;
17'h17dc2:	data_out=16'h1ec;
17'h17dc3:	data_out=16'h20a;
17'h17dc4:	data_out=16'h1a4;
17'h17dc5:	data_out=16'h185;
17'h17dc6:	data_out=16'h3c3;
17'h17dc7:	data_out=16'h22f;
17'h17dc8:	data_out=16'h242;
17'h17dc9:	data_out=16'h1d8;
17'h17dca:	data_out=16'h1d0;
17'h17dcb:	data_out=16'h2b7;
17'h17dcc:	data_out=16'h1ec;
17'h17dcd:	data_out=16'h2ba;
17'h17dce:	data_out=16'h2d6;
17'h17dcf:	data_out=16'h1c5;
17'h17dd0:	data_out=16'h30e;
17'h17dd1:	data_out=16'h33a;
17'h17dd2:	data_out=16'h79;
17'h17dd3:	data_out=16'h3f1;
17'h17dd4:	data_out=16'h3fb;
17'h17dd5:	data_out=16'h3c6;
17'h17dd6:	data_out=16'h157;
17'h17dd7:	data_out=16'h105;
17'h17dd8:	data_out=16'h3bd;
17'h17dd9:	data_out=16'h1d9;
17'h17dda:	data_out=16'h26d;
17'h17ddb:	data_out=16'h23e;
17'h17ddc:	data_out=16'h2bc;
17'h17ddd:	data_out=16'h2f8;
17'h17dde:	data_out=16'h41b;
17'h17ddf:	data_out=16'h150;
17'h17de0:	data_out=16'h14f;
17'h17de1:	data_out=16'h2a5;
17'h17de2:	data_out=16'h265;
17'h17de3:	data_out=16'h2b1;
17'h17de4:	data_out=16'h1cb;
17'h17de5:	data_out=16'h234;
17'h17de6:	data_out=16'h122;
17'h17de7:	data_out=16'h2dd;
17'h17de8:	data_out=16'h10a;
17'h17de9:	data_out=16'h20a;
17'h17dea:	data_out=16'hef;
17'h17deb:	data_out=16'h2c4;
17'h17dec:	data_out=16'h1b2;
17'h17ded:	data_out=16'h2ae;
17'h17dee:	data_out=16'hea;
17'h17def:	data_out=16'h388;
17'h17df0:	data_out=16'hf0;
17'h17df1:	data_out=16'hdb;
17'h17df2:	data_out=16'h2cc;
17'h17df3:	data_out=16'h35a;
17'h17df4:	data_out=16'h287;
17'h17df5:	data_out=16'h310;
17'h17df6:	data_out=16'h19c;
17'h17df7:	data_out=16'h3ce;
17'h17df8:	data_out=16'h22a;
17'h17df9:	data_out=16'h1f9;
17'h17dfa:	data_out=16'h2cd;
17'h17dfb:	data_out=16'h10b;
17'h17dfc:	data_out=16'hb7;
17'h17dfd:	data_out=16'h102;
17'h17dfe:	data_out=16'h21b;
17'h17dff:	data_out=16'h182;
17'h17e00:	data_out=16'h3da;
17'h17e01:	data_out=16'h4fc;
17'h17e02:	data_out=16'h39b;
17'h17e03:	data_out=16'h6d8;
17'h17e04:	data_out=16'h4d1;
17'h17e05:	data_out=16'h5fb;
17'h17e06:	data_out=16'h2ac;
17'h17e07:	data_out=16'h1a9;
17'h17e08:	data_out=16'h311;
17'h17e09:	data_out=16'h107;
17'h17e0a:	data_out=16'h3c3;
17'h17e0b:	data_out=16'h2ff;
17'h17e0c:	data_out=16'h415;
17'h17e0d:	data_out=16'h392;
17'h17e0e:	data_out=16'h125;
17'h17e0f:	data_out=16'h3df;
17'h17e10:	data_out=16'h334;
17'h17e11:	data_out=16'h4e7;
17'h17e12:	data_out=16'h23d;
17'h17e13:	data_out=16'h5af;
17'h17e14:	data_out=16'h3b0;
17'h17e15:	data_out=16'h220;
17'h17e16:	data_out=16'h3e0;
17'h17e17:	data_out=16'h45a;
17'h17e18:	data_out=16'h63;
17'h17e19:	data_out=16'h2fa;
17'h17e1a:	data_out=16'h568;
17'h17e1b:	data_out=16'h495;
17'h17e1c:	data_out=16'h728;
17'h17e1d:	data_out=16'h63b;
17'h17e1e:	data_out=16'h3de;
17'h17e1f:	data_out=16'h23c;
17'h17e20:	data_out=16'h6cc;
17'h17e21:	data_out=16'h135;
17'h17e22:	data_out=16'h3a8;
17'h17e23:	data_out=16'h45;
17'h17e24:	data_out=16'h45;
17'h17e25:	data_out=16'h26a;
17'h17e26:	data_out=16'h12b;
17'h17e27:	data_out=16'h681;
17'h17e28:	data_out=16'h140;
17'h17e29:	data_out=16'h460;
17'h17e2a:	data_out=16'h2d9;
17'h17e2b:	data_out=16'h4bf;
17'h17e2c:	data_out=16'h37f;
17'h17e2d:	data_out=16'h350;
17'h17e2e:	data_out=16'h36b;
17'h17e2f:	data_out=16'h720;
17'h17e30:	data_out=16'h569;
17'h17e31:	data_out=16'h3c2;
17'h17e32:	data_out=16'h5b0;
17'h17e33:	data_out=16'h386;
17'h17e34:	data_out=16'h3cb;
17'h17e35:	data_out=16'h576;
17'h17e36:	data_out=16'h3be;
17'h17e37:	data_out=16'h3a7;
17'h17e38:	data_out=16'h4d2;
17'h17e39:	data_out=16'h382;
17'h17e3a:	data_out=16'h221;
17'h17e3b:	data_out=16'h2c3;
17'h17e3c:	data_out=16'h60a;
17'h17e3d:	data_out=16'h57b;
17'h17e3e:	data_out=16'h140;
17'h17e3f:	data_out=16'h5f9;
17'h17e40:	data_out=16'h483;
17'h17e41:	data_out=16'h3fe;
17'h17e42:	data_out=16'h289;
17'h17e43:	data_out=16'h2b2;
17'h17e44:	data_out=16'h3b3;
17'h17e45:	data_out=16'h1bd;
17'h17e46:	data_out=16'h45d;
17'h17e47:	data_out=16'h271;
17'h17e48:	data_out=16'h309;
17'h17e49:	data_out=16'h274;
17'h17e4a:	data_out=16'h33c;
17'h17e4b:	data_out=16'h3fc;
17'h17e4c:	data_out=16'h29a;
17'h17e4d:	data_out=16'h3c6;
17'h17e4e:	data_out=16'h425;
17'h17e4f:	data_out=16'h261;
17'h17e50:	data_out=16'h483;
17'h17e51:	data_out=16'h44c;
17'h17e52:	data_out=16'h37;
17'h17e53:	data_out=16'h745;
17'h17e54:	data_out=16'h715;
17'h17e55:	data_out=16'h43b;
17'h17e56:	data_out=16'h1c7;
17'h17e57:	data_out=16'h193;
17'h17e58:	data_out=16'h46a;
17'h17e59:	data_out=16'h3b7;
17'h17e5a:	data_out=16'h473;
17'h17e5b:	data_out=16'h4f5;
17'h17e5c:	data_out=16'h586;
17'h17e5d:	data_out=16'h56f;
17'h17e5e:	data_out=16'h723;
17'h17e5f:	data_out=16'h1e7;
17'h17e60:	data_out=16'h16a;
17'h17e61:	data_out=16'h599;
17'h17e62:	data_out=16'h2e1;
17'h17e63:	data_out=16'h3a3;
17'h17e64:	data_out=16'h2d0;
17'h17e65:	data_out=16'h4b6;
17'h17e66:	data_out=16'h214;
17'h17e67:	data_out=16'h321;
17'h17e68:	data_out=16'h137;
17'h17e69:	data_out=16'h281;
17'h17e6a:	data_out=16'h122;
17'h17e6b:	data_out=16'h5fe;
17'h17e6c:	data_out=16'h409;
17'h17e6d:	data_out=16'h3a7;
17'h17e6e:	data_out=16'h111;
17'h17e6f:	data_out=16'h6ff;
17'h17e70:	data_out=16'h129;
17'h17e71:	data_out=16'h113;
17'h17e72:	data_out=16'h602;
17'h17e73:	data_out=16'h6ba;
17'h17e74:	data_out=16'h55e;
17'h17e75:	data_out=16'h57a;
17'h17e76:	data_out=16'h1e0;
17'h17e77:	data_out=16'h4c2;
17'h17e78:	data_out=16'h33a;
17'h17e79:	data_out=16'h314;
17'h17e7a:	data_out=16'h3b6;
17'h17e7b:	data_out=16'h140;
17'h17e7c:	data_out=16'ha8;
17'h17e7d:	data_out=16'h16e;
17'h17e7e:	data_out=16'h289;
17'h17e7f:	data_out=16'h2e7;
17'h17e80:	data_out=16'h538;
17'h17e81:	data_out=16'h779;
17'h17e82:	data_out=16'h4fa;
17'h17e83:	data_out=16'h8ea;
17'h17e84:	data_out=16'h8f7;
17'h17e85:	data_out=16'ha00;
17'h17e86:	data_out=16'h3d9;
17'h17e87:	data_out=16'h4ab;
17'h17e88:	data_out=16'h388;
17'h17e89:	data_out=16'h14d;
17'h17e8a:	data_out=16'h67f;
17'h17e8b:	data_out=16'h2c2;
17'h17e8c:	data_out=16'h5c2;
17'h17e8d:	data_out=16'h503;
17'h17e8e:	data_out=16'h17e;
17'h17e8f:	data_out=16'h58b;
17'h17e90:	data_out=16'h3a6;
17'h17e91:	data_out=16'h866;
17'h17e92:	data_out=16'h359;
17'h17e93:	data_out=16'h7b2;
17'h17e94:	data_out=16'h47c;
17'h17e95:	data_out=16'h32c;
17'h17e96:	data_out=16'h623;
17'h17e97:	data_out=16'h515;
17'h17e98:	data_out=16'he9;
17'h17e99:	data_out=16'h36f;
17'h17e9a:	data_out=16'h9ad;
17'h17e9b:	data_out=16'h59e;
17'h17e9c:	data_out=16'ha00;
17'h17e9d:	data_out=16'h998;
17'h17e9e:	data_out=16'h5d4;
17'h17e9f:	data_out=16'h462;
17'h17ea0:	data_out=16'ha00;
17'h17ea1:	data_out=16'h17f;
17'h17ea2:	data_out=16'h4b0;
17'h17ea3:	data_out=16'h4a;
17'h17ea4:	data_out=16'h4a;
17'h17ea5:	data_out=16'h39b;
17'h17ea6:	data_out=16'h1aa;
17'h17ea7:	data_out=16'h9ec;
17'h17ea8:	data_out=16'h18b;
17'h17ea9:	data_out=16'h515;
17'h17eaa:	data_out=16'h3d5;
17'h17eab:	data_out=16'h519;
17'h17eac:	data_out=16'h589;
17'h17ead:	data_out=16'h308;
17'h17eae:	data_out=16'h53a;
17'h17eaf:	data_out=16'ha00;
17'h17eb0:	data_out=16'h95b;
17'h17eb1:	data_out=16'h6ed;
17'h17eb2:	data_out=16'h9c8;
17'h17eb3:	data_out=16'h4a0;
17'h17eb4:	data_out=16'h537;
17'h17eb5:	data_out=16'h971;
17'h17eb6:	data_out=16'h442;
17'h17eb7:	data_out=16'h4f4;
17'h17eb8:	data_out=16'h8c0;
17'h17eb9:	data_out=16'h4c4;
17'h17eba:	data_out=16'h2f7;
17'h17ebb:	data_out=16'h56e;
17'h17ebc:	data_out=16'h6e7;
17'h17ebd:	data_out=16'h8e5;
17'h17ebe:	data_out=16'h18c;
17'h17ebf:	data_out=16'ha00;
17'h17ec0:	data_out=16'h864;
17'h17ec1:	data_out=16'h402;
17'h17ec2:	data_out=16'h340;
17'h17ec3:	data_out=16'h39d;
17'h17ec4:	data_out=16'h6bd;
17'h17ec5:	data_out=16'h34e;
17'h17ec6:	data_out=16'h336;
17'h17ec7:	data_out=16'h352;
17'h17ec8:	data_out=16'h3e8;
17'h17ec9:	data_out=16'h3b6;
17'h17eca:	data_out=16'h62d;
17'h17ecb:	data_out=16'h532;
17'h17ecc:	data_out=16'h3e8;
17'h17ecd:	data_out=16'h4cf;
17'h17ece:	data_out=16'h61e;
17'h17ecf:	data_out=16'h3a2;
17'h17ed0:	data_out=16'h697;
17'h17ed1:	data_out=16'h5f0;
17'h17ed2:	data_out=16'h67;
17'h17ed3:	data_out=16'ha00;
17'h17ed4:	data_out=16'ha00;
17'h17ed5:	data_out=16'h41c;
17'h17ed6:	data_out=16'h389;
17'h17ed7:	data_out=16'h33d;
17'h17ed8:	data_out=16'h47c;
17'h17ed9:	data_out=16'h73f;
17'h17eda:	data_out=16'h57e;
17'h17edb:	data_out=16'h8b4;
17'h17edc:	data_out=16'h894;
17'h17edd:	data_out=16'h891;
17'h17ede:	data_out=16'ha00;
17'h17edf:	data_out=16'h2ce;
17'h17ee0:	data_out=16'h1ac;
17'h17ee1:	data_out=16'h9a5;
17'h17ee2:	data_out=16'h368;
17'h17ee3:	data_out=16'h4ae;
17'h17ee4:	data_out=16'h401;
17'h17ee5:	data_out=16'h7cb;
17'h17ee6:	data_out=16'h2c7;
17'h17ee7:	data_out=16'h341;
17'h17ee8:	data_out=16'h181;
17'h17ee9:	data_out=16'h303;
17'h17eea:	data_out=16'h17c;
17'h17eeb:	data_out=16'ha00;
17'h17eec:	data_out=16'h6e3;
17'h17eed:	data_out=16'h4c0;
17'h17eee:	data_out=16'h17c;
17'h17eef:	data_out=16'ha00;
17'h17ef0:	data_out=16'h17d;
17'h17ef1:	data_out=16'h32f;
17'h17ef2:	data_out=16'ha00;
17'h17ef3:	data_out=16'ha00;
17'h17ef4:	data_out=16'h951;
17'h17ef5:	data_out=16'h832;
17'h17ef6:	data_out=16'h200;
17'h17ef7:	data_out=16'h605;
17'h17ef8:	data_out=16'h486;
17'h17ef9:	data_out=16'h5db;
17'h17efa:	data_out=16'h49e;
17'h17efb:	data_out=16'h18c;
17'h17efc:	data_out=16'h153;
17'h17efd:	data_out=16'h36e;
17'h17efe:	data_out=16'h324;
17'h17eff:	data_out=16'h61f;
17'h17f00:	data_out=16'h697;
17'h17f01:	data_out=16'h808;
17'h17f02:	data_out=16'h60f;
17'h17f03:	data_out=16'ha00;
17'h17f04:	data_out=16'ha00;
17'h17f05:	data_out=16'ha00;
17'h17f06:	data_out=16'h4b9;
17'h17f07:	data_out=16'h5cc;
17'h17f08:	data_out=16'h4fd;
17'h17f09:	data_out=16'h234;
17'h17f0a:	data_out=16'h79f;
17'h17f0b:	data_out=16'h2b9;
17'h17f0c:	data_out=16'h723;
17'h17f0d:	data_out=16'h67d;
17'h17f0e:	data_out=16'h1c0;
17'h17f0f:	data_out=16'h656;
17'h17f10:	data_out=16'h5d3;
17'h17f11:	data_out=16'ha00;
17'h17f12:	data_out=16'h44d;
17'h17f13:	data_out=16'h9b0;
17'h17f14:	data_out=16'h51b;
17'h17f15:	data_out=16'h403;
17'h17f16:	data_out=16'h7e6;
17'h17f17:	data_out=16'h583;
17'h17f18:	data_out=16'h141;
17'h17f19:	data_out=16'h2b4;
17'h17f1a:	data_out=16'ha00;
17'h17f1b:	data_out=16'h5be;
17'h17f1c:	data_out=16'ha00;
17'h17f1d:	data_out=16'ha00;
17'h17f1e:	data_out=16'h6b1;
17'h17f1f:	data_out=16'h5e1;
17'h17f20:	data_out=16'ha00;
17'h17f21:	data_out=16'h1c1;
17'h17f22:	data_out=16'h590;
17'h17f23:	data_out=16'he5;
17'h17f24:	data_out=16'he5;
17'h17f25:	data_out=16'h521;
17'h17f26:	data_out=16'h378;
17'h17f27:	data_out=16'ha00;
17'h17f28:	data_out=16'h1cf;
17'h17f29:	data_out=16'h6e3;
17'h17f2a:	data_out=16'h46f;
17'h17f2b:	data_out=16'h52f;
17'h17f2c:	data_out=16'h71c;
17'h17f2d:	data_out=16'h427;
17'h17f2e:	data_out=16'h5c6;
17'h17f2f:	data_out=16'ha00;
17'h17f30:	data_out=16'ha00;
17'h17f31:	data_out=16'h7ac;
17'h17f32:	data_out=16'ha00;
17'h17f33:	data_out=16'h54b;
17'h17f34:	data_out=16'h674;
17'h17f35:	data_out=16'ha00;
17'h17f36:	data_out=16'h592;
17'h17f37:	data_out=16'h5f4;
17'h17f38:	data_out=16'ha00;
17'h17f39:	data_out=16'h579;
17'h17f3a:	data_out=16'h2ca;
17'h17f3b:	data_out=16'h6f6;
17'h17f3c:	data_out=16'h79a;
17'h17f3d:	data_out=16'ha00;
17'h17f3e:	data_out=16'h1d0;
17'h17f3f:	data_out=16'ha00;
17'h17f40:	data_out=16'ha00;
17'h17f41:	data_out=16'h55d;
17'h17f42:	data_out=16'h4d8;
17'h17f43:	data_out=16'h432;
17'h17f44:	data_out=16'h84e;
17'h17f45:	data_out=16'h432;
17'h17f46:	data_out=16'h4a7;
17'h17f47:	data_out=16'h48f;
17'h17f48:	data_out=16'h387;
17'h17f49:	data_out=16'h564;
17'h17f4a:	data_out=16'h740;
17'h17f4b:	data_out=16'h66a;
17'h17f4c:	data_out=16'h51a;
17'h17f4d:	data_out=16'h5a0;
17'h17f4e:	data_out=16'h6c3;
17'h17f4f:	data_out=16'h47f;
17'h17f50:	data_out=16'h86d;
17'h17f51:	data_out=16'h876;
17'h17f52:	data_out=16'he2;
17'h17f53:	data_out=16'ha00;
17'h17f54:	data_out=16'ha00;
17'h17f55:	data_out=16'h605;
17'h17f56:	data_out=16'h54e;
17'h17f57:	data_out=16'h4d3;
17'h17f58:	data_out=16'h6c0;
17'h17f59:	data_out=16'h94d;
17'h17f5a:	data_out=16'h548;
17'h17f5b:	data_out=16'ha00;
17'h17f5c:	data_out=16'h972;
17'h17f5d:	data_out=16'h966;
17'h17f5e:	data_out=16'ha00;
17'h17f5f:	data_out=16'h318;
17'h17f60:	data_out=16'h2e5;
17'h17f61:	data_out=16'ha00;
17'h17f62:	data_out=16'h3c3;
17'h17f63:	data_out=16'h53f;
17'h17f64:	data_out=16'h506;
17'h17f65:	data_out=16'h8e6;
17'h17f66:	data_out=16'h261;
17'h17f67:	data_out=16'h32b;
17'h17f68:	data_out=16'h1c4;
17'h17f69:	data_out=16'h487;
17'h17f6a:	data_out=16'h1be;
17'h17f6b:	data_out=16'ha00;
17'h17f6c:	data_out=16'h7c2;
17'h17f6d:	data_out=16'h559;
17'h17f6e:	data_out=16'h1be;
17'h17f6f:	data_out=16'ha00;
17'h17f70:	data_out=16'h1bf;
17'h17f71:	data_out=16'h375;
17'h17f72:	data_out=16'ha00;
17'h17f73:	data_out=16'ha00;
17'h17f74:	data_out=16'ha00;
17'h17f75:	data_out=16'h934;
17'h17f76:	data_out=16'h244;
17'h17f77:	data_out=16'h89d;
17'h17f78:	data_out=16'h514;
17'h17f79:	data_out=16'h6cc;
17'h17f7a:	data_out=16'h531;
17'h17f7b:	data_out=16'h1d0;
17'h17f7c:	data_out=16'h1a6;
17'h17f7d:	data_out=16'h41d;
17'h17f7e:	data_out=16'h511;
17'h17f7f:	data_out=16'h76f;
17'h17f80:	data_out=16'h819;
17'h17f81:	data_out=16'h80d;
17'h17f82:	data_out=16'h5dc;
17'h17f83:	data_out=16'ha00;
17'h17f84:	data_out=16'h9f2;
17'h17f85:	data_out=16'ha00;
17'h17f86:	data_out=16'h4e3;
17'h17f87:	data_out=16'h622;
17'h17f88:	data_out=16'h55d;
17'h17f89:	data_out=16'h2e2;
17'h17f8a:	data_out=16'h6df;
17'h17f8b:	data_out=16'h289;
17'h17f8c:	data_out=16'h6f2;
17'h17f8d:	data_out=16'h67d;
17'h17f8e:	data_out=16'h1c7;
17'h17f8f:	data_out=16'h605;
17'h17f90:	data_out=16'h66e;
17'h17f91:	data_out=16'h913;
17'h17f92:	data_out=16'h492;
17'h17f93:	data_out=16'h998;
17'h17f94:	data_out=16'h536;
17'h17f95:	data_out=16'h421;
17'h17f96:	data_out=16'h80d;
17'h17f97:	data_out=16'h590;
17'h17f98:	data_out=16'h1b7;
17'h17f99:	data_out=16'h15a;
17'h17f9a:	data_out=16'h9e9;
17'h17f9b:	data_out=16'h54b;
17'h17f9c:	data_out=16'ha00;
17'h17f9d:	data_out=16'ha00;
17'h17f9e:	data_out=16'h6ad;
17'h17f9f:	data_out=16'h4ac;
17'h17fa0:	data_out=16'ha00;
17'h17fa1:	data_out=16'h1c7;
17'h17fa2:	data_out=16'h52b;
17'h17fa3:	data_out=16'h129;
17'h17fa4:	data_out=16'h129;
17'h17fa5:	data_out=16'h508;
17'h17fa6:	data_out=16'h3ff;
17'h17fa7:	data_out=16'ha00;
17'h17fa8:	data_out=16'h1d2;
17'h17fa9:	data_out=16'h77e;
17'h17faa:	data_out=16'h56b;
17'h17fab:	data_out=16'h425;
17'h17fac:	data_out=16'h72e;
17'h17fad:	data_out=16'h3ce;
17'h17fae:	data_out=16'h626;
17'h17faf:	data_out=16'ha00;
17'h17fb0:	data_out=16'ha00;
17'h17fb1:	data_out=16'h630;
17'h17fb2:	data_out=16'ha00;
17'h17fb3:	data_out=16'h558;
17'h17fb4:	data_out=16'h73a;
17'h17fb5:	data_out=16'ha00;
17'h17fb6:	data_out=16'h708;
17'h17fb7:	data_out=16'h599;
17'h17fb8:	data_out=16'ha00;
17'h17fb9:	data_out=16'h5ac;
17'h17fba:	data_out=16'h350;
17'h17fbb:	data_out=16'h6fc;
17'h17fbc:	data_out=16'h707;
17'h17fbd:	data_out=16'ha00;
17'h17fbe:	data_out=16'h1d3;
17'h17fbf:	data_out=16'ha00;
17'h17fc0:	data_out=16'h9e5;
17'h17fc1:	data_out=16'h624;
17'h17fc2:	data_out=16'h542;
17'h17fc3:	data_out=16'h313;
17'h17fc4:	data_out=16'h806;
17'h17fc5:	data_out=16'h450;
17'h17fc6:	data_out=16'h46a;
17'h17fc7:	data_out=16'h599;
17'h17fc8:	data_out=16'h2f9;
17'h17fc9:	data_out=16'h552;
17'h17fca:	data_out=16'h83c;
17'h17fcb:	data_out=16'h64c;
17'h17fcc:	data_out=16'h5d7;
17'h17fcd:	data_out=16'h578;
17'h17fce:	data_out=16'h717;
17'h17fcf:	data_out=16'h54d;
17'h17fd0:	data_out=16'h889;
17'h17fd1:	data_out=16'h7f1;
17'h17fd2:	data_out=16'h106;
17'h17fd3:	data_out=16'ha00;
17'h17fd4:	data_out=16'ha00;
17'h17fd5:	data_out=16'h581;
17'h17fd6:	data_out=16'h576;
17'h17fd7:	data_out=16'h48b;
17'h17fd8:	data_out=16'h69a;
17'h17fd9:	data_out=16'h919;
17'h17fda:	data_out=16'h3d3;
17'h17fdb:	data_out=16'h97c;
17'h17fdc:	data_out=16'h904;
17'h17fdd:	data_out=16'h9bb;
17'h17fde:	data_out=16'ha00;
17'h17fdf:	data_out=16'h384;
17'h17fe0:	data_out=16'h390;
17'h17fe1:	data_out=16'ha00;
17'h17fe2:	data_out=16'h345;
17'h17fe3:	data_out=16'h537;
17'h17fe4:	data_out=16'h602;
17'h17fe5:	data_out=16'h7e1;
17'h17fe6:	data_out=16'hef;
17'h17fe7:	data_out=16'h344;
17'h17fe8:	data_out=16'h1c8;
17'h17fe9:	data_out=16'h4c8;
17'h17fea:	data_out=16'h1c6;
17'h17feb:	data_out=16'ha00;
17'h17fec:	data_out=16'h8b5;
17'h17fed:	data_out=16'h559;
17'h17fee:	data_out=16'h1c6;
17'h17fef:	data_out=16'ha00;
17'h17ff0:	data_out=16'h1c7;
17'h17ff1:	data_out=16'h437;
17'h17ff2:	data_out=16'ha00;
17'h17ff3:	data_out=16'ha00;
17'h17ff4:	data_out=16'ha00;
17'h17ff5:	data_out=16'h7dc;
17'h17ff6:	data_out=16'h208;
17'h17ff7:	data_out=16'h943;
17'h17ff8:	data_out=16'h3f3;
17'h17ff9:	data_out=16'h7a9;
17'h17ffa:	data_out=16'h53a;
17'h17ffb:	data_out=16'h1d3;
17'h17ffc:	data_out=16'h20e;
17'h17ffd:	data_out=16'h2d6;
17'h17ffe:	data_out=16'h555;
17'h17fff:	data_out=16'h77b;
17'h18000:	data_out=16'h7b5;
17'h18001:	data_out=16'h692;
17'h18002:	data_out=16'h5fa;
17'h18003:	data_out=16'ha00;
17'h18004:	data_out=16'h82e;
17'h18005:	data_out=16'ha00;
17'h18006:	data_out=16'h63a;
17'h18007:	data_out=16'h502;
17'h18008:	data_out=16'h52c;
17'h18009:	data_out=16'h456;
17'h1800a:	data_out=16'h52c;
17'h1800b:	data_out=16'h5c2;
17'h1800c:	data_out=16'h4a8;
17'h1800d:	data_out=16'h774;
17'h1800e:	data_out=16'h1d6;
17'h1800f:	data_out=16'h5d1;
17'h18010:	data_out=16'h862;
17'h18011:	data_out=16'h736;
17'h18012:	data_out=16'h592;
17'h18013:	data_out=16'ha00;
17'h18014:	data_out=16'h75c;
17'h18015:	data_out=16'h3bd;
17'h18016:	data_out=16'h7ce;
17'h18017:	data_out=16'h800;
17'h18018:	data_out=16'hf2;
17'h18019:	data_out=16'h98;
17'h1801a:	data_out=16'h871;
17'h1801b:	data_out=16'h776;
17'h1801c:	data_out=16'ha00;
17'h1801d:	data_out=16'h9cc;
17'h1801e:	data_out=16'h7ea;
17'h1801f:	data_out=16'h3b3;
17'h18020:	data_out=16'ha00;
17'h18021:	data_out=16'h1d9;
17'h18022:	data_out=16'h792;
17'h18023:	data_out=16'h804c;
17'h18024:	data_out=16'h804d;
17'h18025:	data_out=16'h635;
17'h18026:	data_out=16'h552;
17'h18027:	data_out=16'ha00;
17'h18028:	data_out=16'h1ea;
17'h18029:	data_out=16'h8fb;
17'h1802a:	data_out=16'h50d;
17'h1802b:	data_out=16'h472;
17'h1802c:	data_out=16'h6db;
17'h1802d:	data_out=16'h555;
17'h1802e:	data_out=16'h640;
17'h1802f:	data_out=16'ha00;
17'h18030:	data_out=16'h8a0;
17'h18031:	data_out=16'h4a8;
17'h18032:	data_out=16'h8f3;
17'h18033:	data_out=16'h6f5;
17'h18034:	data_out=16'h655;
17'h18035:	data_out=16'h8df;
17'h18036:	data_out=16'h6fd;
17'h18037:	data_out=16'h5d4;
17'h18038:	data_out=16'ha00;
17'h18039:	data_out=16'h714;
17'h1803a:	data_out=16'h35a;
17'h1803b:	data_out=16'h50e;
17'h1803c:	data_out=16'h842;
17'h1803d:	data_out=16'ha00;
17'h1803e:	data_out=16'h1eb;
17'h1803f:	data_out=16'ha00;
17'h18040:	data_out=16'ha00;
17'h18041:	data_out=16'h6d2;
17'h18042:	data_out=16'h664;
17'h18043:	data_out=16'h505;
17'h18044:	data_out=16'h6c7;
17'h18045:	data_out=16'h3ed;
17'h18046:	data_out=16'h60e;
17'h18047:	data_out=16'h5ab;
17'h18048:	data_out=16'h3a2;
17'h18049:	data_out=16'h67c;
17'h1804a:	data_out=16'h663;
17'h1804b:	data_out=16'h550;
17'h1804c:	data_out=16'h616;
17'h1804d:	data_out=16'h7cc;
17'h1804e:	data_out=16'h6c2;
17'h1804f:	data_out=16'h52f;
17'h18050:	data_out=16'h9b3;
17'h18051:	data_out=16'h7eb;
17'h18052:	data_out=16'h8060;
17'h18053:	data_out=16'h8a2;
17'h18054:	data_out=16'ha00;
17'h18055:	data_out=16'h78e;
17'h18056:	data_out=16'h667;
17'h18057:	data_out=16'h5b5;
17'h18058:	data_out=16'h7c8;
17'h18059:	data_out=16'h9ce;
17'h1805a:	data_out=16'h556;
17'h1805b:	data_out=16'h6ee;
17'h1805c:	data_out=16'h7e7;
17'h1805d:	data_out=16'h956;
17'h1805e:	data_out=16'ha00;
17'h1805f:	data_out=16'h326;
17'h18060:	data_out=16'h420;
17'h18061:	data_out=16'h8d4;
17'h18062:	data_out=16'h518;
17'h18063:	data_out=16'h6d4;
17'h18064:	data_out=16'h5d7;
17'h18065:	data_out=16'h824;
17'h18066:	data_out=16'h45;
17'h18067:	data_out=16'h454;
17'h18068:	data_out=16'h1dc;
17'h18069:	data_out=16'h4e1;
17'h1806a:	data_out=16'h1d4;
17'h1806b:	data_out=16'h972;
17'h1806c:	data_out=16'h6f7;
17'h1806d:	data_out=16'h6f1;
17'h1806e:	data_out=16'h1d4;
17'h1806f:	data_out=16'ha00;
17'h18070:	data_out=16'h1d5;
17'h18071:	data_out=16'h298;
17'h18072:	data_out=16'ha00;
17'h18073:	data_out=16'ha00;
17'h18074:	data_out=16'h899;
17'h18075:	data_out=16'h915;
17'h18076:	data_out=16'h242;
17'h18077:	data_out=16'ha00;
17'h18078:	data_out=16'h5be;
17'h18079:	data_out=16'h745;
17'h1807a:	data_out=16'h715;
17'h1807b:	data_out=16'h1ec;
17'h1807c:	data_out=16'h128;
17'h1807d:	data_out=16'h332;
17'h1807e:	data_out=16'h831;
17'h1807f:	data_out=16'h636;
17'h18080:	data_out=16'ha00;
17'h18081:	data_out=16'ha00;
17'h18082:	data_out=16'h6a8;
17'h18083:	data_out=16'ha00;
17'h18084:	data_out=16'h77d;
17'h18085:	data_out=16'h9ff;
17'h18086:	data_out=16'h24b;
17'h18087:	data_out=16'h65c;
17'h18088:	data_out=16'h67b;
17'h18089:	data_out=16'h3a1;
17'h1808a:	data_out=16'h6eb;
17'h1808b:	data_out=16'h5eb;
17'h1808c:	data_out=16'h4c3;
17'h1808d:	data_out=16'h9d4;
17'h1808e:	data_out=16'h146;
17'h1808f:	data_out=16'h816;
17'h18090:	data_out=16'ha00;
17'h18091:	data_out=16'h733;
17'h18092:	data_out=16'h90c;
17'h18093:	data_out=16'ha00;
17'h18094:	data_out=16'h8e5;
17'h18095:	data_out=16'h335;
17'h18096:	data_out=16'h83e;
17'h18097:	data_out=16'ha00;
17'h18098:	data_out=16'h5d;
17'h18099:	data_out=16'h1a2;
17'h1809a:	data_out=16'h81c;
17'h1809b:	data_out=16'ha00;
17'h1809c:	data_out=16'ha00;
17'h1809d:	data_out=16'ha00;
17'h1809e:	data_out=16'ha00;
17'h1809f:	data_out=16'h105;
17'h180a0:	data_out=16'ha00;
17'h180a1:	data_out=16'h149;
17'h180a2:	data_out=16'ha00;
17'h180a3:	data_out=16'h8192;
17'h180a4:	data_out=16'h8195;
17'h180a5:	data_out=16'h6f3;
17'h180a6:	data_out=16'h3ad;
17'h180a7:	data_out=16'ha00;
17'h180a8:	data_out=16'h158;
17'h180a9:	data_out=16'ha00;
17'h180aa:	data_out=16'h985;
17'h180ab:	data_out=16'h6e2;
17'h180ac:	data_out=16'h6c6;
17'h180ad:	data_out=16'h7bc;
17'h180ae:	data_out=16'ha00;
17'h180af:	data_out=16'ha00;
17'h180b0:	data_out=16'h8d5;
17'h180b1:	data_out=16'h8c0;
17'h180b2:	data_out=16'h961;
17'h180b3:	data_out=16'h909;
17'h180b4:	data_out=16'h98e;
17'h180b5:	data_out=16'h7bb;
17'h180b6:	data_out=16'ha00;
17'h180b7:	data_out=16'h6a2;
17'h180b8:	data_out=16'ha00;
17'h180b9:	data_out=16'h9af;
17'h180ba:	data_out=16'h878;
17'h180bb:	data_out=16'h327;
17'h180bc:	data_out=16'ha00;
17'h180bd:	data_out=16'ha00;
17'h180be:	data_out=16'h159;
17'h180bf:	data_out=16'h9ff;
17'h180c0:	data_out=16'ha00;
17'h180c1:	data_out=16'h624;
17'h180c2:	data_out=16'ha00;
17'h180c3:	data_out=16'h8008;
17'h180c4:	data_out=16'h47a;
17'h180c5:	data_out=16'h369;
17'h180c6:	data_out=16'h76c;
17'h180c7:	data_out=16'h7d2;
17'h180c8:	data_out=16'h9f8;
17'h180c9:	data_out=16'h697;
17'h180ca:	data_out=16'h914;
17'h180cb:	data_out=16'ha00;
17'h180cc:	data_out=16'h9eb;
17'h180cd:	data_out=16'ha00;
17'h180ce:	data_out=16'ha00;
17'h180cf:	data_out=16'h86b;
17'h180d0:	data_out=16'h75a;
17'h180d1:	data_out=16'h363;
17'h180d2:	data_out=16'h81a0;
17'h180d3:	data_out=16'ha00;
17'h180d4:	data_out=16'ha00;
17'h180d5:	data_out=16'h407;
17'h180d6:	data_out=16'h39f;
17'h180d7:	data_out=16'h409;
17'h180d8:	data_out=16'h40c;
17'h180d9:	data_out=16'h8ea;
17'h180da:	data_out=16'ha00;
17'h180db:	data_out=16'h49f;
17'h180dc:	data_out=16'ha00;
17'h180dd:	data_out=16'ha00;
17'h180de:	data_out=16'ha00;
17'h180df:	data_out=16'h661;
17'h180e0:	data_out=16'h39d;
17'h180e1:	data_out=16'h797;
17'h180e2:	data_out=16'h6e7;
17'h180e3:	data_out=16'h906;
17'h180e4:	data_out=16'h649;
17'h180e5:	data_out=16'h9ff;
17'h180e6:	data_out=16'ha0;
17'h180e7:	data_out=16'h698;
17'h180e8:	data_out=16'h14c;
17'h180e9:	data_out=16'h5b0;
17'h180ea:	data_out=16'h142;
17'h180eb:	data_out=16'h974;
17'h180ec:	data_out=16'ha00;
17'h180ed:	data_out=16'h939;
17'h180ee:	data_out=16'h142;
17'h180ef:	data_out=16'ha00;
17'h180f0:	data_out=16'h144;
17'h180f1:	data_out=16'h431;
17'h180f2:	data_out=16'ha00;
17'h180f3:	data_out=16'ha00;
17'h180f4:	data_out=16'h8c9;
17'h180f5:	data_out=16'h5c0;
17'h180f6:	data_out=16'h230;
17'h180f7:	data_out=16'h830;
17'h180f8:	data_out=16'h19e;
17'h180f9:	data_out=16'ha00;
17'h180fa:	data_out=16'h8f9;
17'h180fb:	data_out=16'h15a;
17'h180fc:	data_out=16'h197;
17'h180fd:	data_out=16'h80d1;
17'h180fe:	data_out=16'h5cc;
17'h180ff:	data_out=16'h5c4;
17'h18100:	data_out=16'ha00;
17'h18101:	data_out=16'h9ff;
17'h18102:	data_out=16'h785;
17'h18103:	data_out=16'ha00;
17'h18104:	data_out=16'h8145;
17'h18105:	data_out=16'h262;
17'h18106:	data_out=16'h8165;
17'h18107:	data_out=16'h177;
17'h18108:	data_out=16'h89f;
17'h18109:	data_out=16'h506;
17'h1810a:	data_out=16'h171;
17'h1810b:	data_out=16'ha00;
17'h1810c:	data_out=16'h8044;
17'h1810d:	data_out=16'ha00;
17'h1810e:	data_out=16'hc5;
17'h1810f:	data_out=16'h917;
17'h18110:	data_out=16'ha00;
17'h18111:	data_out=16'h80eb;
17'h18112:	data_out=16'ha00;
17'h18113:	data_out=16'ha00;
17'h18114:	data_out=16'ha00;
17'h18115:	data_out=16'h12b;
17'h18116:	data_out=16'h55f;
17'h18117:	data_out=16'ha00;
17'h18118:	data_out=16'h0;
17'h18119:	data_out=16'h146;
17'h1811a:	data_out=16'h805a;
17'h1811b:	data_out=16'ha00;
17'h1811c:	data_out=16'h658;
17'h1811d:	data_out=16'ha00;
17'h1811e:	data_out=16'ha00;
17'h1811f:	data_out=16'h8556;
17'h18120:	data_out=16'ha00;
17'h18121:	data_out=16'hcc;
17'h18122:	data_out=16'ha00;
17'h18123:	data_out=16'h8307;
17'h18124:	data_out=16'h830a;
17'h18125:	data_out=16'h829;
17'h18126:	data_out=16'h664;
17'h18127:	data_out=16'h9ff;
17'h18128:	data_out=16'hde;
17'h18129:	data_out=16'ha00;
17'h1812a:	data_out=16'h9ff;
17'h1812b:	data_out=16'h621;
17'h1812c:	data_out=16'h3ab;
17'h1812d:	data_out=16'ha00;
17'h1812e:	data_out=16'ha00;
17'h1812f:	data_out=16'ha00;
17'h18130:	data_out=16'h177;
17'h18131:	data_out=16'h213;
17'h18132:	data_out=16'h18a;
17'h18133:	data_out=16'ha00;
17'h18134:	data_out=16'h703;
17'h18135:	data_out=16'h80e3;
17'h18136:	data_out=16'ha00;
17'h18137:	data_out=16'h7a7;
17'h18138:	data_out=16'h6c8;
17'h18139:	data_out=16'ha00;
17'h1813a:	data_out=16'h826;
17'h1813b:	data_out=16'h84b7;
17'h1813c:	data_out=16'ha00;
17'h1813d:	data_out=16'h994;
17'h1813e:	data_out=16'hdf;
17'h1813f:	data_out=16'h187;
17'h18140:	data_out=16'h58b;
17'h18141:	data_out=16'h950;
17'h18142:	data_out=16'ha00;
17'h18143:	data_out=16'h8441;
17'h18144:	data_out=16'h82c0;
17'h18145:	data_out=16'hfc;
17'h18146:	data_out=16'ha00;
17'h18147:	data_out=16'h7ac;
17'h18148:	data_out=16'ha00;
17'h18149:	data_out=16'h77e;
17'h1814a:	data_out=16'h525;
17'h1814b:	data_out=16'ha00;
17'h1814c:	data_out=16'ha00;
17'h1814d:	data_out=16'ha00;
17'h1814e:	data_out=16'ha00;
17'h1814f:	data_out=16'h7d4;
17'h18150:	data_out=16'h501;
17'h18151:	data_out=16'h8205;
17'h18152:	data_out=16'h837e;
17'h18153:	data_out=16'ha00;
17'h18154:	data_out=16'ha00;
17'h18155:	data_out=16'h5d7;
17'h18156:	data_out=16'h289;
17'h18157:	data_out=16'h2c6;
17'h18158:	data_out=16'h54b;
17'h18159:	data_out=16'h529;
17'h1815a:	data_out=16'ha00;
17'h1815b:	data_out=16'h86bc;
17'h1815c:	data_out=16'h870;
17'h1815d:	data_out=16'ha00;
17'h1815e:	data_out=16'ha00;
17'h1815f:	data_out=16'h73d;
17'h18160:	data_out=16'h490;
17'h18161:	data_out=16'h81b8;
17'h18162:	data_out=16'h980;
17'h18163:	data_out=16'ha00;
17'h18164:	data_out=16'h3f5;
17'h18165:	data_out=16'h6b6;
17'h18166:	data_out=16'h8016;
17'h18167:	data_out=16'h8a6;
17'h18168:	data_out=16'hd1;
17'h18169:	data_out=16'h854;
17'h1816a:	data_out=16'hbe;
17'h1816b:	data_out=16'h11f;
17'h1816c:	data_out=16'ha00;
17'h1816d:	data_out=16'ha00;
17'h1816e:	data_out=16'hbe;
17'h1816f:	data_out=16'h9a4;
17'h18170:	data_out=16'hc1;
17'h18171:	data_out=16'h1b2;
17'h18172:	data_out=16'h3f3;
17'h18173:	data_out=16'h49d;
17'h18174:	data_out=16'h166;
17'h18175:	data_out=16'h14f;
17'h18176:	data_out=16'h1ea;
17'h18177:	data_out=16'h8e9;
17'h18178:	data_out=16'h822a;
17'h18179:	data_out=16'ha00;
17'h1817a:	data_out=16'ha00;
17'h1817b:	data_out=16'he0;
17'h1817c:	data_out=16'h111;
17'h1817d:	data_out=16'h86ad;
17'h1817e:	data_out=16'h86c;
17'h1817f:	data_out=16'h801d;
17'h18180:	data_out=16'ha00;
17'h18181:	data_out=16'h9c4;
17'h18182:	data_out=16'h676;
17'h18183:	data_out=16'ha00;
17'h18184:	data_out=16'h281;
17'h18185:	data_out=16'h5a9;
17'h18186:	data_out=16'h343;
17'h18187:	data_out=16'h4b9;
17'h18188:	data_out=16'h628;
17'h18189:	data_out=16'h6b3;
17'h1818a:	data_out=16'h203;
17'h1818b:	data_out=16'h870;
17'h1818c:	data_out=16'hc6;
17'h1818d:	data_out=16'ha00;
17'h1818e:	data_out=16'h131;
17'h1818f:	data_out=16'h8ad;
17'h18190:	data_out=16'ha00;
17'h18191:	data_out=16'h193;
17'h18192:	data_out=16'ha00;
17'h18193:	data_out=16'ha00;
17'h18194:	data_out=16'ha00;
17'h18195:	data_out=16'h229;
17'h18196:	data_out=16'h667;
17'h18197:	data_out=16'ha00;
17'h18198:	data_out=16'hdc;
17'h18199:	data_out=16'haf;
17'h1819a:	data_out=16'h3c2;
17'h1819b:	data_out=16'ha00;
17'h1819c:	data_out=16'h7ec;
17'h1819d:	data_out=16'ha00;
17'h1819e:	data_out=16'ha00;
17'h1819f:	data_out=16'h8038;
17'h181a0:	data_out=16'ha00;
17'h181a1:	data_out=16'h136;
17'h181a2:	data_out=16'ha00;
17'h181a3:	data_out=16'h82c7;
17'h181a4:	data_out=16'h82cb;
17'h181a5:	data_out=16'h779;
17'h181a6:	data_out=16'h682;
17'h181a7:	data_out=16'ha00;
17'h181a8:	data_out=16'h146;
17'h181a9:	data_out=16'ha00;
17'h181aa:	data_out=16'ha00;
17'h181ab:	data_out=16'h3e1;
17'h181ac:	data_out=16'h4f6;
17'h181ad:	data_out=16'h9d4;
17'h181ae:	data_out=16'ha00;
17'h181af:	data_out=16'ha00;
17'h181b0:	data_out=16'h45b;
17'h181b1:	data_out=16'h326;
17'h181b2:	data_out=16'h46e;
17'h181b3:	data_out=16'ha00;
17'h181b4:	data_out=16'h7b8;
17'h181b5:	data_out=16'h135;
17'h181b6:	data_out=16'ha00;
17'h181b7:	data_out=16'h67b;
17'h181b8:	data_out=16'h6e8;
17'h181b9:	data_out=16'ha00;
17'h181ba:	data_out=16'h700;
17'h181bb:	data_out=16'h81de;
17'h181bc:	data_out=16'h9a9;
17'h181bd:	data_out=16'ha00;
17'h181be:	data_out=16'h146;
17'h181bf:	data_out=16'h5a4;
17'h181c0:	data_out=16'h83d;
17'h181c1:	data_out=16'h724;
17'h181c2:	data_out=16'ha00;
17'h181c3:	data_out=16'h72;
17'h181c4:	data_out=16'h151;
17'h181c5:	data_out=16'h253;
17'h181c6:	data_out=16'h7ed;
17'h181c7:	data_out=16'h87f;
17'h181c8:	data_out=16'ha00;
17'h181c9:	data_out=16'h6e9;
17'h181ca:	data_out=16'h760;
17'h181cb:	data_out=16'ha00;
17'h181cc:	data_out=16'h9d8;
17'h181cd:	data_out=16'ha00;
17'h181ce:	data_out=16'h9f9;
17'h181cf:	data_out=16'h7e2;
17'h181d0:	data_out=16'h726;
17'h181d1:	data_out=16'h9c;
17'h181d2:	data_out=16'h82e2;
17'h181d3:	data_out=16'ha00;
17'h181d4:	data_out=16'ha00;
17'h181d5:	data_out=16'h4c2;
17'h181d6:	data_out=16'h3d3;
17'h181d7:	data_out=16'h3cb;
17'h181d8:	data_out=16'h446;
17'h181d9:	data_out=16'h7b3;
17'h181da:	data_out=16'ha00;
17'h181db:	data_out=16'h8112;
17'h181dc:	data_out=16'h792;
17'h181dd:	data_out=16'ha00;
17'h181de:	data_out=16'ha00;
17'h181df:	data_out=16'h5bb;
17'h181e0:	data_out=16'h529;
17'h181e1:	data_out=16'h277;
17'h181e2:	data_out=16'h9a8;
17'h181e3:	data_out=16'ha00;
17'h181e4:	data_out=16'h4c9;
17'h181e5:	data_out=16'h6ae;
17'h181e6:	data_out=16'h27;
17'h181e7:	data_out=16'h795;
17'h181e8:	data_out=16'h13a;
17'h181e9:	data_out=16'h542;
17'h181ea:	data_out=16'h12c;
17'h181eb:	data_out=16'h4d3;
17'h181ec:	data_out=16'ha00;
17'h181ed:	data_out=16'ha00;
17'h181ee:	data_out=16'h12c;
17'h181ef:	data_out=16'h9f8;
17'h181f0:	data_out=16'h12f;
17'h181f1:	data_out=16'h56c;
17'h181f2:	data_out=16'h7bd;
17'h181f3:	data_out=16'h85a;
17'h181f4:	data_out=16'h448;
17'h181f5:	data_out=16'h2e7;
17'h181f6:	data_out=16'h23f;
17'h181f7:	data_out=16'ha00;
17'h181f8:	data_out=16'h192;
17'h181f9:	data_out=16'ha00;
17'h181fa:	data_out=16'ha00;
17'h181fb:	data_out=16'h147;
17'h181fc:	data_out=16'h190;
17'h181fd:	data_out=16'h8009;
17'h181fe:	data_out=16'h932;
17'h181ff:	data_out=16'h31a;
17'h18200:	data_out=16'ha00;
17'h18201:	data_out=16'ha00;
17'h18202:	data_out=16'h652;
17'h18203:	data_out=16'ha00;
17'h18204:	data_out=16'h9a7;
17'h18205:	data_out=16'h9ec;
17'h18206:	data_out=16'h499;
17'h18207:	data_out=16'h9a2;
17'h18208:	data_out=16'h63c;
17'h18209:	data_out=16'h45e;
17'h1820a:	data_out=16'h6e2;
17'h1820b:	data_out=16'h45b;
17'h1820c:	data_out=16'h6bd;
17'h1820d:	data_out=16'h93c;
17'h1820e:	data_out=16'h158;
17'h1820f:	data_out=16'h954;
17'h18210:	data_out=16'h7a3;
17'h18211:	data_out=16'h8f5;
17'h18212:	data_out=16'ha00;
17'h18213:	data_out=16'ha00;
17'h18214:	data_out=16'h79a;
17'h18215:	data_out=16'h37a;
17'h18216:	data_out=16'h872;
17'h18217:	data_out=16'h9e1;
17'h18218:	data_out=16'hfd;
17'h18219:	data_out=16'h241;
17'h1821a:	data_out=16'h9e9;
17'h1821b:	data_out=16'ha00;
17'h1821c:	data_out=16'ha00;
17'h1821d:	data_out=16'ha00;
17'h1821e:	data_out=16'ha00;
17'h1821f:	data_out=16'h31d;
17'h18220:	data_out=16'ha00;
17'h18221:	data_out=16'h15a;
17'h18222:	data_out=16'h8f8;
17'h18223:	data_out=16'h8165;
17'h18224:	data_out=16'h8169;
17'h18225:	data_out=16'h5bb;
17'h18226:	data_out=16'h48d;
17'h18227:	data_out=16'ha00;
17'h18228:	data_out=16'h165;
17'h18229:	data_out=16'h9c9;
17'h1822a:	data_out=16'ha00;
17'h1822b:	data_out=16'h448;
17'h1822c:	data_out=16'h710;
17'h1822d:	data_out=16'h758;
17'h1822e:	data_out=16'ha00;
17'h1822f:	data_out=16'ha00;
17'h18230:	data_out=16'h9ed;
17'h18231:	data_out=16'h948;
17'h18232:	data_out=16'h9f1;
17'h18233:	data_out=16'h843;
17'h18234:	data_out=16'ha00;
17'h18235:	data_out=16'h861;
17'h18236:	data_out=16'h9a0;
17'h18237:	data_out=16'h63e;
17'h18238:	data_out=16'ha00;
17'h18239:	data_out=16'h8e9;
17'h1823a:	data_out=16'h7dd;
17'h1823b:	data_out=16'h3ee;
17'h1823c:	data_out=16'h827;
17'h1823d:	data_out=16'ha00;
17'h1823e:	data_out=16'h166;
17'h1823f:	data_out=16'h9ec;
17'h18240:	data_out=16'h9f8;
17'h18241:	data_out=16'h566;
17'h18242:	data_out=16'ha00;
17'h18243:	data_out=16'h8e;
17'h18244:	data_out=16'h674;
17'h18245:	data_out=16'h3af;
17'h18246:	data_out=16'h48c;
17'h18247:	data_out=16'ha00;
17'h18248:	data_out=16'ha00;
17'h18249:	data_out=16'h55a;
17'h1824a:	data_out=16'ha00;
17'h1824b:	data_out=16'ha00;
17'h1824c:	data_out=16'ha00;
17'h1824d:	data_out=16'h9f0;
17'h1824e:	data_out=16'ha00;
17'h1824f:	data_out=16'h957;
17'h18250:	data_out=16'h863;
17'h18251:	data_out=16'h2c6;
17'h18252:	data_out=16'h81a3;
17'h18253:	data_out=16'ha00;
17'h18254:	data_out=16'ha00;
17'h18255:	data_out=16'h31b;
17'h18256:	data_out=16'h446;
17'h18257:	data_out=16'h374;
17'h18258:	data_out=16'h302;
17'h18259:	data_out=16'h9f8;
17'h1825a:	data_out=16'h8d8;
17'h1825b:	data_out=16'h627;
17'h1825c:	data_out=16'h9fe;
17'h1825d:	data_out=16'ha00;
17'h1825e:	data_out=16'ha00;
17'h1825f:	data_out=16'h5ed;
17'h18260:	data_out=16'h580;
17'h18261:	data_out=16'h958;
17'h18262:	data_out=16'h72d;
17'h18263:	data_out=16'h867;
17'h18264:	data_out=16'h936;
17'h18265:	data_out=16'h9eb;
17'h18266:	data_out=16'h1aa;
17'h18267:	data_out=16'h6e9;
17'h18268:	data_out=16'h15b;
17'h18269:	data_out=16'h4df;
17'h1826a:	data_out=16'h155;
17'h1826b:	data_out=16'h9f9;
17'h1826c:	data_out=16'ha00;
17'h1826d:	data_out=16'h896;
17'h1826e:	data_out=16'h155;
17'h1826f:	data_out=16'h9f9;
17'h18270:	data_out=16'h157;
17'h18271:	data_out=16'h82c;
17'h18272:	data_out=16'h9f9;
17'h18273:	data_out=16'h9f9;
17'h18274:	data_out=16'h9e6;
17'h18275:	data_out=16'h5ff;
17'h18276:	data_out=16'h2e1;
17'h18277:	data_out=16'h980;
17'h18278:	data_out=16'h285;
17'h18279:	data_out=16'ha00;
17'h1827a:	data_out=16'h834;
17'h1827b:	data_out=16'h167;
17'h1827c:	data_out=16'h20f;
17'h1827d:	data_out=16'h30a;
17'h1827e:	data_out=16'h473;
17'h1827f:	data_out=16'h7e9;
17'h18280:	data_out=16'ha00;
17'h18281:	data_out=16'ha00;
17'h18282:	data_out=16'h4f4;
17'h18283:	data_out=16'ha00;
17'h18284:	data_out=16'h7a7;
17'h18285:	data_out=16'h8d5;
17'h18286:	data_out=16'h5e;
17'h18287:	data_out=16'h7fe;
17'h18288:	data_out=16'h5c1;
17'h18289:	data_out=16'h2d1;
17'h1828a:	data_out=16'h770;
17'h1828b:	data_out=16'h1c9;
17'h1828c:	data_out=16'h683;
17'h1828d:	data_out=16'h6e4;
17'h1828e:	data_out=16'hec;
17'h1828f:	data_out=16'h821;
17'h18290:	data_out=16'h5a6;
17'h18291:	data_out=16'h7be;
17'h18292:	data_out=16'h8a4;
17'h18293:	data_out=16'h9dd;
17'h18294:	data_out=16'h589;
17'h18295:	data_out=16'h2ec;
17'h18296:	data_out=16'h6f8;
17'h18297:	data_out=16'h7dd;
17'h18298:	data_out=16'hee;
17'h18299:	data_out=16'h1e1;
17'h1829a:	data_out=16'h7ff;
17'h1829b:	data_out=16'ha00;
17'h1829c:	data_out=16'h950;
17'h1829d:	data_out=16'ha00;
17'h1829e:	data_out=16'h98c;
17'h1829f:	data_out=16'h16;
17'h182a0:	data_out=16'ha00;
17'h182a1:	data_out=16'heb;
17'h182a2:	data_out=16'h6c8;
17'h182a3:	data_out=16'h80ae;
17'h182a4:	data_out=16'h80a9;
17'h182a5:	data_out=16'h351;
17'h182a6:	data_out=16'h2de;
17'h182a7:	data_out=16'ha00;
17'h182a8:	data_out=16'hed;
17'h182a9:	data_out=16'h7c1;
17'h182aa:	data_out=16'ha00;
17'h182ab:	data_out=16'h390;
17'h182ac:	data_out=16'h5bf;
17'h182ad:	data_out=16'h645;
17'h182ae:	data_out=16'h8c1;
17'h182af:	data_out=16'ha00;
17'h182b0:	data_out=16'h8bf;
17'h182b1:	data_out=16'h9b7;
17'h182b2:	data_out=16'h931;
17'h182b3:	data_out=16'h635;
17'h182b4:	data_out=16'ha00;
17'h182b5:	data_out=16'h721;
17'h182b6:	data_out=16'h9cb;
17'h182b7:	data_out=16'h4dd;
17'h182b8:	data_out=16'ha00;
17'h182b9:	data_out=16'h70a;
17'h182ba:	data_out=16'h803;
17'h182bb:	data_out=16'h420;
17'h182bc:	data_out=16'h6c8;
17'h182bd:	data_out=16'ha00;
17'h182be:	data_out=16'hee;
17'h182bf:	data_out=16'h8c1;
17'h182c0:	data_out=16'h850;
17'h182c1:	data_out=16'h513;
17'h182c2:	data_out=16'h958;
17'h182c3:	data_out=16'h833d;
17'h182c4:	data_out=16'h4e1;
17'h182c5:	data_out=16'h315;
17'h182c6:	data_out=16'h402;
17'h182c7:	data_out=16'h877;
17'h182c8:	data_out=16'ha00;
17'h182c9:	data_out=16'h2c2;
17'h182ca:	data_out=16'ha00;
17'h182cb:	data_out=16'ha00;
17'h182cc:	data_out=16'h94b;
17'h182cd:	data_out=16'h78d;
17'h182ce:	data_out=16'h9b4;
17'h182cf:	data_out=16'h864;
17'h182d0:	data_out=16'h52d;
17'h182d1:	data_out=16'h8067;
17'h182d2:	data_out=16'h80a7;
17'h182d3:	data_out=16'ha00;
17'h182d4:	data_out=16'ha00;
17'h182d5:	data_out=16'h12c;
17'h182d6:	data_out=16'h2a9;
17'h182d7:	data_out=16'h9e;
17'h182d8:	data_out=16'h15e;
17'h182d9:	data_out=16'h7e6;
17'h182da:	data_out=16'h7fa;
17'h182db:	data_out=16'h511;
17'h182dc:	data_out=16'h9fc;
17'h182dd:	data_out=16'ha00;
17'h182de:	data_out=16'ha00;
17'h182df:	data_out=16'h60b;
17'h182e0:	data_out=16'h493;
17'h182e1:	data_out=16'h770;
17'h182e2:	data_out=16'h586;
17'h182e3:	data_out=16'h669;
17'h182e4:	data_out=16'h82b;
17'h182e5:	data_out=16'h96b;
17'h182e6:	data_out=16'h13b;
17'h182e7:	data_out=16'h57f;
17'h182e8:	data_out=16'he9;
17'h182e9:	data_out=16'h43b;
17'h182ea:	data_out=16'he9;
17'h182eb:	data_out=16'h8f0;
17'h182ec:	data_out=16'ha00;
17'h182ed:	data_out=16'h698;
17'h182ee:	data_out=16'he9;
17'h182ef:	data_out=16'h9e7;
17'h182f0:	data_out=16'hea;
17'h182f1:	data_out=16'h84b;
17'h182f2:	data_out=16'h9e7;
17'h182f3:	data_out=16'h9e5;
17'h182f4:	data_out=16'h8b2;
17'h182f5:	data_out=16'h384;
17'h182f6:	data_out=16'h1fe;
17'h182f7:	data_out=16'h532;
17'h182f8:	data_out=16'h80e8;
17'h182f9:	data_out=16'ha00;
17'h182fa:	data_out=16'h643;
17'h182fb:	data_out=16'hee;
17'h182fc:	data_out=16'h233;
17'h182fd:	data_out=16'h805e;
17'h182fe:	data_out=16'h39;
17'h182ff:	data_out=16'h5f2;
17'h18300:	data_out=16'h7a8;
17'h18301:	data_out=16'h9fc;
17'h18302:	data_out=16'h41f;
17'h18303:	data_out=16'h877;
17'h18304:	data_out=16'h28f;
17'h18305:	data_out=16'h45a;
17'h18306:	data_out=16'h81c1;
17'h18307:	data_out=16'h3f1;
17'h18308:	data_out=16'h35a;
17'h18309:	data_out=16'hc2;
17'h1830a:	data_out=16'h541;
17'h1830b:	data_out=16'h18c;
17'h1830c:	data_out=16'h1ee;
17'h1830d:	data_out=16'h4ac;
17'h1830e:	data_out=16'h4a;
17'h1830f:	data_out=16'h68d;
17'h18310:	data_out=16'h413;
17'h18311:	data_out=16'h307;
17'h18312:	data_out=16'h727;
17'h18313:	data_out=16'h655;
17'h18314:	data_out=16'h4b1;
17'h18315:	data_out=16'h152;
17'h18316:	data_out=16'h3dc;
17'h18317:	data_out=16'h6f2;
17'h18318:	data_out=16'h80b6;
17'h18319:	data_out=16'h50;
17'h1831a:	data_out=16'h2df;
17'h1831b:	data_out=16'ha00;
17'h1831c:	data_out=16'h4cf;
17'h1831d:	data_out=16'h9fe;
17'h1831e:	data_out=16'h78f;
17'h1831f:	data_out=16'h8280;
17'h18320:	data_out=16'ha00;
17'h18321:	data_out=16'h5a;
17'h18322:	data_out=16'h67f;
17'h18323:	data_out=16'h830e;
17'h18324:	data_out=16'h830f;
17'h18325:	data_out=16'h2dc;
17'h18326:	data_out=16'h122;
17'h18327:	data_out=16'h9f7;
17'h18328:	data_out=16'h82;
17'h18329:	data_out=16'h6b9;
17'h1832a:	data_out=16'h8c9;
17'h1832b:	data_out=16'h216;
17'h1832c:	data_out=16'h30e;
17'h1832d:	data_out=16'h6ab;
17'h1832e:	data_out=16'h63c;
17'h1832f:	data_out=16'ha00;
17'h18330:	data_out=16'h406;
17'h18331:	data_out=16'h66a;
17'h18332:	data_out=16'h42c;
17'h18333:	data_out=16'h50e;
17'h18334:	data_out=16'h6c7;
17'h18335:	data_out=16'h257;
17'h18336:	data_out=16'h712;
17'h18337:	data_out=16'h412;
17'h18338:	data_out=16'h674;
17'h18339:	data_out=16'h5b4;
17'h1833a:	data_out=16'h620;
17'h1833b:	data_out=16'h1a;
17'h1833c:	data_out=16'h686;
17'h1833d:	data_out=16'h5e7;
17'h1833e:	data_out=16'h82;
17'h1833f:	data_out=16'h2da;
17'h18340:	data_out=16'h46f;
17'h18341:	data_out=16'h3f9;
17'h18342:	data_out=16'h754;
17'h18343:	data_out=16'h82db;
17'h18344:	data_out=16'h14f;
17'h18345:	data_out=16'h10;
17'h18346:	data_out=16'h499;
17'h18347:	data_out=16'h536;
17'h18348:	data_out=16'h824;
17'h18349:	data_out=16'h263;
17'h1834a:	data_out=16'h71e;
17'h1834b:	data_out=16'h7ce;
17'h1834c:	data_out=16'h5e7;
17'h1834d:	data_out=16'h6f3;
17'h1834e:	data_out=16'h690;
17'h1834f:	data_out=16'h473;
17'h18350:	data_out=16'h228;
17'h18351:	data_out=16'h81b5;
17'h18352:	data_out=16'h8338;
17'h18353:	data_out=16'ha00;
17'h18354:	data_out=16'ha00;
17'h18355:	data_out=16'h1ba;
17'h18356:	data_out=16'h224;
17'h18357:	data_out=16'h8d;
17'h18358:	data_out=16'h238;
17'h18359:	data_out=16'h4e5;
17'h1835a:	data_out=16'h807;
17'h1835b:	data_out=16'h811b;
17'h1835c:	data_out=16'h790;
17'h1835d:	data_out=16'ha00;
17'h1835e:	data_out=16'ha00;
17'h1835f:	data_out=16'h4af;
17'h18360:	data_out=16'h2eb;
17'h18361:	data_out=16'h256;
17'h18362:	data_out=16'h3f5;
17'h18363:	data_out=16'h53e;
17'h18364:	data_out=16'h4c8;
17'h18365:	data_out=16'h619;
17'h18366:	data_out=16'h6d;
17'h18367:	data_out=16'h408;
17'h18368:	data_out=16'h5e;
17'h18369:	data_out=16'h392;
17'h1836a:	data_out=16'h2d;
17'h1836b:	data_out=16'h3b5;
17'h1836c:	data_out=16'ha00;
17'h1836d:	data_out=16'h562;
17'h1836e:	data_out=16'h3c;
17'h1836f:	data_out=16'h83c;
17'h18370:	data_out=16'h4c;
17'h18371:	data_out=16'h458;
17'h18372:	data_out=16'h41c;
17'h18373:	data_out=16'h57a;
17'h18374:	data_out=16'h3fb;
17'h18375:	data_out=16'h21a;
17'h18376:	data_out=16'hde;
17'h18377:	data_out=16'h23b;
17'h18378:	data_out=16'h81da;
17'h18379:	data_out=16'h754;
17'h1837a:	data_out=16'h52d;
17'h1837b:	data_out=16'h85;
17'h1837c:	data_out=16'h62;
17'h1837d:	data_out=16'h82eb;
17'h1837e:	data_out=16'h80a7;
17'h1837f:	data_out=16'h137;
17'h18380:	data_out=16'h4c9;
17'h18381:	data_out=16'h751;
17'h18382:	data_out=16'h344;
17'h18383:	data_out=16'h641;
17'h18384:	data_out=16'h275;
17'h18385:	data_out=16'h3d2;
17'h18386:	data_out=16'h8025;
17'h18387:	data_out=16'h2d2;
17'h18388:	data_out=16'h27b;
17'h18389:	data_out=16'h55;
17'h1838a:	data_out=16'h3f3;
17'h1838b:	data_out=16'h12d;
17'h1838c:	data_out=16'h1da;
17'h1838d:	data_out=16'h368;
17'h1838e:	data_out=16'h34;
17'h1838f:	data_out=16'h4ae;
17'h18390:	data_out=16'h255;
17'h18391:	data_out=16'h291;
17'h18392:	data_out=16'h4f4;
17'h18393:	data_out=16'h46f;
17'h18394:	data_out=16'h376;
17'h18395:	data_out=16'h161;
17'h18396:	data_out=16'h2ec;
17'h18397:	data_out=16'h4c8;
17'h18398:	data_out=16'h80a0;
17'h18399:	data_out=16'h106;
17'h1839a:	data_out=16'h244;
17'h1839b:	data_out=16'h76b;
17'h1839c:	data_out=16'h454;
17'h1839d:	data_out=16'h75b;
17'h1839e:	data_out=16'h515;
17'h1839f:	data_out=16'h80cd;
17'h183a0:	data_out=16'h8eb;
17'h183a1:	data_out=16'h35;
17'h183a2:	data_out=16'h41b;
17'h183a3:	data_out=16'h81e9;
17'h183a4:	data_out=16'h81d6;
17'h183a5:	data_out=16'h25d;
17'h183a6:	data_out=16'h49;
17'h183a7:	data_out=16'h7b7;
17'h183a8:	data_out=16'h41;
17'h183a9:	data_out=16'h45c;
17'h183aa:	data_out=16'h4f0;
17'h183ab:	data_out=16'h244;
17'h183ac:	data_out=16'h270;
17'h183ad:	data_out=16'h3f8;
17'h183ae:	data_out=16'h480;
17'h183af:	data_out=16'h9d6;
17'h183b0:	data_out=16'h334;
17'h183b1:	data_out=16'h476;
17'h183b2:	data_out=16'h367;
17'h183b3:	data_out=16'h3a8;
17'h183b4:	data_out=16'h3d8;
17'h183b5:	data_out=16'h23c;
17'h183b6:	data_out=16'h461;
17'h183b7:	data_out=16'h33d;
17'h183b8:	data_out=16'h3df;
17'h183b9:	data_out=16'h406;
17'h183ba:	data_out=16'h3ff;
17'h183bb:	data_out=16'h72;
17'h183bc:	data_out=16'h533;
17'h183bd:	data_out=16'h427;
17'h183be:	data_out=16'h4f;
17'h183bf:	data_out=16'h293;
17'h183c0:	data_out=16'h2b4;
17'h183c1:	data_out=16'h329;
17'h183c2:	data_out=16'h4b0;
17'h183c3:	data_out=16'h80ed;
17'h183c4:	data_out=16'h178;
17'h183c5:	data_out=16'h29;
17'h183c6:	data_out=16'h347;
17'h183c7:	data_out=16'h325;
17'h183c8:	data_out=16'h553;
17'h183c9:	data_out=16'h224;
17'h183ca:	data_out=16'h422;
17'h183cb:	data_out=16'h58b;
17'h183cc:	data_out=16'h3f2;
17'h183cd:	data_out=16'h46b;
17'h183ce:	data_out=16'h484;
17'h183cf:	data_out=16'h287;
17'h183d0:	data_out=16'h1b9;
17'h183d1:	data_out=16'h70;
17'h183d2:	data_out=16'h81ab;
17'h183d3:	data_out=16'ha00;
17'h183d4:	data_out=16'h971;
17'h183d5:	data_out=16'h1be;
17'h183d6:	data_out=16'h1f3;
17'h183d7:	data_out=16'h101;
17'h183d8:	data_out=16'h234;
17'h183d9:	data_out=16'h35e;
17'h183da:	data_out=16'h601;
17'h183db:	data_out=16'h7b;
17'h183dc:	data_out=16'h602;
17'h183dd:	data_out=16'h725;
17'h183de:	data_out=16'h9bc;
17'h183df:	data_out=16'h33b;
17'h183e0:	data_out=16'h18d;
17'h183e1:	data_out=16'h21c;
17'h183e2:	data_out=16'h30f;
17'h183e3:	data_out=16'h3c0;
17'h183e4:	data_out=16'h330;
17'h183e5:	data_out=16'h47f;
17'h183e6:	data_out=16'hce;
17'h183e7:	data_out=16'h2f1;
17'h183e8:	data_out=16'h3a;
17'h183e9:	data_out=16'h2a8;
17'h183ea:	data_out=16'h17;
17'h183eb:	data_out=16'h347;
17'h183ec:	data_out=16'ha00;
17'h183ed:	data_out=16'h3d4;
17'h183ee:	data_out=16'h20;
17'h183ef:	data_out=16'h5f1;
17'h183f0:	data_out=16'h27;
17'h183f1:	data_out=16'h249;
17'h183f2:	data_out=16'h35e;
17'h183f3:	data_out=16'h40f;
17'h183f4:	data_out=16'h32b;
17'h183f5:	data_out=16'h1f7;
17'h183f6:	data_out=16'h11a;
17'h183f7:	data_out=16'h10c;
17'h183f8:	data_out=16'h806d;
17'h183f9:	data_out=16'h487;
17'h183fa:	data_out=16'h3b7;
17'h183fb:	data_out=16'h4c;
17'h183fc:	data_out=16'h7c;
17'h183fd:	data_out=16'h81c5;
17'h183fe:	data_out=16'h8027;
17'h183ff:	data_out=16'h14a;
17'h18400:	data_out=16'h10f;
17'h18401:	data_out=16'h224;
17'h18402:	data_out=16'h284;
17'h18403:	data_out=16'h2f3;
17'h18404:	data_out=16'h816b;
17'h18405:	data_out=16'h74;
17'h18406:	data_out=16'h8167;
17'h18407:	data_out=16'h66;
17'h18408:	data_out=16'had;
17'h18409:	data_out=16'ha;
17'h1840a:	data_out=16'h801f;
17'h1840b:	data_out=16'hb1;
17'h1840c:	data_out=16'h80dd;
17'h1840d:	data_out=16'hdc;
17'h1840e:	data_out=16'h8025;
17'h1840f:	data_out=16'h236;
17'h18410:	data_out=16'h1b2;
17'h18411:	data_out=16'h81d3;
17'h18412:	data_out=16'h43e;
17'h18413:	data_out=16'h175;
17'h18414:	data_out=16'h32d;
17'h18415:	data_out=16'h80d0;
17'h18416:	data_out=16'h2d;
17'h18417:	data_out=16'h3ff;
17'h18418:	data_out=16'h8055;
17'h18419:	data_out=16'h818d;
17'h1841a:	data_out=16'h820b;
17'h1841b:	data_out=16'h4cd;
17'h1841c:	data_out=16'he1;
17'h1841d:	data_out=16'h2db;
17'h1841e:	data_out=16'h3db;
17'h1841f:	data_out=16'h80c5;
17'h18420:	data_out=16'h4a9;
17'h18421:	data_out=16'h8022;
17'h18422:	data_out=16'h256;
17'h18423:	data_out=16'h81fc;
17'h18424:	data_out=16'h81fd;
17'h18425:	data_out=16'hd8;
17'h18426:	data_out=16'hb0;
17'h18427:	data_out=16'h34d;
17'h18428:	data_out=16'h8015;
17'h18429:	data_out=16'h1ca;
17'h1842a:	data_out=16'h323;
17'h1842b:	data_out=16'h804a;
17'h1842c:	data_out=16'h2d;
17'h1842d:	data_out=16'h157;
17'h1842e:	data_out=16'h414;
17'h1842f:	data_out=16'h529;
17'h18430:	data_out=16'h81ba;
17'h18431:	data_out=16'h813a;
17'h18432:	data_out=16'h81b0;
17'h18433:	data_out=16'h325;
17'h18434:	data_out=16'h8097;
17'h18435:	data_out=16'h8242;
17'h18436:	data_out=16'h260;
17'h18437:	data_out=16'h283;
17'h18438:	data_out=16'h80c5;
17'h18439:	data_out=16'h2bf;
17'h1843a:	data_out=16'h287;
17'h1843b:	data_out=16'h8267;
17'h1843c:	data_out=16'h3d2;
17'h1843d:	data_out=16'hba;
17'h1843e:	data_out=16'h8017;
17'h1843f:	data_out=16'h80ef;
17'h18440:	data_out=16'hd7;
17'h18441:	data_out=16'h321;
17'h18442:	data_out=16'h12a;
17'h18443:	data_out=16'h810c;
17'h18444:	data_out=16'h80ee;
17'h18445:	data_out=16'h811d;
17'h18446:	data_out=16'h267;
17'h18447:	data_out=16'h126;
17'h18448:	data_out=16'h40e;
17'h18449:	data_out=16'he1;
17'h1844a:	data_out=16'h2f;
17'h1844b:	data_out=16'hb7;
17'h1844c:	data_out=16'hf0;
17'h1844d:	data_out=16'h26c;
17'h1844e:	data_out=16'h28c;
17'h1844f:	data_out=16'h8014;
17'h18450:	data_out=16'h148;
17'h18451:	data_out=16'h81da;
17'h18452:	data_out=16'h8215;
17'h18453:	data_out=16'h541;
17'h18454:	data_out=16'h42d;
17'h18455:	data_out=16'h1f0;
17'h18456:	data_out=16'h22e;
17'h18457:	data_out=16'h15f;
17'h18458:	data_out=16'h227;
17'h18459:	data_out=16'h133;
17'h1845a:	data_out=16'h4b9;
17'h1845b:	data_out=16'h82d4;
17'h1845c:	data_out=16'h173;
17'h1845d:	data_out=16'h3d5;
17'h1845e:	data_out=16'h499;
17'h1845f:	data_out=16'h1af;
17'h18460:	data_out=16'h8005;
17'h18461:	data_out=16'h8246;
17'h18462:	data_out=16'h2bb;
17'h18463:	data_out=16'h335;
17'h18464:	data_out=16'h8072;
17'h18465:	data_out=16'h4e;
17'h18466:	data_out=16'h80f8;
17'h18467:	data_out=16'h24f;
17'h18468:	data_out=16'h8019;
17'h18469:	data_out=16'h17e;
17'h1846a:	data_out=16'h802d;
17'h1846b:	data_out=16'h8159;
17'h1846c:	data_out=16'h531;
17'h1846d:	data_out=16'h33d;
17'h1846e:	data_out=16'h8033;
17'h1846f:	data_out=16'h190;
17'h18470:	data_out=16'h8020;
17'h18471:	data_out=16'h1a1;
17'h18472:	data_out=16'h8004;
17'h18473:	data_out=16'h8085;
17'h18474:	data_out=16'h81c6;
17'h18475:	data_out=16'h8106;
17'h18476:	data_out=16'h808f;
17'h18477:	data_out=16'h8001;
17'h18478:	data_out=16'h81d3;
17'h18479:	data_out=16'h40a;
17'h1847a:	data_out=16'h34a;
17'h1847b:	data_out=16'h8010;
17'h1847c:	data_out=16'h77;
17'h1847d:	data_out=16'h821c;
17'h1847e:	data_out=16'h8012;
17'h1847f:	data_out=16'h80c5;
17'h18480:	data_out=16'h12b;
17'h18481:	data_out=16'h19c;
17'h18482:	data_out=16'h1da;
17'h18483:	data_out=16'h78;
17'h18484:	data_out=16'h84e1;
17'h18485:	data_out=16'h833f;
17'h18486:	data_out=16'h83bc;
17'h18487:	data_out=16'h81e9;
17'h18488:	data_out=16'h92;
17'h18489:	data_out=16'h8097;
17'h1848a:	data_out=16'h81d2;
17'h1848b:	data_out=16'h94;
17'h1848c:	data_out=16'h8379;
17'h1848d:	data_out=16'ha4;
17'h1848e:	data_out=16'h80a8;
17'h1848f:	data_out=16'h90;
17'h18490:	data_out=16'h189;
17'h18491:	data_out=16'h85ba;
17'h18492:	data_out=16'h38c;
17'h18493:	data_out=16'h8041;
17'h18494:	data_out=16'h2da;
17'h18495:	data_out=16'h81d8;
17'h18496:	data_out=16'h81fc;
17'h18497:	data_out=16'h3b5;
17'h18498:	data_out=16'h80c3;
17'h18499:	data_out=16'h820c;
17'h1849a:	data_out=16'h853f;
17'h1849b:	data_out=16'h526;
17'h1849c:	data_out=16'h8278;
17'h1849d:	data_out=16'h181;
17'h1849e:	data_out=16'h397;
17'h1849f:	data_out=16'h835c;
17'h184a0:	data_out=16'h43d;
17'h184a1:	data_out=16'h80a6;
17'h184a2:	data_out=16'h26b;
17'h184a3:	data_out=16'h81fd;
17'h184a4:	data_out=16'h81fe;
17'h184a5:	data_out=16'h91;
17'h184a6:	data_out=16'h809e;
17'h184a7:	data_out=16'h212;
17'h184a8:	data_out=16'h80a9;
17'h184a9:	data_out=16'h1ec;
17'h184aa:	data_out=16'h25f;
17'h184ab:	data_out=16'h808d;
17'h184ac:	data_out=16'h81e4;
17'h184ad:	data_out=16'h19f;
17'h184ae:	data_out=16'h39d;
17'h184af:	data_out=16'h469;
17'h184b0:	data_out=16'h8572;
17'h184b1:	data_out=16'h82e9;
17'h184b2:	data_out=16'h8570;
17'h184b3:	data_out=16'h2da;
17'h184b4:	data_out=16'h8269;
17'h184b5:	data_out=16'h855c;
17'h184b6:	data_out=16'h262;
17'h184b7:	data_out=16'h1d0;
17'h184b8:	data_out=16'h8385;
17'h184b9:	data_out=16'h1ff;
17'h184ba:	data_out=16'h20a;
17'h184bb:	data_out=16'h84ab;
17'h184bc:	data_out=16'h3ba;
17'h184bd:	data_out=16'h8205;
17'h184be:	data_out=16'h80b1;
17'h184bf:	data_out=16'h8414;
17'h184c0:	data_out=16'h81ed;
17'h184c1:	data_out=16'h2d3;
17'h184c2:	data_out=16'h24;
17'h184c3:	data_out=16'h8394;
17'h184c4:	data_out=16'h83b6;
17'h184c5:	data_out=16'h81e0;
17'h184c6:	data_out=16'h2aa;
17'h184c7:	data_out=16'h8012;
17'h184c8:	data_out=16'h326;
17'h184c9:	data_out=16'h76;
17'h184ca:	data_out=16'h812f;
17'h184cb:	data_out=16'h8080;
17'h184cc:	data_out=16'h8082;
17'h184cd:	data_out=16'h2a2;
17'h184ce:	data_out=16'h228;
17'h184cf:	data_out=16'h80ca;
17'h184d0:	data_out=16'h8125;
17'h184d1:	data_out=16'h8447;
17'h184d2:	data_out=16'h81e7;
17'h184d3:	data_out=16'h51a;
17'h184d4:	data_out=16'h3de;
17'h184d5:	data_out=16'h55;
17'h184d6:	data_out=16'h13d;
17'h184d7:	data_out=16'h120;
17'h184d8:	data_out=16'h120;
17'h184d9:	data_out=16'h8110;
17'h184da:	data_out=16'h613;
17'h184db:	data_out=16'h85a9;
17'h184dc:	data_out=16'h8063;
17'h184dd:	data_out=16'h32d;
17'h184de:	data_out=16'h431;
17'h184df:	data_out=16'h169;
17'h184e0:	data_out=16'h8103;
17'h184e1:	data_out=16'h8552;
17'h184e2:	data_out=16'h2b7;
17'h184e3:	data_out=16'h2ef;
17'h184e4:	data_out=16'h8337;
17'h184e5:	data_out=16'h82c4;
17'h184e6:	data_out=16'h821d;
17'h184e7:	data_out=16'h20e;
17'h184e8:	data_out=16'h80af;
17'h184e9:	data_out=16'hfe;
17'h184ea:	data_out=16'h80b2;
17'h184eb:	data_out=16'h8504;
17'h184ec:	data_out=16'h604;
17'h184ed:	data_out=16'h2f5;
17'h184ee:	data_out=16'h80ae;
17'h184ef:	data_out=16'h8153;
17'h184f0:	data_out=16'h80ac;
17'h184f1:	data_out=16'h22;
17'h184f2:	data_out=16'h83cb;
17'h184f3:	data_out=16'h8472;
17'h184f4:	data_out=16'h8574;
17'h184f5:	data_out=16'h83fd;
17'h184f6:	data_out=16'h81a5;
17'h184f7:	data_out=16'h8214;
17'h184f8:	data_out=16'h8462;
17'h184f9:	data_out=16'h304;
17'h184fa:	data_out=16'h301;
17'h184fb:	data_out=16'h80a1;
17'h184fc:	data_out=16'h8015;
17'h184fd:	data_out=16'h8477;
17'h184fe:	data_out=16'h80cf;
17'h184ff:	data_out=16'h82c1;
17'h18500:	data_out=16'h96;
17'h18501:	data_out=16'hba;
17'h18502:	data_out=16'h239;
17'h18503:	data_out=16'h32;
17'h18504:	data_out=16'h8777;
17'h18505:	data_out=16'h850a;
17'h18506:	data_out=16'h8403;
17'h18507:	data_out=16'h8472;
17'h18508:	data_out=16'h130;
17'h18509:	data_out=16'h809d;
17'h1850a:	data_out=16'h83f8;
17'h1850b:	data_out=16'hf3;
17'h1850c:	data_out=16'h85e0;
17'h1850d:	data_out=16'hed;
17'h1850e:	data_out=16'h80cf;
17'h1850f:	data_out=16'h116;
17'h18510:	data_out=16'h1c8;
17'h18511:	data_out=16'h884c;
17'h18512:	data_out=16'h349;
17'h18513:	data_out=16'h8035;
17'h18514:	data_out=16'h387;
17'h18515:	data_out=16'h8232;
17'h18516:	data_out=16'h82ad;
17'h18517:	data_out=16'h495;
17'h18518:	data_out=16'h80b5;
17'h18519:	data_out=16'h8278;
17'h1851a:	data_out=16'h870f;
17'h1851b:	data_out=16'h63f;
17'h1851c:	data_out=16'h83c0;
17'h1851d:	data_out=16'h8049;
17'h1851e:	data_out=16'h3dc;
17'h1851f:	data_out=16'h8422;
17'h18520:	data_out=16'h371;
17'h18521:	data_out=16'h80ca;
17'h18522:	data_out=16'h246;
17'h18523:	data_out=16'h8241;
17'h18524:	data_out=16'h8241;
17'h18525:	data_out=16'h8089;
17'h18526:	data_out=16'h8059;
17'h18527:	data_out=16'h8d;
17'h18528:	data_out=16'h80cb;
17'h18529:	data_out=16'h343;
17'h1852a:	data_out=16'h231;
17'h1852b:	data_out=16'h80f0;
17'h1852c:	data_out=16'h82ec;
17'h1852d:	data_out=16'h1f2;
17'h1852e:	data_out=16'h4a2;
17'h1852f:	data_out=16'h4d5;
17'h18530:	data_out=16'h8777;
17'h18531:	data_out=16'h85a7;
17'h18532:	data_out=16'h8769;
17'h18533:	data_out=16'h36f;
17'h18534:	data_out=16'h83ea;
17'h18535:	data_out=16'h876a;
17'h18536:	data_out=16'h387;
17'h18537:	data_out=16'h21f;
17'h18538:	data_out=16'h8457;
17'h18539:	data_out=16'h29d;
17'h1853a:	data_out=16'h151;
17'h1853b:	data_out=16'h86dc;
17'h1853c:	data_out=16'h455;
17'h1853d:	data_out=16'h8308;
17'h1853e:	data_out=16'h80c0;
17'h1853f:	data_out=16'h85a1;
17'h18540:	data_out=16'h8308;
17'h18541:	data_out=16'h387;
17'h18542:	data_out=16'h805d;
17'h18543:	data_out=16'h83c5;
17'h18544:	data_out=16'h8604;
17'h18545:	data_out=16'h823f;
17'h18546:	data_out=16'h30e;
17'h18547:	data_out=16'h8065;
17'h18548:	data_out=16'h342;
17'h18549:	data_out=16'h8095;
17'h1854a:	data_out=16'h830e;
17'h1854b:	data_out=16'h81d7;
17'h1854c:	data_out=16'h8120;
17'h1854d:	data_out=16'h277;
17'h1854e:	data_out=16'h243;
17'h1854f:	data_out=16'h81b9;
17'h18550:	data_out=16'h81b4;
17'h18551:	data_out=16'h84b4;
17'h18552:	data_out=16'h8255;
17'h18553:	data_out=16'h4c4;
17'h18554:	data_out=16'h473;
17'h18555:	data_out=16'hc2;
17'h18556:	data_out=16'haa;
17'h18557:	data_out=16'hb9;
17'h18558:	data_out=16'h1ac;
17'h18559:	data_out=16'h8246;
17'h1855a:	data_out=16'h769;
17'h1855b:	data_out=16'h874f;
17'h1855c:	data_out=16'h820d;
17'h1855d:	data_out=16'h261;
17'h1855e:	data_out=16'h4e7;
17'h1855f:	data_out=16'h124;
17'h18560:	data_out=16'h814f;
17'h18561:	data_out=16'h873b;
17'h18562:	data_out=16'h30b;
17'h18563:	data_out=16'h38f;
17'h18564:	data_out=16'h84ad;
17'h18565:	data_out=16'h84e8;
17'h18566:	data_out=16'h82d1;
17'h18567:	data_out=16'h23d;
17'h18568:	data_out=16'h80c9;
17'h18569:	data_out=16'h10d;
17'h1856a:	data_out=16'h80cf;
17'h1856b:	data_out=16'h86d1;
17'h1856c:	data_out=16'h4c0;
17'h1856d:	data_out=16'h390;
17'h1856e:	data_out=16'h80d0;
17'h1856f:	data_out=16'h82ef;
17'h18570:	data_out=16'h80ca;
17'h18571:	data_out=16'h8061;
17'h18572:	data_out=16'h85c1;
17'h18573:	data_out=16'h8629;
17'h18574:	data_out=16'h877a;
17'h18575:	data_out=16'h8478;
17'h18576:	data_out=16'h81e9;
17'h18577:	data_out=16'h8240;
17'h18578:	data_out=16'h84b1;
17'h18579:	data_out=16'h37a;
17'h1857a:	data_out=16'h3ad;
17'h1857b:	data_out=16'h80cb;
17'h1857c:	data_out=16'h8088;
17'h1857d:	data_out=16'h8504;
17'h1857e:	data_out=16'h803b;
17'h1857f:	data_out=16'h846a;
17'h18580:	data_out=16'hc;
17'h18581:	data_out=16'h2c;
17'h18582:	data_out=16'h8e;
17'h18583:	data_out=16'h47;
17'h18584:	data_out=16'h80d0;
17'h18585:	data_out=16'h8067;
17'h18586:	data_out=16'h80c0;
17'h18587:	data_out=16'h8083;
17'h18588:	data_out=16'h11;
17'h18589:	data_out=16'h803e;
17'h1858a:	data_out=16'h806e;
17'h1858b:	data_out=16'h804a;
17'h1858c:	data_out=16'h80a5;
17'h1858d:	data_out=16'hd;
17'h1858e:	data_out=16'h801c;
17'h1858f:	data_out=16'h2c;
17'h18590:	data_out=16'h3b;
17'h18591:	data_out=16'h811d;
17'h18592:	data_out=16'hbf;
17'h18593:	data_out=16'h8027;
17'h18594:	data_out=16'h116;
17'h18595:	data_out=16'h806f;
17'h18596:	data_out=16'h8076;
17'h18597:	data_out=16'h143;
17'h18598:	data_out=16'h803a;
17'h18599:	data_out=16'h80b3;
17'h1859a:	data_out=16'h80f9;
17'h1859b:	data_out=16'hd0;
17'h1859c:	data_out=16'h32;
17'h1859d:	data_out=16'h8e;
17'h1859e:	data_out=16'h11a;
17'h1859f:	data_out=16'h8082;
17'h185a0:	data_out=16'h105;
17'h185a1:	data_out=16'h801b;
17'h185a2:	data_out=16'h91;
17'h185a3:	data_out=16'h80a5;
17'h185a4:	data_out=16'h80af;
17'h185a5:	data_out=16'h8014;
17'h185a6:	data_out=16'h803b;
17'h185a7:	data_out=16'h9c;
17'h185a8:	data_out=16'h8017;
17'h185a9:	data_out=16'h83;
17'h185aa:	data_out=16'h64;
17'h185ab:	data_out=16'h804b;
17'h185ac:	data_out=16'h8050;
17'h185ad:	data_out=16'h8007;
17'h185ae:	data_out=16'hd9;
17'h185af:	data_out=16'hbf;
17'h185b0:	data_out=16'h812e;
17'h185b1:	data_out=16'h80ca;
17'h185b2:	data_out=16'h811a;
17'h185b3:	data_out=16'h11d;
17'h185b4:	data_out=16'h80ab;
17'h185b5:	data_out=16'h8119;
17'h185b6:	data_out=16'h84;
17'h185b7:	data_out=16'hb3;
17'h185b8:	data_out=16'h809c;
17'h185b9:	data_out=16'h7a;
17'h185ba:	data_out=16'h7c;
17'h185bb:	data_out=16'h811a;
17'h185bc:	data_out=16'hc0;
17'h185bd:	data_out=16'h802f;
17'h185be:	data_out=16'h801f;
17'h185bf:	data_out=16'h80c9;
17'h185c0:	data_out=16'h802f;
17'h185c1:	data_out=16'hfa;
17'h185c2:	data_out=16'h8048;
17'h185c3:	data_out=16'h8092;
17'h185c4:	data_out=16'h80e7;
17'h185c5:	data_out=16'h808d;
17'h185c6:	data_out=16'hc3;
17'h185c7:	data_out=16'h20;
17'h185c8:	data_out=16'h89;
17'h185c9:	data_out=16'h802b;
17'h185ca:	data_out=16'h807d;
17'h185cb:	data_out=16'h8040;
17'h185cc:	data_out=16'h803e;
17'h185cd:	data_out=16'h91;
17'h185ce:	data_out=16'h59;
17'h185cf:	data_out=16'h8065;
17'h185d0:	data_out=16'h8008;
17'h185d1:	data_out=16'h80db;
17'h185d2:	data_out=16'h80a7;
17'h185d3:	data_out=16'h197;
17'h185d4:	data_out=16'ha7;
17'h185d5:	data_out=16'h801c;
17'h185d6:	data_out=16'h70;
17'h185d7:	data_out=16'h36;
17'h185d8:	data_out=16'h2c;
17'h185d9:	data_out=16'h800d;
17'h185da:	data_out=16'h12e;
17'h185db:	data_out=16'h810f;
17'h185dc:	data_out=16'h801d;
17'h185dd:	data_out=16'h85;
17'h185de:	data_out=16'ha6;
17'h185df:	data_out=16'h4b;
17'h185e0:	data_out=16'h8073;
17'h185e1:	data_out=16'h8106;
17'h185e2:	data_out=16'h74;
17'h185e3:	data_out=16'h122;
17'h185e4:	data_out=16'h80ce;
17'h185e5:	data_out=16'h80d4;
17'h185e6:	data_out=16'h80ac;
17'h185e7:	data_out=16'h59;
17'h185e8:	data_out=16'h8021;
17'h185e9:	data_out=16'h26;
17'h185ea:	data_out=16'h8013;
17'h185eb:	data_out=16'h80e6;
17'h185ec:	data_out=16'h104;
17'h185ed:	data_out=16'h123;
17'h185ee:	data_out=16'h8011;
17'h185ef:	data_out=16'h800a;
17'h185f0:	data_out=16'h8013;
17'h185f1:	data_out=16'h17;
17'h185f2:	data_out=16'h80af;
17'h185f3:	data_out=16'h80db;
17'h185f4:	data_out=16'h812f;
17'h185f5:	data_out=16'h80bb;
17'h185f6:	data_out=16'h8071;
17'h185f7:	data_out=16'h809a;
17'h185f8:	data_out=16'h80f7;
17'h185f9:	data_out=16'hba;
17'h185fa:	data_out=16'h126;
17'h185fb:	data_out=16'h8018;
17'h185fc:	data_out=16'h801c;
17'h185fd:	data_out=16'h80fe;
17'h185fe:	data_out=16'h804d;
17'h185ff:	data_out=16'h8094;
17'h18600:	data_out=16'h8004;
17'h18601:	data_out=16'h8001;
17'h18602:	data_out=16'h1;
17'h18603:	data_out=16'h8002;
17'h18604:	data_out=16'h8006;
17'h18605:	data_out=16'h7;
17'h18606:	data_out=16'h2;
17'h18607:	data_out=16'h8006;
17'h18608:	data_out=16'h7;
17'h18609:	data_out=16'h8002;
17'h1860a:	data_out=16'h2;
17'h1860b:	data_out=16'h8003;
17'h1860c:	data_out=16'h5;
17'h1860d:	data_out=16'h8001;
17'h1860e:	data_out=16'h0;
17'h1860f:	data_out=16'h1;
17'h18610:	data_out=16'h9;
17'h18611:	data_out=16'h1;
17'h18612:	data_out=16'h3;
17'h18613:	data_out=16'h8008;
17'h18614:	data_out=16'h8005;
17'h18615:	data_out=16'h8006;
17'h18616:	data_out=16'h8004;
17'h18617:	data_out=16'h8003;
17'h18618:	data_out=16'h2;
17'h18619:	data_out=16'h9;
17'h1861a:	data_out=16'h5;
17'h1861b:	data_out=16'h8007;
17'h1861c:	data_out=16'h6;
17'h1861d:	data_out=16'h8009;
17'h1861e:	data_out=16'h8008;
17'h1861f:	data_out=16'h8007;
17'h18620:	data_out=16'h8001;
17'h18621:	data_out=16'h2;
17'h18622:	data_out=16'h8000;
17'h18623:	data_out=16'h2;
17'h18624:	data_out=16'h0;
17'h18625:	data_out=16'h8007;
17'h18626:	data_out=16'h5;
17'h18627:	data_out=16'h8002;
17'h18628:	data_out=16'h0;
17'h18629:	data_out=16'h8002;
17'h1862a:	data_out=16'h5;
17'h1862b:	data_out=16'h8004;
17'h1862c:	data_out=16'h6;
17'h1862d:	data_out=16'h8004;
17'h1862e:	data_out=16'h6;
17'h1862f:	data_out=16'h6;
17'h18630:	data_out=16'h6;
17'h18631:	data_out=16'h8000;
17'h18632:	data_out=16'h7;
17'h18633:	data_out=16'h8008;
17'h18634:	data_out=16'h3;
17'h18635:	data_out=16'h8006;
17'h18636:	data_out=16'h8003;
17'h18637:	data_out=16'h8005;
17'h18638:	data_out=16'h8006;
17'h18639:	data_out=16'h8006;
17'h1863a:	data_out=16'h8003;
17'h1863b:	data_out=16'h9;
17'h1863c:	data_out=16'h8006;
17'h1863d:	data_out=16'h8002;
17'h1863e:	data_out=16'h8008;
17'h1863f:	data_out=16'h2;
17'h18640:	data_out=16'h8009;
17'h18641:	data_out=16'h1;
17'h18642:	data_out=16'h8006;
17'h18643:	data_out=16'h0;
17'h18644:	data_out=16'h4;
17'h18645:	data_out=16'h9;
17'h18646:	data_out=16'h8;
17'h18647:	data_out=16'h8005;
17'h18648:	data_out=16'h8003;
17'h18649:	data_out=16'h4;
17'h1864a:	data_out=16'h8000;
17'h1864b:	data_out=16'h8005;
17'h1864c:	data_out=16'h9;
17'h1864d:	data_out=16'h8004;
17'h1864e:	data_out=16'h8009;
17'h1864f:	data_out=16'h6;
17'h18650:	data_out=16'h5;
17'h18651:	data_out=16'h8;
17'h18652:	data_out=16'h6;
17'h18653:	data_out=16'h8002;
17'h18654:	data_out=16'h8007;
17'h18655:	data_out=16'h8005;
17'h18656:	data_out=16'h3;
17'h18657:	data_out=16'h8004;
17'h18658:	data_out=16'h8003;
17'h18659:	data_out=16'h8009;
17'h1865a:	data_out=16'h8004;
17'h1865b:	data_out=16'h8000;
17'h1865c:	data_out=16'h8001;
17'h1865d:	data_out=16'h8003;
17'h1865e:	data_out=16'h8008;
17'h1865f:	data_out=16'h8001;
17'h18660:	data_out=16'h8;
17'h18661:	data_out=16'h8004;
17'h18662:	data_out=16'h9;
17'h18663:	data_out=16'h2;
17'h18664:	data_out=16'h8005;
17'h18665:	data_out=16'h7;
17'h18666:	data_out=16'h6;
17'h18667:	data_out=16'h2;
17'h18668:	data_out=16'h2;
17'h18669:	data_out=16'h8004;
17'h1866a:	data_out=16'h6;
17'h1866b:	data_out=16'h1;
17'h1866c:	data_out=16'h2;
17'h1866d:	data_out=16'h6;
17'h1866e:	data_out=16'h8002;
17'h1866f:	data_out=16'h8002;
17'h18670:	data_out=16'h5;
17'h18671:	data_out=16'h8005;
17'h18672:	data_out=16'h5;
17'h18673:	data_out=16'h7;
17'h18674:	data_out=16'h8001;
17'h18675:	data_out=16'h8001;
17'h18676:	data_out=16'h8007;
17'h18677:	data_out=16'h5;
17'h18678:	data_out=16'h8001;
17'h18679:	data_out=16'h8002;
17'h1867a:	data_out=16'h8004;
17'h1867b:	data_out=16'h7;
17'h1867c:	data_out=16'h5;
17'h1867d:	data_out=16'h8002;
17'h1867e:	data_out=16'h8003;
17'h1867f:	data_out=16'h3;
17'h18680:	data_out=16'h2;
17'h18681:	data_out=16'h8004;
17'h18682:	data_out=16'h8004;
17'h18683:	data_out=16'h7;
17'h18684:	data_out=16'h8005;
17'h18685:	data_out=16'h8007;
17'h18686:	data_out=16'h8000;
17'h18687:	data_out=16'h6;
17'h18688:	data_out=16'h8001;
17'h18689:	data_out=16'h8004;
17'h1868a:	data_out=16'h8002;
17'h1868b:	data_out=16'h8009;
17'h1868c:	data_out=16'h8007;
17'h1868d:	data_out=16'h5;
17'h1868e:	data_out=16'h8002;
17'h1868f:	data_out=16'h7;
17'h18690:	data_out=16'h9;
17'h18691:	data_out=16'h8006;
17'h18692:	data_out=16'h5;
17'h18693:	data_out=16'h8001;
17'h18694:	data_out=16'h2;
17'h18695:	data_out=16'h7;
17'h18696:	data_out=16'h8005;
17'h18697:	data_out=16'h8007;
17'h18698:	data_out=16'h8004;
17'h18699:	data_out=16'h8000;
17'h1869a:	data_out=16'h9;
17'h1869b:	data_out=16'h8008;
17'h1869c:	data_out=16'h6;
17'h1869d:	data_out=16'h8003;
17'h1869e:	data_out=16'h4;
17'h1869f:	data_out=16'h8000;
17'h186a0:	data_out=16'h2;
17'h186a1:	data_out=16'h8009;
17'h186a2:	data_out=16'h8003;
17'h186a3:	data_out=16'h6;
17'h186a4:	data_out=16'h8006;
17'h186a5:	data_out=16'h6;
17'h186a6:	data_out=16'h2;
17'h186a7:	data_out=16'h1;
17'h186a8:	data_out=16'h8007;
17'h186a9:	data_out=16'h9;
17'h186aa:	data_out=16'h2;
17'h186ab:	data_out=16'h8005;
17'h186ac:	data_out=16'h5;
17'h186ad:	data_out=16'h9;
17'h186ae:	data_out=16'h8007;
17'h186af:	data_out=16'h5;
17'h186b0:	data_out=16'h8006;
17'h186b1:	data_out=16'h7;
17'h186b2:	data_out=16'h8006;
17'h186b3:	data_out=16'h6;
17'h186b4:	data_out=16'h5;
17'h186b5:	data_out=16'h8002;
17'h186b6:	data_out=16'h7;
17'h186b7:	data_out=16'h8007;
17'h186b8:	data_out=16'h7;
17'h186b9:	data_out=16'h7;
17'h186ba:	data_out=16'h8006;
17'h186bb:	data_out=16'h4;
17'h186bc:	data_out=16'h8006;
17'h186bd:	data_out=16'h7;
17'h186be:	data_out=16'h8006;
17'h186bf:	data_out=16'h6;
17'h186c0:	data_out=16'h7;
17'h186c1:	data_out=16'h1;
17'h186c2:	data_out=16'h2;
17'h186c3:	data_out=16'h8008;
17'h186c4:	data_out=16'h8003;
17'h186c5:	data_out=16'h8005;
17'h186c6:	data_out=16'h2;
17'h186c7:	data_out=16'h8000;
17'h186c8:	data_out=16'h8005;
17'h186c9:	data_out=16'h8005;
17'h186ca:	data_out=16'h4;
17'h186cb:	data_out=16'h8009;
17'h186cc:	data_out=16'h8005;
17'h186cd:	data_out=16'h6;
17'h186ce:	data_out=16'h5;
17'h186cf:	data_out=16'h8002;
17'h186d0:	data_out=16'h4;
17'h186d1:	data_out=16'h8;
17'h186d2:	data_out=16'h8006;
17'h186d3:	data_out=16'h0;
17'h186d4:	data_out=16'h8003;
17'h186d5:	data_out=16'h8007;
17'h186d6:	data_out=16'h2;
17'h186d7:	data_out=16'h8006;
17'h186d8:	data_out=16'h9;
17'h186d9:	data_out=16'h5;
17'h186da:	data_out=16'h7;
17'h186db:	data_out=16'h8006;
17'h186dc:	data_out=16'h3;
17'h186dd:	data_out=16'h8008;
17'h186de:	data_out=16'h9;
17'h186df:	data_out=16'h1;
17'h186e0:	data_out=16'h2;
17'h186e1:	data_out=16'h2;
17'h186e2:	data_out=16'h2;
17'h186e3:	data_out=16'h8;
17'h186e4:	data_out=16'h6;
17'h186e5:	data_out=16'h8005;
17'h186e6:	data_out=16'h8001;
17'h186e7:	data_out=16'h8008;
17'h186e8:	data_out=16'h8001;
17'h186e9:	data_out=16'h8007;
17'h186ea:	data_out=16'h8007;
17'h186eb:	data_out=16'h3;
17'h186ec:	data_out=16'h8;
17'h186ed:	data_out=16'h6;
17'h186ee:	data_out=16'h8008;
17'h186ef:	data_out=16'h3;
17'h186f0:	data_out=16'h5;
17'h186f1:	data_out=16'h8004;
17'h186f2:	data_out=16'h8006;
17'h186f3:	data_out=16'h8007;
17'h186f4:	data_out=16'h8003;
17'h186f5:	data_out=16'h5;
17'h186f6:	data_out=16'h8004;
17'h186f7:	data_out=16'h8003;
17'h186f8:	data_out=16'h1;
17'h186f9:	data_out=16'h8006;
17'h186fa:	data_out=16'h8000;
17'h186fb:	data_out=16'h8005;
17'h186fc:	data_out=16'h8005;
17'h186fd:	data_out=16'h8001;
17'h186fe:	data_out=16'h5;
17'h186ff:	data_out=16'h6;
17'h18700:	data_out=16'h8008;
17'h18701:	data_out=16'h8002;
17'h18702:	data_out=16'h5;
17'h18703:	data_out=16'h7;
17'h18704:	data_out=16'h2;
17'h18705:	data_out=16'h8006;
17'h18706:	data_out=16'h9;
17'h18707:	data_out=16'h8008;
17'h18708:	data_out=16'h8003;
17'h18709:	data_out=16'h8008;
17'h1870a:	data_out=16'h4;
17'h1870b:	data_out=16'h8004;
17'h1870c:	data_out=16'h8;
17'h1870d:	data_out=16'h5;
17'h1870e:	data_out=16'h8;
17'h1870f:	data_out=16'h4;
17'h18710:	data_out=16'h8008;
17'h18711:	data_out=16'h8007;
17'h18712:	data_out=16'h6;
17'h18713:	data_out=16'h8002;
17'h18714:	data_out=16'h8;
17'h18715:	data_out=16'h8007;
17'h18716:	data_out=16'h4;
17'h18717:	data_out=16'h8000;
17'h18718:	data_out=16'h8004;
17'h18719:	data_out=16'h8005;
17'h1871a:	data_out=16'h3;
17'h1871b:	data_out=16'h8000;
17'h1871c:	data_out=16'h3;
17'h1871d:	data_out=16'h8001;
17'h1871e:	data_out=16'h8004;
17'h1871f:	data_out=16'h5;
17'h18720:	data_out=16'h6;
17'h18721:	data_out=16'h8008;
17'h18722:	data_out=16'h3;
17'h18723:	data_out=16'h8002;
17'h18724:	data_out=16'h8005;
17'h18725:	data_out=16'h3;
17'h18726:	data_out=16'h8001;
17'h18727:	data_out=16'h1;
17'h18728:	data_out=16'h4;
17'h18729:	data_out=16'h8006;
17'h1872a:	data_out=16'h6;
17'h1872b:	data_out=16'h3;
17'h1872c:	data_out=16'h9;
17'h1872d:	data_out=16'h5;
17'h1872e:	data_out=16'h8002;
17'h1872f:	data_out=16'h8009;
17'h18730:	data_out=16'h7;
17'h18731:	data_out=16'h8005;
17'h18732:	data_out=16'h8001;
17'h18733:	data_out=16'h6;
17'h18734:	data_out=16'h8003;
17'h18735:	data_out=16'h8006;
17'h18736:	data_out=16'h8004;
17'h18737:	data_out=16'h1;
17'h18738:	data_out=16'h8002;
17'h18739:	data_out=16'h9;
17'h1873a:	data_out=16'h8008;
17'h1873b:	data_out=16'h8008;
17'h1873c:	data_out=16'h8001;
17'h1873d:	data_out=16'h8003;
17'h1873e:	data_out=16'h6;
17'h1873f:	data_out=16'h8005;
17'h18740:	data_out=16'h8002;
17'h18741:	data_out=16'h8001;
17'h18742:	data_out=16'h3;
17'h18743:	data_out=16'h2;
17'h18744:	data_out=16'h8007;
17'h18745:	data_out=16'h8007;
17'h18746:	data_out=16'h8007;
17'h18747:	data_out=16'h6;
17'h18748:	data_out=16'h8004;
17'h18749:	data_out=16'h8;
17'h1874a:	data_out=16'h8000;
17'h1874b:	data_out=16'h8005;
17'h1874c:	data_out=16'h4;
17'h1874d:	data_out=16'h7;
17'h1874e:	data_out=16'h8004;
17'h1874f:	data_out=16'h2;
17'h18750:	data_out=16'h8008;
17'h18751:	data_out=16'h3;
17'h18752:	data_out=16'h8002;
17'h18753:	data_out=16'h8002;
17'h18754:	data_out=16'h6;
17'h18755:	data_out=16'h4;
17'h18756:	data_out=16'h8;
17'h18757:	data_out=16'h8005;
17'h18758:	data_out=16'h3;
17'h18759:	data_out=16'h8009;
17'h1875a:	data_out=16'h8004;
17'h1875b:	data_out=16'h8007;
17'h1875c:	data_out=16'h8003;
17'h1875d:	data_out=16'h8008;
17'h1875e:	data_out=16'h8003;
17'h1875f:	data_out=16'h4;
17'h18760:	data_out=16'h1;
17'h18761:	data_out=16'h9;
17'h18762:	data_out=16'h8003;
17'h18763:	data_out=16'h2;
17'h18764:	data_out=16'h8008;
17'h18765:	data_out=16'h8001;
17'h18766:	data_out=16'h8001;
17'h18767:	data_out=16'h8003;
17'h18768:	data_out=16'h8002;
17'h18769:	data_out=16'h8;
17'h1876a:	data_out=16'h1;
17'h1876b:	data_out=16'h8007;
17'h1876c:	data_out=16'h6;
17'h1876d:	data_out=16'h6;
17'h1876e:	data_out=16'h4;
17'h1876f:	data_out=16'h7;
17'h18770:	data_out=16'h1;
17'h18771:	data_out=16'h8007;
17'h18772:	data_out=16'h8004;
17'h18773:	data_out=16'h8002;
17'h18774:	data_out=16'h6;
17'h18775:	data_out=16'h8005;
17'h18776:	data_out=16'h2;
17'h18777:	data_out=16'h8000;
17'h18778:	data_out=16'h8005;
17'h18779:	data_out=16'h7;
17'h1877a:	data_out=16'h2;
17'h1877b:	data_out=16'h2;
17'h1877c:	data_out=16'h8;
17'h1877d:	data_out=16'h8;
17'h1877e:	data_out=16'h8003;
17'h1877f:	data_out=16'h8001;
17'h18780:	data_out=16'h8;
17'h18781:	data_out=16'h3;
17'h18782:	data_out=16'h8007;
17'h18783:	data_out=16'h9;
17'h18784:	data_out=16'h8007;
17'h18785:	data_out=16'h1;
17'h18786:	data_out=16'h8003;
17'h18787:	data_out=16'h0;
17'h18788:	data_out=16'h0;
17'h18789:	data_out=16'h7;
17'h1878a:	data_out=16'h2;
17'h1878b:	data_out=16'h8003;
17'h1878c:	data_out=16'h5;
17'h1878d:	data_out=16'h8003;
17'h1878e:	data_out=16'h8005;
17'h1878f:	data_out=16'h8004;
17'h18790:	data_out=16'h8001;
17'h18791:	data_out=16'h0;
17'h18792:	data_out=16'h3;
17'h18793:	data_out=16'h8005;
17'h18794:	data_out=16'h5;
17'h18795:	data_out=16'h8005;
17'h18796:	data_out=16'h4;
17'h18797:	data_out=16'h8009;
17'h18798:	data_out=16'h8007;
17'h18799:	data_out=16'h8003;
17'h1879a:	data_out=16'h2;
17'h1879b:	data_out=16'h8008;
17'h1879c:	data_out=16'h8004;
17'h1879d:	data_out=16'h8;
17'h1879e:	data_out=16'h0;
17'h1879f:	data_out=16'h8006;
17'h187a0:	data_out=16'h1;
17'h187a1:	data_out=16'h2;
17'h187a2:	data_out=16'h8006;
17'h187a3:	data_out=16'h3;
17'h187a4:	data_out=16'h8006;
17'h187a5:	data_out=16'h8000;
17'h187a6:	data_out=16'h8006;
17'h187a7:	data_out=16'h4;
17'h187a8:	data_out=16'h8002;
17'h187a9:	data_out=16'h5;
17'h187aa:	data_out=16'h8008;
17'h187ab:	data_out=16'h8007;
17'h187ac:	data_out=16'h8007;
17'h187ad:	data_out=16'h8004;
17'h187ae:	data_out=16'h8002;
17'h187af:	data_out=16'h1;
17'h187b0:	data_out=16'h6;
17'h187b1:	data_out=16'h8008;
17'h187b2:	data_out=16'h5;
17'h187b3:	data_out=16'h1;
17'h187b4:	data_out=16'h8003;
17'h187b5:	data_out=16'h0;
17'h187b6:	data_out=16'h2;
17'h187b7:	data_out=16'h8001;
17'h187b8:	data_out=16'h6;
17'h187b9:	data_out=16'h8006;
17'h187ba:	data_out=16'h8000;
17'h187bb:	data_out=16'h8007;
17'h187bc:	data_out=16'h8007;
17'h187bd:	data_out=16'h9;
17'h187be:	data_out=16'h8004;
17'h187bf:	data_out=16'h3;
17'h187c0:	data_out=16'h2;
17'h187c1:	data_out=16'h8002;
17'h187c2:	data_out=16'h8003;
17'h187c3:	data_out=16'h6;
17'h187c4:	data_out=16'h7;
17'h187c5:	data_out=16'h0;
17'h187c6:	data_out=16'h0;
17'h187c7:	data_out=16'h8004;
17'h187c8:	data_out=16'h8003;
17'h187c9:	data_out=16'h1;
17'h187ca:	data_out=16'h8002;
17'h187cb:	data_out=16'h8001;
17'h187cc:	data_out=16'h6;
17'h187cd:	data_out=16'h6;
17'h187ce:	data_out=16'h9;
17'h187cf:	data_out=16'h3;
17'h187d0:	data_out=16'h7;
17'h187d1:	data_out=16'h5;
17'h187d2:	data_out=16'h8005;
17'h187d3:	data_out=16'h8005;
17'h187d4:	data_out=16'h8004;
17'h187d5:	data_out=16'h6;
17'h187d6:	data_out=16'h2;
17'h187d7:	data_out=16'h8007;
17'h187d8:	data_out=16'h8009;
17'h187d9:	data_out=16'h8007;
17'h187da:	data_out=16'h8006;
17'h187db:	data_out=16'h8007;
17'h187dc:	data_out=16'h8007;
17'h187dd:	data_out=16'h8001;
17'h187de:	data_out=16'h6;
17'h187df:	data_out=16'h4;
17'h187e0:	data_out=16'h7;
17'h187e1:	data_out=16'h8006;
17'h187e2:	data_out=16'h0;
17'h187e3:	data_out=16'h5;
17'h187e4:	data_out=16'h3;
17'h187e5:	data_out=16'h8009;
17'h187e6:	data_out=16'h8008;
17'h187e7:	data_out=16'h9;
17'h187e8:	data_out=16'h2;
17'h187e9:	data_out=16'h8001;
17'h187ea:	data_out=16'h8001;
17'h187eb:	data_out=16'h8001;
17'h187ec:	data_out=16'h8004;
17'h187ed:	data_out=16'h8002;
17'h187ee:	data_out=16'h8008;
17'h187ef:	data_out=16'h8006;
17'h187f0:	data_out=16'h8006;
17'h187f1:	data_out=16'h8004;
17'h187f2:	data_out=16'h8002;
17'h187f3:	data_out=16'h8001;
17'h187f4:	data_out=16'h8007;
17'h187f5:	data_out=16'h8009;
17'h187f6:	data_out=16'h1;
17'h187f7:	data_out=16'h8007;
17'h187f8:	data_out=16'h8007;
17'h187f9:	data_out=16'h4;
17'h187fa:	data_out=16'h8004;
17'h187fb:	data_out=16'h8005;
17'h187fc:	data_out=16'h8006;
17'h187fd:	data_out=16'h8007;
		default: #7 data_out=32'hFFFF;
	endcase
end
endmodule


module ReadOnlyMemory_WHO(output reg [15:0] data_out, input [16:0] address);
always@(address)begin
	case(address) 
17'h0:	data_out=16'h266;
17'h1:	data_out=16'h720;
17'h2:	data_out=16'h1c4;
17'h3:	data_out=16'h864f;
17'h4:	data_out=16'h8a00;
17'h5:	data_out=16'h7ca;
17'h6:	data_out=16'h8a00;
17'h7:	data_out=16'h6cc;
17'h8:	data_out=16'h84ca;
17'h9:	data_out=16'h8406;
17'ha:	data_out=16'h221;
17'hb:	data_out=16'h1d0;
17'hc:	data_out=16'h828e;
17'hd:	data_out=16'h3f;
17'he:	data_out=16'h8a00;
17'hf:	data_out=16'h2c;
17'h10:	data_out=16'h8a00;
17'h11:	data_out=16'h99;
17'h12:	data_out=16'h20;
17'h13:	data_out=16'h89fc;
17'h14:	data_out=16'h8a00;
17'h15:	data_out=16'h8a00;
17'h16:	data_out=16'h8a00;
17'h17:	data_out=16'h8309;
17'h18:	data_out=16'h14e;
17'h19:	data_out=16'h3c5;
17'h1a:	data_out=16'h8a00;
17'h1b:	data_out=16'h136;
17'h1c:	data_out=16'h8577;
17'h1d:	data_out=16'h825f;
17'h1e:	data_out=16'h8a00;
17'h1f:	data_out=16'h94d;
17'h20:	data_out=16'h88ca;
17'h21:	data_out=16'h8a00;
17'h22:	data_out=16'h8597;
17'h23:	data_out=16'h865d;
17'h24:	data_out=16'h8763;
17'h25:	data_out=16'h81ee;
17'h26:	data_out=16'h8a00;
17'h27:	data_out=16'h4c3;
17'h28:	data_out=16'h838b;
17'h29:	data_out=16'h8484;
17'h2a:	data_out=16'h8d2;
17'h2b:	data_out=16'h8277;
17'h2c:	data_out=16'h8a00;
17'h2d:	data_out=16'h82d;
17'h2e:	data_out=16'h2c3;
17'h2f:	data_out=16'h8a00;
17'h30:	data_out=16'h86ec;
17'h31:	data_out=16'h8a00;
17'h32:	data_out=16'h8a00;
17'h33:	data_out=16'h9ff;
17'h34:	data_out=16'h8420;
17'h35:	data_out=16'h2fd;
17'h36:	data_out=16'h8a00;
17'h37:	data_out=16'hd0;
17'h38:	data_out=16'h5e;
17'h39:	data_out=16'h8a00;
17'h3a:	data_out=16'h825e;
17'h3b:	data_out=16'h8a00;
17'h3c:	data_out=16'h8a00;
17'h3d:	data_out=16'h8551;
17'h3e:	data_out=16'h806a;
17'h3f:	data_out=16'h8135;
17'h40:	data_out=16'h7f6;
17'h41:	data_out=16'h899e;
17'h42:	data_out=16'h69a;
17'h43:	data_out=16'h85f2;
17'h44:	data_out=16'h845f;
17'h45:	data_out=16'h81ec;
17'h46:	data_out=16'h86b;
17'h47:	data_out=16'h8a00;
17'h48:	data_out=16'h88be;
17'h49:	data_out=16'h817f;
17'h4a:	data_out=16'h697;
17'h4b:	data_out=16'h8081;
17'h4c:	data_out=16'h96a;
17'h4d:	data_out=16'h8154;
17'h4e:	data_out=16'h8a00;
17'h4f:	data_out=16'h86d2;
17'h50:	data_out=16'h843e;
17'h51:	data_out=16'h8a00;
17'h52:	data_out=16'h864a;
17'h53:	data_out=16'h2d7;
17'h54:	data_out=16'h85bb;
17'h55:	data_out=16'h4a6;
17'h56:	data_out=16'h8a00;
17'h57:	data_out=16'h8e2;
17'h58:	data_out=16'h8a00;
17'h59:	data_out=16'h81be;
17'h5a:	data_out=16'h84d4;
17'h5b:	data_out=16'h8a00;
17'h5c:	data_out=16'h13;
17'h5d:	data_out=16'h8a00;
17'h5e:	data_out=16'h74b;
17'h5f:	data_out=16'h899b;
17'h60:	data_out=16'h521;
17'h61:	data_out=16'h85b3;
17'h62:	data_out=16'h8a00;
17'h63:	data_out=16'h8049;
17'h64:	data_out=16'ha00;
17'h65:	data_out=16'h142;
17'h66:	data_out=16'h2;
17'h67:	data_out=16'h8888;
17'h68:	data_out=16'h8a00;
17'h69:	data_out=16'h11e;
17'h6a:	data_out=16'h869d;
17'h6b:	data_out=16'h8a00;
17'h6c:	data_out=16'h759;
17'h6d:	data_out=16'h89ff;
17'h6e:	data_out=16'h7bf;
17'h6f:	data_out=16'h8a00;
17'h70:	data_out=16'h815e;
17'h71:	data_out=16'h8282;
17'h72:	data_out=16'h8526;
17'h73:	data_out=16'h8a00;
17'h74:	data_out=16'h8a00;
17'h75:	data_out=16'h4f6;
17'h76:	data_out=16'h89ff;
17'h77:	data_out=16'h6ce;
17'h78:	data_out=16'h8e7;
17'h79:	data_out=16'h8a00;
17'h7a:	data_out=16'h8a00;
17'h7b:	data_out=16'h835a;
17'h7c:	data_out=16'h83ba;
17'h7d:	data_out=16'h85b5;
17'h7e:	data_out=16'h866;
17'h7f:	data_out=16'h612;
17'h80:	data_out=16'h8a00;
17'h81:	data_out=16'h82c6;
17'h82:	data_out=16'h8791;
17'h83:	data_out=16'h89a;
17'h84:	data_out=16'h8a00;
17'h85:	data_out=16'h8409;
17'h86:	data_out=16'h376;
17'h87:	data_out=16'h2d4;
17'h88:	data_out=16'h829f;
17'h89:	data_out=16'h60;
17'h8a:	data_out=16'h8990;
17'h8b:	data_out=16'h2f8;
17'h8c:	data_out=16'h8691;
17'h8d:	data_out=16'h84a6;
17'h8e:	data_out=16'h825a;
17'h8f:	data_out=16'h8198;
17'h90:	data_out=16'h204;
17'h91:	data_out=16'h396;
17'h92:	data_out=16'h83fc;
17'h93:	data_out=16'h8387;
17'h94:	data_out=16'h2a2;
17'h95:	data_out=16'h8056;
17'h96:	data_out=16'h8a00;
17'h97:	data_out=16'h8a00;
17'h98:	data_out=16'h89fd;
17'h99:	data_out=16'h8732;
17'h9a:	data_out=16'h3ac;
17'h9b:	data_out=16'h8053;
17'h9c:	data_out=16'h8a00;
17'h9d:	data_out=16'h61a;
17'h9e:	data_out=16'h8a00;
17'h9f:	data_out=16'h865c;
17'ha0:	data_out=16'h89b6;
17'ha1:	data_out=16'h8a00;
17'ha2:	data_out=16'h73d;
17'ha3:	data_out=16'h8a00;
17'ha4:	data_out=16'h876f;
17'ha5:	data_out=16'h87c0;
17'ha6:	data_out=16'h66c;
17'ha7:	data_out=16'h49;
17'ha8:	data_out=16'h8a00;
17'ha9:	data_out=16'h63d;
17'haa:	data_out=16'h64d;
17'hab:	data_out=16'h8a00;
17'hac:	data_out=16'h9f5;
17'had:	data_out=16'h811f;
17'hae:	data_out=16'h8a00;
17'haf:	data_out=16'h8367;
17'hb0:	data_out=16'h8a00;
17'hb1:	data_out=16'h87ec;
17'hb2:	data_out=16'h13f;
17'hb3:	data_out=16'h870c;
17'hb4:	data_out=16'h8856;
17'hb5:	data_out=16'h81cc;
17'hb6:	data_out=16'h8526;
17'hb7:	data_out=16'h8220;
17'hb8:	data_out=16'h4d8;
17'hb9:	data_out=16'h181;
17'hba:	data_out=16'h89fd;
17'hbb:	data_out=16'h8d9;
17'hbc:	data_out=16'h896b;
17'hbd:	data_out=16'h8230;
17'hbe:	data_out=16'h89f7;
17'hbf:	data_out=16'h9f4;
17'hc0:	data_out=16'h85d8;
17'hc1:	data_out=16'h887c;
17'hc2:	data_out=16'h168;
17'hc3:	data_out=16'h826e;
17'hc4:	data_out=16'h893b;
17'hc5:	data_out=16'h8222;
17'hc6:	data_out=16'h8867;
17'hc7:	data_out=16'h107;
17'hc8:	data_out=16'h8a00;
17'hc9:	data_out=16'h40f;
17'hca:	data_out=16'h85c3;
17'hcb:	data_out=16'h820f;
17'hcc:	data_out=16'h8127;
17'hcd:	data_out=16'h8751;
17'hce:	data_out=16'h8a00;
17'hcf:	data_out=16'h82dc;
17'hd0:	data_out=16'h8a00;
17'hd1:	data_out=16'h2a7;
17'hd2:	data_out=16'h81e7;
17'hd3:	data_out=16'h2a3;
17'hd4:	data_out=16'h19;
17'hd5:	data_out=16'h8237;
17'hd6:	data_out=16'h81fa;
17'hd7:	data_out=16'h236;
17'hd8:	data_out=16'h81fc;
17'hd9:	data_out=16'h820b;
17'hda:	data_out=16'h82b2;
17'hdb:	data_out=16'h8217;
17'hdc:	data_out=16'h8433;
17'hdd:	data_out=16'ha00;
17'hde:	data_out=16'h8464;
17'hdf:	data_out=16'h862c;
17'he0:	data_out=16'h8471;
17'he1:	data_out=16'h81;
17'he2:	data_out=16'h8337;
17'he3:	data_out=16'h8413;
17'he4:	data_out=16'h87c1;
17'he5:	data_out=16'h8429;
17'he6:	data_out=16'h8a00;
17'he7:	data_out=16'h8c3;
17'he8:	data_out=16'h8a00;
17'he9:	data_out=16'h81c1;
17'hea:	data_out=16'h82bc;
17'heb:	data_out=16'h8a00;
17'hec:	data_out=16'h8a00;
17'hed:	data_out=16'h8118;
17'hee:	data_out=16'h8a00;
17'hef:	data_out=16'h299;
17'hf0:	data_out=16'h81cb;
17'hf1:	data_out=16'h8163;
17'hf2:	data_out=16'h8022;
17'hf3:	data_out=16'hf;
17'hf4:	data_out=16'h1bd;
17'hf5:	data_out=16'h200;
17'hf6:	data_out=16'h81f4;
17'hf7:	data_out=16'hf2;
17'hf8:	data_out=16'h8214;
17'hf9:	data_out=16'h814a;
17'hfa:	data_out=16'h9fe;
17'hfb:	data_out=16'h8a00;
17'hfc:	data_out=16'ha00;
17'hfd:	data_out=16'ha00;
17'hfe:	data_out=16'h8a00;
17'hff:	data_out=16'h89fd;
17'h100:	data_out=16'h5e2;
17'h101:	data_out=16'h831e;
17'h102:	data_out=16'h5ad;
17'h103:	data_out=16'h82c0;
17'h104:	data_out=16'h8a00;
17'h105:	data_out=16'h34f;
17'h106:	data_out=16'hd8;
17'h107:	data_out=16'h372;
17'h108:	data_out=16'h8a00;
17'h109:	data_out=16'h5a;
17'h10a:	data_out=16'h4b8;
17'h10b:	data_out=16'h8a00;
17'h10c:	data_out=16'h8177;
17'h10d:	data_out=16'h8a00;
17'h10e:	data_out=16'h89e6;
17'h10f:	data_out=16'h85cc;
17'h110:	data_out=16'h8a00;
17'h111:	data_out=16'h8011;
17'h112:	data_out=16'h833f;
17'h113:	data_out=16'h8262;
17'h114:	data_out=16'h8a00;
17'h115:	data_out=16'h8012;
17'h116:	data_out=16'h89d0;
17'h117:	data_out=16'h4cc;
17'h118:	data_out=16'h8a00;
17'h119:	data_out=16'h9f9;
17'h11a:	data_out=16'h8712;
17'h11b:	data_out=16'h81ba;
17'h11c:	data_out=16'h87e2;
17'h11d:	data_out=16'h815f;
17'h11e:	data_out=16'h8a00;
17'h11f:	data_out=16'h8120;
17'h120:	data_out=16'h8519;
17'h121:	data_out=16'h4af;
17'h122:	data_out=16'h998;
17'h123:	data_out=16'h81f6;
17'h124:	data_out=16'h159;
17'h125:	data_out=16'h8037;
17'h126:	data_out=16'h8a00;
17'h127:	data_out=16'h8423;
17'h128:	data_out=16'h8a00;
17'h129:	data_out=16'h63;
17'h12a:	data_out=16'h8094;
17'h12b:	data_out=16'h89f9;
17'h12c:	data_out=16'h8a00;
17'h12d:	data_out=16'hca;
17'h12e:	data_out=16'h83eb;
17'h12f:	data_out=16'h85d7;
17'h130:	data_out=16'h80ba;
17'h131:	data_out=16'h82d8;
17'h132:	data_out=16'h8a00;
17'h133:	data_out=16'h7;
17'h134:	data_out=16'h8a00;
17'h135:	data_out=16'h820d;
17'h136:	data_out=16'h8a00;
17'h137:	data_out=16'h8104;
17'h138:	data_out=16'h60;
17'h139:	data_out=16'h807d;
17'h13a:	data_out=16'ha00;
17'h13b:	data_out=16'h87ca;
17'h13c:	data_out=16'h8917;
17'h13d:	data_out=16'h8a00;
17'h13e:	data_out=16'h8a00;
17'h13f:	data_out=16'h86a6;
17'h140:	data_out=16'h888c;
17'h141:	data_out=16'hcc;
17'h142:	data_out=16'h83f;
17'h143:	data_out=16'h80d0;
17'h144:	data_out=16'h8a00;
17'h145:	data_out=16'h263;
17'h146:	data_out=16'h8931;
17'h147:	data_out=16'h276;
17'h148:	data_out=16'h8a00;
17'h149:	data_out=16'h89fe;
17'h14a:	data_out=16'h86cd;
17'h14b:	data_out=16'h849d;
17'h14c:	data_out=16'h8270;
17'h14d:	data_out=16'h8141;
17'h14e:	data_out=16'h226;
17'h14f:	data_out=16'h328;
17'h150:	data_out=16'h8374;
17'h151:	data_out=16'h837b;
17'h152:	data_out=16'h27a;
17'h153:	data_out=16'h8040;
17'h154:	data_out=16'h8a00;
17'h155:	data_out=16'h8a00;
17'h156:	data_out=16'h1dd;
17'h157:	data_out=16'h886b;
17'h158:	data_out=16'h815a;
17'h159:	data_out=16'h85fc;
17'h15a:	data_out=16'h309;
17'h15b:	data_out=16'h119;
17'h15c:	data_out=16'h80dd;
17'h15d:	data_out=16'h3aa;
17'h15e:	data_out=16'h9ff;
17'h15f:	data_out=16'h8a00;
17'h160:	data_out=16'h8280;
17'h161:	data_out=16'h851b;
17'h162:	data_out=16'h62;
17'h163:	data_out=16'ha00;
17'h164:	data_out=16'h240;
17'h165:	data_out=16'h8715;
17'h166:	data_out=16'hd4;
17'h167:	data_out=16'h8264;
17'h168:	data_out=16'h9ff;
17'h169:	data_out=16'h8a00;
17'h16a:	data_out=16'h827e;
17'h16b:	data_out=16'h8507;
17'h16c:	data_out=16'h57;
17'h16d:	data_out=16'ha00;
17'h16e:	data_out=16'h242;
17'h16f:	data_out=16'h8712;
17'h170:	data_out=16'hbe;
17'h171:	data_out=16'h825c;
17'h172:	data_out=16'h880b;
17'h173:	data_out=16'h8a00;
17'h174:	data_out=16'ha8;
17'h175:	data_out=16'h8a00;
17'h176:	data_out=16'h430;
17'h177:	data_out=16'h8146;
17'h178:	data_out=16'h21e;
17'h179:	data_out=16'h8a00;
17'h17a:	data_out=16'h8385;
17'h17b:	data_out=16'h8064;
17'h17c:	data_out=16'h540;
17'h17d:	data_out=16'h8a00;
17'h17e:	data_out=16'h8a00;
17'h17f:	data_out=16'h8a00;
17'h180:	data_out=16'h80dc;
17'h181:	data_out=16'h122;
17'h182:	data_out=16'h8a00;
17'h183:	data_out=16'h8319;
17'h184:	data_out=16'h833f;
17'h185:	data_out=16'h425;
17'h186:	data_out=16'h291;
17'h187:	data_out=16'h8a00;
17'h188:	data_out=16'h41b;
17'h189:	data_out=16'h34c;
17'h18a:	data_out=16'h8a00;
17'h18b:	data_out=16'h72;
17'h18c:	data_out=16'h8a00;
17'h18d:	data_out=16'h8118;
17'h18e:	data_out=16'h8a00;
17'h18f:	data_out=16'h89fe;
17'h190:	data_out=16'h879f;
17'h191:	data_out=16'h84fd;
17'h192:	data_out=16'h82e0;
17'h193:	data_out=16'h8074;
17'h194:	data_out=16'h215;
17'h195:	data_out=16'h281;
17'h196:	data_out=16'h8331;
17'h197:	data_out=16'h83c0;
17'h198:	data_out=16'h22c;
17'h199:	data_out=16'h8027;
17'h19a:	data_out=16'h8819;
17'h19b:	data_out=16'h87ad;
17'h19c:	data_out=16'h89fc;
17'h19d:	data_out=16'h885d;
17'h19e:	data_out=16'h6b8;
17'h19f:	data_out=16'h88a4;
17'h1a0:	data_out=16'h8a00;
17'h1a1:	data_out=16'h9fa;
17'h1a2:	data_out=16'h853;
17'h1a3:	data_out=16'ha00;
17'h1a4:	data_out=16'h889c;
17'h1a5:	data_out=16'h8a00;
17'h1a6:	data_out=16'h8a00;
17'h1a7:	data_out=16'h89ff;
17'h1a8:	data_out=16'h82a0;
17'h1a9:	data_out=16'h80f5;
17'h1aa:	data_out=16'h8a00;
17'h1ab:	data_out=16'ha00;
17'h1ac:	data_out=16'h89fe;
17'h1ad:	data_out=16'h89c1;
17'h1ae:	data_out=16'h9ff;
17'h1af:	data_out=16'h8a00;
17'h1b0:	data_out=16'ha00;
17'h1b1:	data_out=16'ha00;
17'h1b2:	data_out=16'h88bb;
17'h1b3:	data_out=16'h88d2;
17'h1b4:	data_out=16'h8a00;
17'h1b5:	data_out=16'h4ce;
17'h1b6:	data_out=16'h89f7;
17'h1b7:	data_out=16'h81ae;
17'h1b8:	data_out=16'h83b9;
17'h1b9:	data_out=16'h9ed;
17'h1ba:	data_out=16'h82b1;
17'h1bb:	data_out=16'h859d;
17'h1bc:	data_out=16'h8425;
17'h1bd:	data_out=16'h81;
17'h1be:	data_out=16'h82de;
17'h1bf:	data_out=16'h845e;
17'h1c0:	data_out=16'h8720;
17'h1c1:	data_out=16'h83e9;
17'h1c2:	data_out=16'h9ff;
17'h1c3:	data_out=16'h83b7;
17'h1c4:	data_out=16'h82a7;
17'h1c5:	data_out=16'h861a;
17'h1c6:	data_out=16'h848c;
17'h1c7:	data_out=16'h8458;
17'h1c8:	data_out=16'h8a00;
17'h1c9:	data_out=16'ha00;
17'h1ca:	data_out=16'h391;
17'h1cb:	data_out=16'h8032;
17'h1cc:	data_out=16'h8a00;
17'h1cd:	data_out=16'h89a3;
17'h1ce:	data_out=16'h8813;
17'h1cf:	data_out=16'h858a;
17'h1d0:	data_out=16'h573;
17'h1d1:	data_out=16'h8a00;
17'h1d2:	data_out=16'h8a00;
17'h1d3:	data_out=16'h5a4;
17'h1d4:	data_out=16'h8861;
17'h1d5:	data_out=16'h8786;
17'h1d6:	data_out=16'h8a00;
17'h1d7:	data_out=16'h2d8;
17'h1d8:	data_out=16'h821d;
17'h1d9:	data_out=16'h8188;
17'h1da:	data_out=16'h8a00;
17'h1db:	data_out=16'h83c2;
17'h1dc:	data_out=16'h86c5;
17'h1dd:	data_out=16'h4c8;
17'h1de:	data_out=16'h8a00;
17'h1df:	data_out=16'h8752;
17'h1e0:	data_out=16'h81fe;
17'h1e1:	data_out=16'h878e;
17'h1e2:	data_out=16'h8568;
17'h1e3:	data_out=16'h8111;
17'h1e4:	data_out=16'h8759;
17'h1e5:	data_out=16'h19c;
17'h1e6:	data_out=16'ha00;
17'h1e7:	data_out=16'h8a00;
17'h1e8:	data_out=16'h1b2;
17'h1e9:	data_out=16'h85a7;
17'h1ea:	data_out=16'h9fd;
17'h1eb:	data_out=16'h98f;
17'h1ec:	data_out=16'h8072;
17'h1ed:	data_out=16'h34d;
17'h1ee:	data_out=16'h8a00;
17'h1ef:	data_out=16'h8108;
17'h1f0:	data_out=16'h89bf;
17'h1f1:	data_out=16'h8a00;
17'h1f2:	data_out=16'h846f;
17'h1f3:	data_out=16'h8a00;
17'h1f4:	data_out=16'h85b9;
17'h1f5:	data_out=16'h883b;
17'h1f6:	data_out=16'h844f;
17'h1f7:	data_out=16'h8104;
17'h1f8:	data_out=16'h8a00;
17'h1f9:	data_out=16'h805c;
17'h1fa:	data_out=16'ha00;
17'h1fb:	data_out=16'h8a00;
17'h1fc:	data_out=16'h24d;
17'h1fd:	data_out=16'h8a00;
17'h1fe:	data_out=16'h8a00;
17'h1ff:	data_out=16'h23a;
17'h200:	data_out=16'h80fa;
17'h201:	data_out=16'hdd;
17'h202:	data_out=16'h32;
17'h203:	data_out=16'h852e;
17'h204:	data_out=16'h8a00;
17'h205:	data_out=16'h132;
17'h206:	data_out=16'h8a00;
17'h207:	data_out=16'h198;
17'h208:	data_out=16'h9fd;
17'h209:	data_out=16'h57c;
17'h20a:	data_out=16'h81b7;
17'h20b:	data_out=16'h819f;
17'h20c:	data_out=16'h8a00;
17'h20d:	data_out=16'h81a9;
17'h20e:	data_out=16'h8a00;
17'h20f:	data_out=16'h497;
17'h210:	data_out=16'hc6;
17'h211:	data_out=16'h8a00;
17'h212:	data_out=16'h28e;
17'h213:	data_out=16'h8827;
17'h214:	data_out=16'h8038;
17'h215:	data_out=16'h8457;
17'h216:	data_out=16'h8a00;
17'h217:	data_out=16'h478;
17'h218:	data_out=16'h8a00;
17'h219:	data_out=16'h8a00;
17'h21a:	data_out=16'h8a00;
17'h21b:	data_out=16'h8a00;
17'h21c:	data_out=16'h86f1;
17'h21d:	data_out=16'h8a00;
17'h21e:	data_out=16'h84b5;
17'h21f:	data_out=16'h8205;
17'h220:	data_out=16'h8643;
17'h221:	data_out=16'h2a9;
17'h222:	data_out=16'h8a00;
17'h223:	data_out=16'h829;
17'h224:	data_out=16'h89ff;
17'h225:	data_out=16'h8586;
17'h226:	data_out=16'h89fb;
17'h227:	data_out=16'h8a00;
17'h228:	data_out=16'h8a00;
17'h229:	data_out=16'h82d0;
17'h22a:	data_out=16'h1b6;
17'h22b:	data_out=16'h14f;
17'h22c:	data_out=16'h8a00;
17'h22d:	data_out=16'h8005;
17'h22e:	data_out=16'h8539;
17'h22f:	data_out=16'h8278;
17'h230:	data_out=16'h8a00;
17'h231:	data_out=16'h42a;
17'h232:	data_out=16'h9f4;
17'h233:	data_out=16'h22f;
17'h234:	data_out=16'h8926;
17'h235:	data_out=16'h8631;
17'h236:	data_out=16'h89df;
17'h237:	data_out=16'h71e;
17'h238:	data_out=16'hfd;
17'h239:	data_out=16'h85de;
17'h23a:	data_out=16'h8a00;
17'h23b:	data_out=16'h1ef;
17'h23c:	data_out=16'h6d;
17'h23d:	data_out=16'h803e;
17'h23e:	data_out=16'h8001;
17'h23f:	data_out=16'h8362;
17'h240:	data_out=16'h8a00;
17'h241:	data_out=16'h22f;
17'h242:	data_out=16'h8a00;
17'h243:	data_out=16'h1e7;
17'h244:	data_out=16'h813c;
17'h245:	data_out=16'h8a00;
17'h246:	data_out=16'h541;
17'h247:	data_out=16'h8a00;
17'h248:	data_out=16'h568;
17'h249:	data_out=16'h83cf;
17'h24a:	data_out=16'h367;
17'h24b:	data_out=16'h833e;
17'h24c:	data_out=16'h8a00;
17'h24d:	data_out=16'h81cc;
17'h24e:	data_out=16'h9d2;
17'h24f:	data_out=16'h8a00;
17'h250:	data_out=16'h8873;
17'h251:	data_out=16'h374;
17'h252:	data_out=16'h8a00;
17'h253:	data_out=16'h68d;
17'h254:	data_out=16'h430;
17'h255:	data_out=16'h8a00;
17'h256:	data_out=16'h88c1;
17'h257:	data_out=16'h8a00;
17'h258:	data_out=16'h8a00;
17'h259:	data_out=16'h8083;
17'h25a:	data_out=16'h89fe;
17'h25b:	data_out=16'h3c;
17'h25c:	data_out=16'h8a00;
17'h25d:	data_out=16'h84e5;
17'h25e:	data_out=16'h8a00;
17'h25f:	data_out=16'h8322;
17'h260:	data_out=16'h3af;
17'h261:	data_out=16'h4e3;
17'h262:	data_out=16'h8a00;
17'h263:	data_out=16'h95;
17'h264:	data_out=16'h77c;
17'h265:	data_out=16'h899b;
17'h266:	data_out=16'h88a6;
17'h267:	data_out=16'h516;
17'h268:	data_out=16'h8a00;
17'h269:	data_out=16'h8150;
17'h26a:	data_out=16'h895e;
17'h26b:	data_out=16'h887c;
17'h26c:	data_out=16'h87a9;
17'h26d:	data_out=16'h8502;
17'h26e:	data_out=16'h82e8;
17'h26f:	data_out=16'h806f;
17'h270:	data_out=16'h212;
17'h271:	data_out=16'h27f;
17'h272:	data_out=16'h8336;
17'h273:	data_out=16'h83c4;
17'h274:	data_out=16'h228;
17'h275:	data_out=16'h8029;
17'h276:	data_out=16'h8a00;
17'h277:	data_out=16'h9ff;
17'h278:	data_out=16'h8411;
17'h279:	data_out=16'h2d7;
17'h27a:	data_out=16'h8a00;
17'h27b:	data_out=16'h104;
17'h27c:	data_out=16'h58;
17'h27d:	data_out=16'h8a00;
17'h27e:	data_out=16'h824e;
17'h27f:	data_out=16'h8a00;
17'h280:	data_out=16'h89f5;
17'h281:	data_out=16'h866d;
17'h282:	data_out=16'h288;
17'h283:	data_out=16'h8520;
17'h284:	data_out=16'h8a00;
17'h285:	data_out=16'h197;
17'h286:	data_out=16'h8d6;
17'h287:	data_out=16'h8a00;
17'h288:	data_out=16'h83c9;
17'h289:	data_out=16'h8a00;
17'h28a:	data_out=16'h850c;
17'h28b:	data_out=16'h83c9;
17'h28c:	data_out=16'h8a00;
17'h28d:	data_out=16'h4e;
17'h28e:	data_out=16'h89a7;
17'h28f:	data_out=16'h713;
17'h290:	data_out=16'h89e7;
17'h291:	data_out=16'h39d;
17'h292:	data_out=16'h8942;
17'h293:	data_out=16'h168;
17'h294:	data_out=16'ha00;
17'h295:	data_out=16'h86f5;
17'h296:	data_out=16'h89fc;
17'h297:	data_out=16'h8a00;
17'h298:	data_out=16'h8922;
17'h299:	data_out=16'h84b2;
17'h29a:	data_out=16'h492;
17'h29b:	data_out=16'h1a4;
17'h29c:	data_out=16'h83f7;
17'h29d:	data_out=16'h140;
17'h29e:	data_out=16'h89fc;
17'h29f:	data_out=16'h9bc;
17'h2a0:	data_out=16'h8086;
17'h2a1:	data_out=16'h8079;
17'h2a2:	data_out=16'h803a;
17'h2a3:	data_out=16'h8a00;
17'h2a4:	data_out=16'h80ed;
17'h2a5:	data_out=16'h8a00;
17'h2a6:	data_out=16'h859a;
17'h2a7:	data_out=16'h304;
17'h2a8:	data_out=16'h1bf;
17'h2a9:	data_out=16'h10c;
17'h2aa:	data_out=16'h3fe;
17'h2ab:	data_out=16'h50e;
17'h2ac:	data_out=16'h8a00;
17'h2ad:	data_out=16'h32d;
17'h2ae:	data_out=16'h8991;
17'h2af:	data_out=16'h8a00;
17'h2b0:	data_out=16'h89f7;
17'h2b1:	data_out=16'h8a00;
17'h2b2:	data_out=16'h81fa;
17'h2b3:	data_out=16'h2fd;
17'h2b4:	data_out=16'h800a;
17'h2b5:	data_out=16'h825b;
17'h2b6:	data_out=16'h8211;
17'h2b7:	data_out=16'h231;
17'h2b8:	data_out=16'h8210;
17'h2b9:	data_out=16'h8225;
17'h2ba:	data_out=16'h82de;
17'h2bb:	data_out=16'h8230;
17'h2bc:	data_out=16'h219;
17'h2bd:	data_out=16'h8a00;
17'h2be:	data_out=16'h880e;
17'h2bf:	data_out=16'h80b0;
17'h2c0:	data_out=16'h8a00;
17'h2c1:	data_out=16'h26a;
17'h2c2:	data_out=16'h8a00;
17'h2c3:	data_out=16'h772;
17'h2c4:	data_out=16'h384;
17'h2c5:	data_out=16'h79d;
17'h2c6:	data_out=16'h102;
17'h2c7:	data_out=16'h8a00;
17'h2c8:	data_out=16'h2c9;
17'h2c9:	data_out=16'h8a00;
17'h2ca:	data_out=16'h85f;
17'h2cb:	data_out=16'h8293;
17'h2cc:	data_out=16'h838e;
17'h2cd:	data_out=16'h6f8;
17'h2ce:	data_out=16'h8a00;
17'h2cf:	data_out=16'h8358;
17'h2d0:	data_out=16'h89ff;
17'h2d1:	data_out=16'h8624;
17'h2d2:	data_out=16'h80e3;
17'h2d3:	data_out=16'h8422;
17'h2d4:	data_out=16'h14;
17'h2d5:	data_out=16'h8677;
17'h2d6:	data_out=16'h1a8;
17'h2d7:	data_out=16'h736;
17'h2d8:	data_out=16'h8a00;
17'h2d9:	data_out=16'h8698;
17'h2da:	data_out=16'h8736;
17'h2db:	data_out=16'h8a00;
17'h2dc:	data_out=16'hba;
17'h2dd:	data_out=16'h8a00;
17'h2de:	data_out=16'h6c;
17'h2df:	data_out=16'h804e;
17'h2e0:	data_out=16'h39a;
17'h2e1:	data_out=16'h89f8;
17'h2e2:	data_out=16'h8407;
17'h2e3:	data_out=16'hf1;
17'h2e4:	data_out=16'h188;
17'h2e5:	data_out=16'h89fe;
17'h2e6:	data_out=16'h8043;
17'h2e7:	data_out=16'h64b;
17'h2e8:	data_out=16'h8505;
17'h2e9:	data_out=16'h805e;
17'h2ea:	data_out=16'h2f6;
17'h2eb:	data_out=16'h680;
17'h2ec:	data_out=16'h8a00;
17'h2ed:	data_out=16'h8a00;
17'h2ee:	data_out=16'ha00;
17'h2ef:	data_out=16'h88dc;
17'h2f0:	data_out=16'h89fc;
17'h2f1:	data_out=16'h8a00;
17'h2f2:	data_out=16'h89e0;
17'h2f3:	data_out=16'h89f5;
17'h2f4:	data_out=16'ha00;
17'h2f5:	data_out=16'h728;
17'h2f6:	data_out=16'h88b7;
17'h2f7:	data_out=16'h80d7;
17'h2f8:	data_out=16'h85fb;
17'h2f9:	data_out=16'h8a00;
17'h2fa:	data_out=16'h81bc;
17'h2fb:	data_out=16'h8a00;
17'h2fc:	data_out=16'h447;
17'h2fd:	data_out=16'hbd;
17'h2fe:	data_out=16'h4c9;
17'h2ff:	data_out=16'h800a;
17'h300:	data_out=16'h2ab;
17'h301:	data_out=16'h8156;
17'h302:	data_out=16'h8a00;
17'h303:	data_out=16'h8a00;
17'h304:	data_out=16'h4bd;
17'h305:	data_out=16'h8716;
17'h306:	data_out=16'h8315;
17'h307:	data_out=16'h855a;
17'h308:	data_out=16'h496;
17'h309:	data_out=16'h44f;
17'h30a:	data_out=16'h8056;
17'h30b:	data_out=16'h63;
17'h30c:	data_out=16'h8653;
17'h30d:	data_out=16'h89fb;
17'h30e:	data_out=16'h88f3;
17'h30f:	data_out=16'h440;
17'h310:	data_out=16'h38b;
17'h311:	data_out=16'h335;
17'h312:	data_out=16'h89f9;
17'h313:	data_out=16'ha00;
17'h314:	data_out=16'h8459;
17'h315:	data_out=16'h8198;
17'h316:	data_out=16'h80f9;
17'h317:	data_out=16'h8a00;
17'h318:	data_out=16'h92;
17'h319:	data_out=16'h8a00;
17'h31a:	data_out=16'h2de;
17'h31b:	data_out=16'h8219;
17'h31c:	data_out=16'h5c3;
17'h31d:	data_out=16'h815f;
17'h31e:	data_out=16'h8110;
17'h31f:	data_out=16'h8129;
17'h320:	data_out=16'h8a00;
17'h321:	data_out=16'h9fc;
17'h322:	data_out=16'h57;
17'h323:	data_out=16'h85a4;
17'h324:	data_out=16'h86fe;
17'h325:	data_out=16'h86c1;
17'h326:	data_out=16'h32d;
17'h327:	data_out=16'h8578;
17'h328:	data_out=16'h89ed;
17'h329:	data_out=16'h82eb;
17'h32a:	data_out=16'h8a00;
17'h32b:	data_out=16'h832;
17'h32c:	data_out=16'h89ff;
17'h32d:	data_out=16'h8247;
17'h32e:	data_out=16'h6c5;
17'h32f:	data_out=16'h1e5;
17'h330:	data_out=16'h8a00;
17'h331:	data_out=16'h8768;
17'h332:	data_out=16'h8768;
17'h333:	data_out=16'h234;
17'h334:	data_out=16'ha00;
17'h335:	data_out=16'h8a00;
17'h336:	data_out=16'h8385;
17'h337:	data_out=16'h8a00;
17'h338:	data_out=16'h804d;
17'h339:	data_out=16'h5a2;
17'h33a:	data_out=16'h2c8;
17'h33b:	data_out=16'h88e9;
17'h33c:	data_out=16'h8004;
17'h33d:	data_out=16'h83a8;
17'h33e:	data_out=16'h89cf;
17'h33f:	data_out=16'h89fe;
17'h340:	data_out=16'h81f4;
17'h341:	data_out=16'ha00;
17'h342:	data_out=16'h8a00;
17'h343:	data_out=16'h83c6;
17'h344:	data_out=16'h8a00;
17'h345:	data_out=16'h53a;
17'h346:	data_out=16'h89fe;
17'h347:	data_out=16'h89fa;
17'h348:	data_out=16'h8a00;
17'h349:	data_out=16'h8502;
17'h34a:	data_out=16'h465;
17'h34b:	data_out=16'h827b;
17'h34c:	data_out=16'h8a00;
17'h34d:	data_out=16'hbe;
17'h34e:	data_out=16'h8a00;
17'h34f:	data_out=16'h994;
17'h350:	data_out=16'h8a00;
17'h351:	data_out=16'h89ff;
17'h352:	data_out=16'h8a00;
17'h353:	data_out=16'h80e4;
17'h354:	data_out=16'h8a00;
17'h355:	data_out=16'h861b;
17'h356:	data_out=16'h4d5;
17'h357:	data_out=16'h83db;
17'h358:	data_out=16'h8a00;
17'h359:	data_out=16'h8819;
17'h35a:	data_out=16'h8a00;
17'h35b:	data_out=16'h116;
17'h35c:	data_out=16'h857d;
17'h35d:	data_out=16'h8a00;
17'h35e:	data_out=16'h867a;
17'h35f:	data_out=16'h868b;
17'h360:	data_out=16'h836e;
17'h361:	data_out=16'ha00;
17'h362:	data_out=16'h89d2;
17'h363:	data_out=16'h868d;
17'h364:	data_out=16'h8482;
17'h365:	data_out=16'h1a6;
17'h366:	data_out=16'h8a00;
17'h367:	data_out=16'h8a00;
17'h368:	data_out=16'h25f;
17'h369:	data_out=16'h8a00;
17'h36a:	data_out=16'h472;
17'h36b:	data_out=16'h6db;
17'h36c:	data_out=16'h8a00;
17'h36d:	data_out=16'h8a00;
17'h36e:	data_out=16'h8346;
17'h36f:	data_out=16'h817a;
17'h370:	data_out=16'h8a00;
17'h371:	data_out=16'h1c0;
17'h372:	data_out=16'h8a00;
17'h373:	data_out=16'h2cc;
17'h374:	data_out=16'h815c;
17'h375:	data_out=16'h28a;
17'h376:	data_out=16'h8a00;
17'h377:	data_out=16'h81ad;
17'h378:	data_out=16'h84f6;
17'h379:	data_out=16'h5b9;
17'h37a:	data_out=16'h8a00;
17'h37b:	data_out=16'h84c5;
17'h37c:	data_out=16'h8b6;
17'h37d:	data_out=16'h8a00;
17'h37e:	data_out=16'h8a00;
17'h37f:	data_out=16'h158;
17'h380:	data_out=16'h5eb;
17'h381:	data_out=16'h8a00;
17'h382:	data_out=16'h8025;
17'h383:	data_out=16'h8a00;
17'h384:	data_out=16'h87b2;
17'h385:	data_out=16'h291;
17'h386:	data_out=16'h8a00;
17'h387:	data_out=16'h74a;
17'h388:	data_out=16'h802e;
17'h389:	data_out=16'h8369;
17'h38a:	data_out=16'h8a00;
17'h38b:	data_out=16'h30f;
17'h38c:	data_out=16'h8647;
17'h38d:	data_out=16'h4c9;
17'h38e:	data_out=16'h82e5;
17'h38f:	data_out=16'h8664;
17'h390:	data_out=16'h6e8;
17'h391:	data_out=16'h3d9;
17'h392:	data_out=16'h8a00;
17'h393:	data_out=16'h356;
17'h394:	data_out=16'h8a00;
17'h395:	data_out=16'h8a00;
17'h396:	data_out=16'h8552;
17'h397:	data_out=16'h8a00;
17'h398:	data_out=16'h8a00;
17'h399:	data_out=16'ha00;
17'h39a:	data_out=16'h89a6;
17'h39b:	data_out=16'h952;
17'h39c:	data_out=16'h88f6;
17'h39d:	data_out=16'h823b;
17'h39e:	data_out=16'h8a00;
17'h39f:	data_out=16'h831f;
17'h3a0:	data_out=16'h8313;
17'h3a1:	data_out=16'h8258;
17'h3a2:	data_out=16'h8972;
17'h3a3:	data_out=16'h1ba;
17'h3a4:	data_out=16'h8165;
17'h3a5:	data_out=16'h8832;
17'h3a6:	data_out=16'h89c6;
17'h3a7:	data_out=16'h80b6;
17'h3a8:	data_out=16'h848c;
17'h3a9:	data_out=16'h3a8;
17'h3aa:	data_out=16'h8706;
17'h3ab:	data_out=16'h88d0;
17'h3ac:	data_out=16'h8a00;
17'h3ad:	data_out=16'h3ce;
17'h3ae:	data_out=16'h82dd;
17'h3af:	data_out=16'h83bd;
17'h3b0:	data_out=16'h89f2;
17'h3b1:	data_out=16'h8527;
17'h3b2:	data_out=16'h851b;
17'h3b3:	data_out=16'h3ae;
17'h3b4:	data_out=16'h8972;
17'h3b5:	data_out=16'h86b9;
17'h3b6:	data_out=16'h81d7;
17'h3b7:	data_out=16'h818b;
17'h3b8:	data_out=16'hfe;
17'h3b9:	data_out=16'h8191;
17'h3ba:	data_out=16'h808a;
17'h3bb:	data_out=16'h1b;
17'h3bc:	data_out=16'h81ae;
17'h3bd:	data_out=16'h28f;
17'h3be:	data_out=16'h81ee;
17'h3bf:	data_out=16'h82a1;
17'h3c0:	data_out=16'ha00;
17'h3c1:	data_out=16'h8a00;
17'h3c2:	data_out=16'h8a00;
17'h3c3:	data_out=16'h8a00;
17'h3c4:	data_out=16'h8223;
17'h3c5:	data_out=16'h836a;
17'h3c6:	data_out=16'h8a00;
17'h3c7:	data_out=16'h832b;
17'h3c8:	data_out=16'h825b;
17'h3c9:	data_out=16'h150;
17'h3ca:	data_out=16'h88b4;
17'h3cb:	data_out=16'h8219;
17'h3cc:	data_out=16'h8352;
17'h3cd:	data_out=16'h806d;
17'h3ce:	data_out=16'h8a00;
17'h3cf:	data_out=16'h274;
17'h3d0:	data_out=16'h8337;
17'h3d1:	data_out=16'h8a00;
17'h3d2:	data_out=16'h20d;
17'h3d3:	data_out=16'h8a00;
17'h3d4:	data_out=16'h89a6;
17'h3d5:	data_out=16'h8167;
17'h3d6:	data_out=16'h89f9;
17'h3d7:	data_out=16'h873d;
17'h3d8:	data_out=16'h85f3;
17'h3d9:	data_out=16'h8a00;
17'h3da:	data_out=16'h8a00;
17'h3db:	data_out=16'h3c9;
17'h3dc:	data_out=16'h8a00;
17'h3dd:	data_out=16'h252;
17'h3de:	data_out=16'h8a00;
17'h3df:	data_out=16'h1b3;
17'h3e0:	data_out=16'h825e;
17'h3e1:	data_out=16'h245;
17'h3e2:	data_out=16'h80cf;
17'h3e3:	data_out=16'h8610;
17'h3e4:	data_out=16'h8a00;
17'h3e5:	data_out=16'h24f;
17'h3e6:	data_out=16'h8a00;
17'h3e7:	data_out=16'h8008;
17'h3e8:	data_out=16'ha00;
17'h3e9:	data_out=16'h37f;
17'h3ea:	data_out=16'h64f;
17'h3eb:	data_out=16'h8334;
17'h3ec:	data_out=16'h8a00;
17'h3ed:	data_out=16'h4f;
17'h3ee:	data_out=16'h8a00;
17'h3ef:	data_out=16'h7e9;
17'h3f0:	data_out=16'h81e4;
17'h3f1:	data_out=16'h8265;
17'h3f2:	data_out=16'h9c2;
17'h3f3:	data_out=16'h8786;
17'h3f4:	data_out=16'h7d8;
17'h3f5:	data_out=16'h6c;
17'h3f6:	data_out=16'h8a00;
17'h3f7:	data_out=16'h89fd;
17'h3f8:	data_out=16'ha00;
17'h3f9:	data_out=16'h8a00;
17'h3fa:	data_out=16'h8404;
17'h3fb:	data_out=16'h8a00;
17'h3fc:	data_out=16'h9c5;
17'h3fd:	data_out=16'h8a00;
17'h3fe:	data_out=16'h52e;
17'h3ff:	data_out=16'ha00;
17'h400:	data_out=16'h85a7;
17'h401:	data_out=16'h89f5;
17'h402:	data_out=16'h368;
17'h403:	data_out=16'h898c;
17'h404:	data_out=16'h8a00;
17'h405:	data_out=16'h8300;
17'h406:	data_out=16'h89fd;
17'h407:	data_out=16'h8a00;
17'h408:	data_out=16'ha00;
17'h409:	data_out=16'h89fd;
17'h40a:	data_out=16'h324;
17'h40b:	data_out=16'h89fa;
17'h40c:	data_out=16'h88c0;
17'h40d:	data_out=16'h498;
17'h40e:	data_out=16'h83d7;
17'h40f:	data_out=16'h8651;
17'h410:	data_out=16'h8704;
17'h411:	data_out=16'h84ad;
17'h412:	data_out=16'h8288;
17'h413:	data_out=16'h8104;
17'h414:	data_out=16'h23c;
17'h415:	data_out=16'h2d7;
17'h416:	data_out=16'h8333;
17'h417:	data_out=16'h8396;
17'h418:	data_out=16'h25d;
17'h419:	data_out=16'h802c;
17'h41a:	data_out=16'h8182;
17'h41b:	data_out=16'h8a00;
17'h41c:	data_out=16'h8789;
17'h41d:	data_out=16'h814b;
17'h41e:	data_out=16'h80a6;
17'h41f:	data_out=16'h4f7;
17'h420:	data_out=16'h8a00;
17'h421:	data_out=16'h945;
17'h422:	data_out=16'h8a00;
17'h423:	data_out=16'h438;
17'h424:	data_out=16'h8689;
17'h425:	data_out=16'h84ac;
17'h426:	data_out=16'h825e;
17'h427:	data_out=16'h81d9;
17'h428:	data_out=16'h206;
17'h429:	data_out=16'h3cf;
17'h42a:	data_out=16'h846b;
17'h42b:	data_out=16'h8393;
17'h42c:	data_out=16'h2c7;
17'h42d:	data_out=16'h8059;
17'h42e:	data_out=16'h8a00;
17'h42f:	data_out=16'h9fa;
17'h430:	data_out=16'h480;
17'h431:	data_out=16'h838a;
17'h432:	data_out=16'h8a00;
17'h433:	data_out=16'h82f2;
17'h434:	data_out=16'h8260;
17'h435:	data_out=16'h8a00;
17'h436:	data_out=16'h89f8;
17'h437:	data_out=16'h8a00;
17'h438:	data_out=16'h8;
17'h439:	data_out=16'h870;
17'h43a:	data_out=16'h8017;
17'h43b:	data_out=16'h89ad;
17'h43c:	data_out=16'h8a00;
17'h43d:	data_out=16'h73b;
17'h43e:	data_out=16'h89ff;
17'h43f:	data_out=16'h758;
17'h440:	data_out=16'h8345;
17'h441:	data_out=16'h885e;
17'h442:	data_out=16'h8a00;
17'h443:	data_out=16'h199;
17'h444:	data_out=16'h81fc;
17'h445:	data_out=16'h1c1;
17'h446:	data_out=16'h80ce;
17'h447:	data_out=16'h85d1;
17'h448:	data_out=16'h8a00;
17'h449:	data_out=16'h254;
17'h44a:	data_out=16'h8a00;
17'h44b:	data_out=16'h18;
17'h44c:	data_out=16'h8689;
17'h44d:	data_out=16'h84ac;
17'h44e:	data_out=16'h825f;
17'h44f:	data_out=16'h81d8;
17'h450:	data_out=16'h205;
17'h451:	data_out=16'h3cf;
17'h452:	data_out=16'h8468;
17'h453:	data_out=16'h8393;
17'h454:	data_out=16'h2c7;
17'h455:	data_out=16'h8059;
17'h456:	data_out=16'h8a00;
17'h457:	data_out=16'h9f2;
17'h458:	data_out=16'h8726;
17'h459:	data_out=16'h7;
17'h45a:	data_out=16'h8a00;
17'h45b:	data_out=16'h8519;
17'h45c:	data_out=16'h9ff;
17'h45d:	data_out=16'h8a00;
17'h45e:	data_out=16'h853b;
17'h45f:	data_out=16'h8a00;
17'h460:	data_out=16'h868c;
17'h461:	data_out=16'h84ab;
17'h462:	data_out=16'h825e;
17'h463:	data_out=16'h81af;
17'h464:	data_out=16'h201;
17'h465:	data_out=16'h3b3;
17'h466:	data_out=16'h8427;
17'h467:	data_out=16'h838e;
17'h468:	data_out=16'h2b2;
17'h469:	data_out=16'h8059;
17'h46a:	data_out=16'h87ed;
17'h46b:	data_out=16'h85dd;
17'h46c:	data_out=16'h88a9;
17'h46d:	data_out=16'h8475;
17'h46e:	data_out=16'h538;
17'h46f:	data_out=16'h80c3;
17'h470:	data_out=16'h8a00;
17'h471:	data_out=16'h4c3;
17'h472:	data_out=16'h8a00;
17'h473:	data_out=16'h8a00;
17'h474:	data_out=16'h8a00;
17'h475:	data_out=16'h9fa;
17'h476:	data_out=16'h508;
17'h477:	data_out=16'h896c;
17'h478:	data_out=16'h8a00;
17'h479:	data_out=16'h8230;
17'h47a:	data_out=16'h808e;
17'h47b:	data_out=16'h8a00;
17'h47c:	data_out=16'h1a;
17'h47d:	data_out=16'h8a00;
17'h47e:	data_out=16'h8a00;
17'h47f:	data_out=16'h9fb;
17'h480:	data_out=16'hc3;
17'h481:	data_out=16'h85b0;
17'h482:	data_out=16'h8a00;
17'h483:	data_out=16'h82f6;
17'h484:	data_out=16'h82b0;
17'h485:	data_out=16'h8a00;
17'h486:	data_out=16'h40a;
17'h487:	data_out=16'h8a00;
17'h488:	data_out=16'h8196;
17'h489:	data_out=16'h8757;
17'h48a:	data_out=16'h8725;
17'h48b:	data_out=16'h8127;
17'h48c:	data_out=16'h877b;
17'h48d:	data_out=16'h31c;
17'h48e:	data_out=16'ha00;
17'h48f:	data_out=16'h8a00;
17'h490:	data_out=16'h1d4;
17'h491:	data_out=16'h85b3;
17'h492:	data_out=16'h8a00;
17'h493:	data_out=16'ha00;
17'h494:	data_out=16'h89ff;
17'h495:	data_out=16'h836;
17'h496:	data_out=16'h874b;
17'h497:	data_out=16'h801b;
17'h498:	data_out=16'h85aa;
17'h499:	data_out=16'h8a00;
17'h49a:	data_out=16'h28e;
17'h49b:	data_out=16'h820b;
17'h49c:	data_out=16'h9fd;
17'h49d:	data_out=16'h8a00;
17'h49e:	data_out=16'h90e;
17'h49f:	data_out=16'h16a;
17'h4a0:	data_out=16'h844f;
17'h4a1:	data_out=16'h89ff;
17'h4a2:	data_out=16'h89fb;
17'h4a3:	data_out=16'h8401;
17'h4a4:	data_out=16'h85d7;
17'h4a5:	data_out=16'h8036;
17'h4a6:	data_out=16'h8a00;
17'h4a7:	data_out=16'h8a00;
17'h4a8:	data_out=16'h83f0;
17'h4a9:	data_out=16'h8a00;
17'h4aa:	data_out=16'h8076;
17'h4ab:	data_out=16'h84e0;
17'h4ac:	data_out=16'h2ee;
17'h4ad:	data_out=16'h808e;
17'h4ae:	data_out=16'h8a00;
17'h4af:	data_out=16'h20;
17'h4b0:	data_out=16'h8a00;
17'h4b1:	data_out=16'h9f7;
17'h4b2:	data_out=16'h8282;
17'h4b3:	data_out=16'h4e7;
17'h4b4:	data_out=16'h8a00;
17'h4b5:	data_out=16'h89eb;
17'h4b6:	data_out=16'h9fa;
17'h4b7:	data_out=16'h8820;
17'h4b8:	data_out=16'h9b9;
17'h4b9:	data_out=16'hc8;
17'h4ba:	data_out=16'h8895;
17'h4bb:	data_out=16'h8985;
17'h4bc:	data_out=16'h87fa;
17'h4bd:	data_out=16'h827a;
17'h4be:	data_out=16'h172;
17'h4bf:	data_out=16'h7c2;
17'h4c0:	data_out=16'h89d1;
17'h4c1:	data_out=16'h9fe;
17'h4c2:	data_out=16'h8706;
17'h4c3:	data_out=16'he2;
17'h4c4:	data_out=16'h8a00;
17'h4c5:	data_out=16'h23d;
17'h4c6:	data_out=16'h84f8;
17'h4c7:	data_out=16'h13;
17'h4c8:	data_out=16'h81a0;
17'h4c9:	data_out=16'h865c;
17'h4ca:	data_out=16'h8a00;
17'h4cb:	data_out=16'h92;
17'h4cc:	data_out=16'h8a00;
17'h4cd:	data_out=16'h2c;
17'h4ce:	data_out=16'h87ad;
17'h4cf:	data_out=16'h8504;
17'h4d0:	data_out=16'h82ed;
17'h4d1:	data_out=16'h806e;
17'h4d2:	data_out=16'h211;
17'h4d3:	data_out=16'h27d;
17'h4d4:	data_out=16'h8337;
17'h4d5:	data_out=16'h83c4;
17'h4d6:	data_out=16'h227;
17'h4d7:	data_out=16'h802a;
17'h4d8:	data_out=16'h8148;
17'h4d9:	data_out=16'h8146;
17'h4da:	data_out=16'h60;
17'h4db:	data_out=16'h90;
17'h4dc:	data_out=16'h131;
17'h4dd:	data_out=16'h1b8;
17'h4de:	data_out=16'h817b;
17'h4df:	data_out=16'h148;
17'h4e0:	data_out=16'h81a1;
17'h4e1:	data_out=16'h81cf;
17'h4e2:	data_out=16'h8a00;
17'h4e3:	data_out=16'h109;
17'h4e4:	data_out=16'h785;
17'h4e5:	data_out=16'h40a;
17'h4e6:	data_out=16'h5de;
17'h4e7:	data_out=16'h81b4;
17'h4e8:	data_out=16'h83ac;
17'h4e9:	data_out=16'h89ff;
17'h4ea:	data_out=16'h89fe;
17'h4eb:	data_out=16'h874c;
17'h4ec:	data_out=16'h89fd;
17'h4ed:	data_out=16'h8a00;
17'h4ee:	data_out=16'hd7;
17'h4ef:	data_out=16'h8779;
17'h4f0:	data_out=16'h66c;
17'h4f1:	data_out=16'h881a;
17'h4f2:	data_out=16'h8374;
17'h4f3:	data_out=16'h84f1;
17'h4f4:	data_out=16'h8616;
17'h4f5:	data_out=16'h4bb;
17'h4f6:	data_out=16'h8a00;
17'h4f7:	data_out=16'h693;
17'h4f8:	data_out=16'h515;
17'h4f9:	data_out=16'h8110;
17'h4fa:	data_out=16'h833e;
17'h4fb:	data_out=16'h2d4;
17'h4fc:	data_out=16'h31d;
17'h4fd:	data_out=16'h824e;
		default: #7 data_out=32'hFFFF;
	endcase
end
endmodule
